library ieee;
use ieee.std_logic_1164.all;

package myTypes is
    
    type aluOp is (LLS, LRS, ADDS, SUBS, ANDS, ORS, XORS, SNES, SLES, SGES, NOP);

end myTypes;
