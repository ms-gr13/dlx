
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_dlx is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (LLS, LRS, ADDS, SUBS, ANDS, ORS, XORS, SNES, SLES, SGES, NOP);
attribute ENUM_ENCODING of aluOp : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";

end CONV_PACK_dlx;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_6;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n13);
   U2 : INV_X1 port map( A => n16, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => S, B1 => B(2), B2 => n13, ZN => 
                           n16);
   U4 : INV_X1 port map( A => n17, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => S, A2 => A(3), B1 => B(3), B2 => n13, ZN => 
                           n17);
   U6 : INV_X1 port map( A => n15, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => S, B1 => B(1), B2 => n13, ZN => 
                           n15);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => S, B1 => B(0), B2 => n13, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_5;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n13);
   U2 : INV_X1 port map( A => n16, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => S, B1 => B(2), B2 => n13, ZN => 
                           n16);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => S, B1 => B(1), B2 => n13, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n17, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => S, A2 => A(3), B1 => B(3), B2 => n13, ZN => 
                           n17);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => S, B1 => B(0), B2 => n13, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_4;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n13);
   U2 : INV_X1 port map( A => n16, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => S, B1 => B(2), B2 => n13, ZN => 
                           n16);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => S, B1 => B(1), B2 => n13, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n17, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => S, A2 => A(3), B1 => B(3), B2 => n13, ZN => 
                           n17);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => S, B1 => B(0), B2 => n13, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_3;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n13);
   U2 : INV_X1 port map( A => n16, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => S, B1 => B(2), B2 => n13, ZN => 
                           n16);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => S, B1 => B(1), B2 => n13, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n17, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => S, A2 => A(3), B1 => B(3), B2 => n13, ZN => 
                           n17);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => S, B1 => B(0), B2 => n13, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_2;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n13);
   U2 : INV_X1 port map( A => n16, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => S, B1 => B(2), B2 => n13, ZN => 
                           n16);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => S, B1 => B(1), B2 => n13, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n17, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => S, A2 => A(3), B1 => B(3), B2 => n13, ZN => 
                           n17);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => S, B1 => B(0), B2 => n13, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_1;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n13);
   U2 : INV_X1 port map( A => n16, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => S, B1 => B(2), B2 => n13, ZN => 
                           n16);
   U4 : INV_X1 port map( A => n17, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => S, A2 => A(3), B1 => B(3), B2 => n13, ZN => 
                           n17);
   U6 : INV_X1 port map( A => n15, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => S, B1 => B(1), B2 => n13, ZN => 
                           n15);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => S, B1 => B(0), B2 => n13, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_15;

architecture SYN_BEHAVIORAL of RCA_NBITS4_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n23, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n29, A2 => n26, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n23);
   U4 : AOI21_X1 port map( B1 => n26, B2 => n29, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n28, B2 => n23, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n25, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n25);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n27, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n27);
   U11 : AOI21_X1 port map( B1 => n24, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n24);
   U13 : INV_X1 port map( A => A(0), ZN => n26);
   U14 : INV_X1 port map( A => B(0), ZN => n29);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n28);
   U20 : XNOR2_X1 port map( A => n30, B => B(2), ZN => n41);
   U21 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U22 : OAI22_X1 port map( A1 => n36, A2 => n30, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U23 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U24 : INV_X1 port map( A => Ci, ZN => n30);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_14;

architecture SYN_BEHAVIORAL of RCA_NBITS4_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n23, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n29, A2 => n26, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n23);
   U4 : AOI21_X1 port map( B1 => n26, B2 => n29, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n28, B2 => n23, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n25, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n25);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n27, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n27);
   U11 : AOI21_X1 port map( B1 => n24, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n24);
   U13 : INV_X1 port map( A => B(0), ZN => n29);
   U14 : INV_X1 port map( A => A(0), ZN => n26);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n28);
   U20 : XNOR2_X1 port map( A => n30, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n30, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U23 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U24 : INV_X1 port map( A => Ci, ZN => n30);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_13;

architecture SYN_BEHAVIORAL of RCA_NBITS4_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n23, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n29, A2 => n26, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n23);
   U4 : AOI21_X1 port map( B1 => n26, B2 => n29, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n28, B2 => n23, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n25, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n25);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n27, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n27);
   U11 : AOI21_X1 port map( B1 => n24, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n24);
   U13 : INV_X1 port map( A => B(0), ZN => n29);
   U14 : INV_X1 port map( A => A(0), ZN => n26);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n28);
   U20 : XNOR2_X1 port map( A => n30, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n30, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U23 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U24 : INV_X1 port map( A => Ci, ZN => n30);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_12;

architecture SYN_BEHAVIORAL of RCA_NBITS4_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U23 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_11;

architecture SYN_BEHAVIORAL of RCA_NBITS4_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U23 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_10;

architecture SYN_BEHAVIORAL of RCA_NBITS4_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U23 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_9;

architecture SYN_BEHAVIORAL of RCA_NBITS4_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U23 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_8;

architecture SYN_BEHAVIORAL of RCA_NBITS4_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U23 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_7;

architecture SYN_BEHAVIORAL of RCA_NBITS4_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U23 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_6;

architecture SYN_BEHAVIORAL of RCA_NBITS4_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U23 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_5;

architecture SYN_BEHAVIORAL of RCA_NBITS4_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U23 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_4;

architecture SYN_BEHAVIORAL of RCA_NBITS4_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U23 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_3;

architecture SYN_BEHAVIORAL of RCA_NBITS4_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U23 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_2;

architecture SYN_BEHAVIORAL of RCA_NBITS4_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U23 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_1;

architecture SYN_BEHAVIORAL of RCA_NBITS4_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n44, B => n43, Z => S(3));
   U26 : XOR2_X1 port map( A => n24, B => A(3), Z => n43);
   U27 : XOR2_X1 port map( A => n42, B => n41, Z => S(2));
   U28 : XOR2_X1 port map( A => n39, B => n38, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n30, A2 => n27, ZN => n37);
   U3 : INV_X1 port map( A => n33, ZN => n24);
   U4 : AOI21_X1 port map( B1 => n27, B2 => n30, A => n37, ZN => n36);
   U5 : OAI21_X1 port map( B1 => n29, B2 => n24, A => n34, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n37, B2 => A(1), A => n26, ZN => n40);
   U7 : INV_X1 port map( A => n31, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n37, B2 => A(1), A => B(1), ZN => n31);
   U9 : AOI21_X1 port map( B1 => n28, B2 => n40, A => n32, ZN => n33);
   U10 : INV_X1 port map( A => A(2), ZN => n28);
   U11 : AOI21_X1 port map( B1 => n25, B2 => A(2), A => B(2), ZN => n32);
   U12 : INV_X1 port map( A => n40, ZN => n25);
   U13 : INV_X1 port map( A => B(0), ZN => n30);
   U14 : INV_X1 port map( A => A(0), ZN => n27);
   U15 : XNOR2_X1 port map( A => A(2), B => n40, ZN => n42);
   U16 : XNOR2_X1 port map( A => n37, B => A(1), ZN => n38);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n35);
   U18 : OAI21_X1 port map( B1 => n33, B2 => A(3), A => B(3), ZN => n34);
   U19 : INV_X1 port map( A => A(3), ZN => n29);
   U20 : XNOR2_X1 port map( A => n23, B => B(2), ZN => n41);
   U21 : OAI22_X1 port map( A1 => n36, A2 => n23, B1 => Ci, B2 => n35, ZN => 
                           S(0));
   U22 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n44);
   U23 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n39);
   U24 : INV_X1 port map( A => Ci, ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_26 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_26;

architecture SYN_BEHAVIORAL of PG_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_25 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_25;

architecture SYN_BEHAVIORAL of PG_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_24 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_24;

architecture SYN_BEHAVIORAL of PG_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_23 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_23;

architecture SYN_BEHAVIORAL of PG_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_22 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_22;

architecture SYN_BEHAVIORAL of PG_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_21 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_21;

architecture SYN_BEHAVIORAL of PG_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_20 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_20;

architecture SYN_BEHAVIORAL of PG_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_19 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_19;

architecture SYN_BEHAVIORAL of PG_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_18 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_18;

architecture SYN_BEHAVIORAL of PG_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_17 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_17;

architecture SYN_BEHAVIORAL of PG_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_16 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_16;

architecture SYN_BEHAVIORAL of PG_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_15 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_15;

architecture SYN_BEHAVIORAL of PG_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_14 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_14;

architecture SYN_BEHAVIORAL of PG_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_13 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_13;

architecture SYN_BEHAVIORAL of PG_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_12 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_12;

architecture SYN_BEHAVIORAL of PG_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);
   U2 : INV_X1 port map( A => n4, ZN => G_ij);
   U3 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_11 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_11;

architecture SYN_BEHAVIORAL of PG_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_10 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_10;

architecture SYN_BEHAVIORAL of PG_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_9 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_9;

architecture SYN_BEHAVIORAL of PG_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_8 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_8;

architecture SYN_BEHAVIORAL of PG_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_7 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_7;

architecture SYN_BEHAVIORAL of PG_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_6 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_6;

architecture SYN_BEHAVIORAL of PG_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_5 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_5;

architecture SYN_BEHAVIORAL of PG_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);
   U2 : INV_X1 port map( A => n4, ZN => G_ij);
   U3 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_4 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_4;

architecture SYN_BEHAVIORAL of PG_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_3 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_3;

architecture SYN_BEHAVIORAL of PG_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_2 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_2;

architecture SYN_BEHAVIORAL of PG_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);
   U2 : INV_X1 port map( A => n4, ZN => G_ij);
   U3 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_1 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_1;

architecture SYN_BEHAVIORAL of PG_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);
   U2 : INV_X1 port map( A => n4, ZN => G_ij);
   U3 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_8 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_8;

architecture SYN_BEHAVIORAL of G_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_7 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_7;

architecture SYN_BEHAVIORAL of G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_6 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_6;

architecture SYN_BEHAVIORAL of G_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_5 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_5;

architecture SYN_BEHAVIORAL of G_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_4 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_4;

architecture SYN_BEHAVIORAL of G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_3 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_3;

architecture SYN_BEHAVIORAL of G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_2 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_2;

architecture SYN_BEHAVIORAL of G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_1 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_1;

architecture SYN_BEHAVIORAL of G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_31 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_31;

architecture SYN_BEHAVIORAL of pg_generator_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_30 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_30;

architecture SYN_BEHAVIORAL of pg_generator_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_29 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_29;

architecture SYN_BEHAVIORAL of pg_generator_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_28 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_28;

architecture SYN_BEHAVIORAL of pg_generator_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_27 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_27;

architecture SYN_BEHAVIORAL of pg_generator_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_26 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_26;

architecture SYN_BEHAVIORAL of pg_generator_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_25 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_25;

architecture SYN_BEHAVIORAL of pg_generator_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_24 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_24;

architecture SYN_BEHAVIORAL of pg_generator_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_23 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_23;

architecture SYN_BEHAVIORAL of pg_generator_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_22 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_22;

architecture SYN_BEHAVIORAL of pg_generator_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_21 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_21;

architecture SYN_BEHAVIORAL of pg_generator_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_20 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_20;

architecture SYN_BEHAVIORAL of pg_generator_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_19 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_19;

architecture SYN_BEHAVIORAL of pg_generator_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_18 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_18;

architecture SYN_BEHAVIORAL of pg_generator_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_17 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_17;

architecture SYN_BEHAVIORAL of pg_generator_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_16 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_16;

architecture SYN_BEHAVIORAL of pg_generator_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_15 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_15;

architecture SYN_BEHAVIORAL of pg_generator_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_14 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_14;

architecture SYN_BEHAVIORAL of pg_generator_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_13 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_13;

architecture SYN_BEHAVIORAL of pg_generator_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_12 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_12;

architecture SYN_BEHAVIORAL of pg_generator_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_11 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_11;

architecture SYN_BEHAVIORAL of pg_generator_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_10 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_10;

architecture SYN_BEHAVIORAL of pg_generator_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_9 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_9;

architecture SYN_BEHAVIORAL of pg_generator_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_8 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_8;

architecture SYN_BEHAVIORAL of pg_generator_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_7 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_7;

architecture SYN_BEHAVIORAL of pg_generator_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_6 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_6;

architecture SYN_BEHAVIORAL of pg_generator_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_5 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_5;

architecture SYN_BEHAVIORAL of pg_generator_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_4 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_4;

architecture SYN_BEHAVIORAL of pg_generator_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_3 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_3;

architecture SYN_BEHAVIORAL of pg_generator_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_2 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_2;

architecture SYN_BEHAVIORAL of pg_generator_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_1 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_1;

architecture SYN_BEHAVIORAL of pg_generator_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_6;

architecture SYN_STRUCTURAL of CarrySelect_6 is

   component MUX21_GENERIC_bits4_6
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1000, n_1001 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1000);
   RCA2 : RCA_NBITS4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1001);
   MUX21_GEN : MUX21_GENERIC_bits4_6 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_5;

architecture SYN_STRUCTURAL of CarrySelect_5 is

   component MUX21_GENERIC_bits4_5
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1002, n_1003 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1002);
   RCA2 : RCA_NBITS4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1003);
   MUX21_GEN : MUX21_GENERIC_bits4_5 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_4;

architecture SYN_STRUCTURAL of CarrySelect_4 is

   component MUX21_GENERIC_bits4_4
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1004, n_1005 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1004);
   RCA2 : RCA_NBITS4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1005);
   MUX21_GEN : MUX21_GENERIC_bits4_4 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_3;

architecture SYN_STRUCTURAL of CarrySelect_3 is

   component MUX21_GENERIC_bits4_3
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1006, n_1007 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1006);
   RCA2 : RCA_NBITS4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1007);
   MUX21_GEN : MUX21_GENERIC_bits4_3 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_2;

architecture SYN_STRUCTURAL of CarrySelect_2 is

   component MUX21_GENERIC_bits4_2
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1008, n_1009 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1008);
   RCA2 : RCA_NBITS4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1009);
   MUX21_GEN : MUX21_GENERIC_bits4_2 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_1;

architecture SYN_STRUCTURAL of CarrySelect_1 is

   component MUX21_GENERIC_bits4_1
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1010, n_1011 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1010);
   RCA2 : RCA_NBITS4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1011);
   MUX21_GEN : MUX21_GENERIC_bits4_1 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_351 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_351;

architecture SYN_ASYNCH_FD of FD_351 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_350 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_350;

architecture SYN_ASYNCH_FD of FD_350 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_349 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_349;

architecture SYN_ASYNCH_FD of FD_349 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_348 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_348;

architecture SYN_ASYNCH_FD of FD_348 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_347 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_347;

architecture SYN_ASYNCH_FD of FD_347 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_346 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_346;

architecture SYN_ASYNCH_FD of FD_346 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_345 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_345;

architecture SYN_ASYNCH_FD of FD_345 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_344 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_344;

architecture SYN_ASYNCH_FD of FD_344 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_343 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_343;

architecture SYN_ASYNCH_FD of FD_343 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_342 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_342;

architecture SYN_ASYNCH_FD of FD_342 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_341 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_341;

architecture SYN_ASYNCH_FD of FD_341 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_340 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_340;

architecture SYN_ASYNCH_FD of FD_340 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_339 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_339;

architecture SYN_ASYNCH_FD of FD_339 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_338 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_338;

architecture SYN_ASYNCH_FD of FD_338 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_337 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_337;

architecture SYN_ASYNCH_FD of FD_337 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_336 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_336;

architecture SYN_ASYNCH_FD of FD_336 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_335 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_335;

architecture SYN_ASYNCH_FD of FD_335 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_334 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_334;

architecture SYN_ASYNCH_FD of FD_334 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_333 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_333;

architecture SYN_ASYNCH_FD of FD_333 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_332 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_332;

architecture SYN_ASYNCH_FD of FD_332 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_331 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_331;

architecture SYN_ASYNCH_FD of FD_331 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_330 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_330;

architecture SYN_ASYNCH_FD of FD_330 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_329 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_329;

architecture SYN_ASYNCH_FD of FD_329 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_328 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_328;

architecture SYN_ASYNCH_FD of FD_328 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_327 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_327;

architecture SYN_ASYNCH_FD of FD_327 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_326 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_326;

architecture SYN_ASYNCH_FD of FD_326 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_325 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_325;

architecture SYN_ASYNCH_FD of FD_325 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_324 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_324;

architecture SYN_ASYNCH_FD of FD_324 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_323 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_323;

architecture SYN_ASYNCH_FD of FD_323 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_322 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_322;

architecture SYN_ASYNCH_FD of FD_322 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_321 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_321;

architecture SYN_ASYNCH_FD of FD_321 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6, n7 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n6);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OR2_X1 port map( A1 => n6, A2 => ENABLE, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n7, A2 => n5, ZN => n1);
   U5 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n7);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_320 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_320;

architecture SYN_ASYNCH_FD of FD_320 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_319 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_319;

architecture SYN_ASYNCH_FD of FD_319 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_318 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_318;

architecture SYN_ASYNCH_FD of FD_318 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_317 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_317;

architecture SYN_ASYNCH_FD of FD_317 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_316 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_316;

architecture SYN_ASYNCH_FD of FD_316 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_315 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_315;

architecture SYN_ASYNCH_FD of FD_315 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_314 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_314;

architecture SYN_ASYNCH_FD of FD_314 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_313 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_313;

architecture SYN_ASYNCH_FD of FD_313 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_312 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_312;

architecture SYN_ASYNCH_FD of FD_312 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_311 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_311;

architecture SYN_ASYNCH_FD of FD_311 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_310 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_310;

architecture SYN_ASYNCH_FD of FD_310 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_309 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_309;

architecture SYN_ASYNCH_FD of FD_309 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_308 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_308;

architecture SYN_ASYNCH_FD of FD_308 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_307 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_307;

architecture SYN_ASYNCH_FD of FD_307 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_306 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_306;

architecture SYN_ASYNCH_FD of FD_306 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_305 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_305;

architecture SYN_ASYNCH_FD of FD_305 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_304 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_304;

architecture SYN_ASYNCH_FD of FD_304 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_303 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_303;

architecture SYN_ASYNCH_FD of FD_303 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_302 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_302;

architecture SYN_ASYNCH_FD of FD_302 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_301 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_301;

architecture SYN_ASYNCH_FD of FD_301 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_300 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_300;

architecture SYN_ASYNCH_FD of FD_300 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_299 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_299;

architecture SYN_ASYNCH_FD of FD_299 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_298 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_298;

architecture SYN_ASYNCH_FD of FD_298 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_297 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_297;

architecture SYN_ASYNCH_FD of FD_297 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_296 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_296;

architecture SYN_ASYNCH_FD of FD_296 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_295 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_295;

architecture SYN_ASYNCH_FD of FD_295 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_294 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_294;

architecture SYN_ASYNCH_FD of FD_294 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_293 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_293;

architecture SYN_ASYNCH_FD of FD_293 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_292 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_292;

architecture SYN_ASYNCH_FD of FD_292 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_291 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_291;

architecture SYN_ASYNCH_FD of FD_291 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_290 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_290;

architecture SYN_ASYNCH_FD of FD_290 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_289 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_289;

architecture SYN_ASYNCH_FD of FD_289 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_288 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_288;

architecture SYN_ASYNCH_FD of FD_288 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_287 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_287;

architecture SYN_ASYNCH_FD of FD_287 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_286 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_286;

architecture SYN_ASYNCH_FD of FD_286 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_285 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_285;

architecture SYN_ASYNCH_FD of FD_285 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_284 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_284;

architecture SYN_ASYNCH_FD of FD_284 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_283 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_283;

architecture SYN_ASYNCH_FD of FD_283 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_282 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_282;

architecture SYN_ASYNCH_FD of FD_282 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_281 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_281;

architecture SYN_ASYNCH_FD of FD_281 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_280 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_280;

architecture SYN_ASYNCH_FD of FD_280 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_279 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_279;

architecture SYN_ASYNCH_FD of FD_279 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_278 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_278;

architecture SYN_ASYNCH_FD of FD_278 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_277 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_277;

architecture SYN_ASYNCH_FD of FD_277 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_276 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_276;

architecture SYN_ASYNCH_FD of FD_276 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_275 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_275;

architecture SYN_ASYNCH_FD of FD_275 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_274 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_274;

architecture SYN_ASYNCH_FD of FD_274 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_273 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_273;

architecture SYN_ASYNCH_FD of FD_273 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_272 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_272;

architecture SYN_ASYNCH_FD of FD_272 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_271 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_271;

architecture SYN_ASYNCH_FD of FD_271 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_270 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_270;

architecture SYN_ASYNCH_FD of FD_270 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_269 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_269;

architecture SYN_ASYNCH_FD of FD_269 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_268 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_268;

architecture SYN_ASYNCH_FD of FD_268 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_267 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_267;

architecture SYN_ASYNCH_FD of FD_267 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_266 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_266;

architecture SYN_ASYNCH_FD of FD_266 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_265 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_265;

architecture SYN_ASYNCH_FD of FD_265 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_264 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_264;

architecture SYN_ASYNCH_FD of FD_264 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_263 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_263;

architecture SYN_ASYNCH_FD of FD_263 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_262 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_262;

architecture SYN_ASYNCH_FD of FD_262 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_261 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_261;

architecture SYN_ASYNCH_FD of FD_261 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_260 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_260;

architecture SYN_ASYNCH_FD of FD_260 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_259 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_259;

architecture SYN_ASYNCH_FD of FD_259 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_258 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_258;

architecture SYN_ASYNCH_FD of FD_258 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_257 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_257;

architecture SYN_ASYNCH_FD of FD_257 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_256 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_256;

architecture SYN_ASYNCH_FD of FD_256 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_255 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_255;

architecture SYN_ASYNCH_FD of FD_255 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_254 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_254;

architecture SYN_ASYNCH_FD of FD_254 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_253 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_253;

architecture SYN_ASYNCH_FD of FD_253 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_252 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_252;

architecture SYN_ASYNCH_FD of FD_252 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_251 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_251;

architecture SYN_ASYNCH_FD of FD_251 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_250 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_250;

architecture SYN_ASYNCH_FD of FD_250 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_249 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_249;

architecture SYN_ASYNCH_FD of FD_249 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_248 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_248;

architecture SYN_ASYNCH_FD of FD_248 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_247 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_247;

architecture SYN_ASYNCH_FD of FD_247 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_246 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_246;

architecture SYN_ASYNCH_FD of FD_246 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_245 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_245;

architecture SYN_ASYNCH_FD of FD_245 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_244 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_244;

architecture SYN_ASYNCH_FD of FD_244 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_243 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_243;

architecture SYN_ASYNCH_FD of FD_243 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_242 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_242;

architecture SYN_ASYNCH_FD of FD_242 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_241 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_241;

architecture SYN_ASYNCH_FD of FD_241 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_240 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_240;

architecture SYN_ASYNCH_FD of FD_240 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_239 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_239;

architecture SYN_ASYNCH_FD of FD_239 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_238 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_238;

architecture SYN_ASYNCH_FD of FD_238 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_237 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_237;

architecture SYN_ASYNCH_FD of FD_237 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_236 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_236;

architecture SYN_ASYNCH_FD of FD_236 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_235 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_235;

architecture SYN_ASYNCH_FD of FD_235 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_234 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_234;

architecture SYN_ASYNCH_FD of FD_234 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_233 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_233;

architecture SYN_ASYNCH_FD of FD_233 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_232 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_232;

architecture SYN_ASYNCH_FD of FD_232 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_231 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_231;

architecture SYN_ASYNCH_FD of FD_231 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_230 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_230;

architecture SYN_ASYNCH_FD of FD_230 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_229 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_229;

architecture SYN_ASYNCH_FD of FD_229 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_228 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_228;

architecture SYN_ASYNCH_FD of FD_228 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_227 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_227;

architecture SYN_ASYNCH_FD of FD_227 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_226 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_226;

architecture SYN_ASYNCH_FD of FD_226 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_225 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_225;

architecture SYN_ASYNCH_FD of FD_225 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_224 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_224;

architecture SYN_ASYNCH_FD of FD_224 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_223 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_223;

architecture SYN_ASYNCH_FD of FD_223 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_222 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_222;

architecture SYN_ASYNCH_FD of FD_222 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_221 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_221;

architecture SYN_ASYNCH_FD of FD_221 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_220 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_220;

architecture SYN_ASYNCH_FD of FD_220 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_219 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_219;

architecture SYN_ASYNCH_FD of FD_219 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_218 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_218;

architecture SYN_ASYNCH_FD of FD_218 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_217 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_217;

architecture SYN_ASYNCH_FD of FD_217 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_216 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_216;

architecture SYN_ASYNCH_FD of FD_216 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_215 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_215;

architecture SYN_ASYNCH_FD of FD_215 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_214 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_214;

architecture SYN_ASYNCH_FD of FD_214 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_213 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_213;

architecture SYN_ASYNCH_FD of FD_213 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_212 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_212;

architecture SYN_ASYNCH_FD of FD_212 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_211 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_211;

architecture SYN_ASYNCH_FD of FD_211 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_210 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_210;

architecture SYN_ASYNCH_FD of FD_210 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_209 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_209;

architecture SYN_ASYNCH_FD of FD_209 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_208 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_208;

architecture SYN_ASYNCH_FD of FD_208 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_207 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_207;

architecture SYN_ASYNCH_FD of FD_207 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_206 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_206;

architecture SYN_ASYNCH_FD of FD_206 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_205 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_205;

architecture SYN_ASYNCH_FD of FD_205 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_204 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_204;

architecture SYN_ASYNCH_FD of FD_204 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_203 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_203;

architecture SYN_ASYNCH_FD of FD_203 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_202 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_202;

architecture SYN_ASYNCH_FD of FD_202 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_201 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_201;

architecture SYN_ASYNCH_FD of FD_201 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_200 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_200;

architecture SYN_ASYNCH_FD of FD_200 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_199 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_199;

architecture SYN_ASYNCH_FD of FD_199 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_198 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_198;

architecture SYN_ASYNCH_FD of FD_198 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_197 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_197;

architecture SYN_ASYNCH_FD of FD_197 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_196 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_196;

architecture SYN_ASYNCH_FD of FD_196 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_195 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_195;

architecture SYN_ASYNCH_FD of FD_195 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_194 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_194;

architecture SYN_ASYNCH_FD of FD_194 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_193 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_193;

architecture SYN_ASYNCH_FD of FD_193 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_192 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_192;

architecture SYN_ASYNCH_FD of FD_192 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_191 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_191;

architecture SYN_ASYNCH_FD of FD_191 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_190 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_190;

architecture SYN_ASYNCH_FD of FD_190 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_189 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_189;

architecture SYN_ASYNCH_FD of FD_189 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_188 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_188;

architecture SYN_ASYNCH_FD of FD_188 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_187 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_187;

architecture SYN_ASYNCH_FD of FD_187 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_186 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_186;

architecture SYN_ASYNCH_FD of FD_186 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_185 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_185;

architecture SYN_ASYNCH_FD of FD_185 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_184 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_184;

architecture SYN_ASYNCH_FD of FD_184 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_183 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_183;

architecture SYN_ASYNCH_FD of FD_183 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_182 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_182;

architecture SYN_ASYNCH_FD of FD_182 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_181 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_181;

architecture SYN_ASYNCH_FD of FD_181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_180 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_180;

architecture SYN_ASYNCH_FD of FD_180 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_179 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_179;

architecture SYN_ASYNCH_FD of FD_179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_178 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_178;

architecture SYN_ASYNCH_FD of FD_178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_177 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_177;

architecture SYN_ASYNCH_FD of FD_177 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_176 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_176;

architecture SYN_ASYNCH_FD of FD_176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_175 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_175;

architecture SYN_ASYNCH_FD of FD_175 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_174 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_174;

architecture SYN_ASYNCH_FD of FD_174 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_173 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_173;

architecture SYN_ASYNCH_FD of FD_173 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_172 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_172;

architecture SYN_ASYNCH_FD of FD_172 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_171 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_171;

architecture SYN_ASYNCH_FD of FD_171 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_170 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_170;

architecture SYN_ASYNCH_FD of FD_170 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_169 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_169;

architecture SYN_ASYNCH_FD of FD_169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_168 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_168;

architecture SYN_ASYNCH_FD of FD_168 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_167 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_167;

architecture SYN_ASYNCH_FD of FD_167 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_166 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_166;

architecture SYN_ASYNCH_FD of FD_166 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_165 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_165;

architecture SYN_ASYNCH_FD of FD_165 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_164 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_164;

architecture SYN_ASYNCH_FD of FD_164 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_163 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_163;

architecture SYN_ASYNCH_FD of FD_163 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_162 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_162;

architecture SYN_ASYNCH_FD of FD_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_161 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_161;

architecture SYN_ASYNCH_FD of FD_161 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_160 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_160;

architecture SYN_ASYNCH_FD of FD_160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_159 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_159;

architecture SYN_ASYNCH_FD of FD_159 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_158 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_158;

architecture SYN_ASYNCH_FD of FD_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_157 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_157;

architecture SYN_ASYNCH_FD of FD_157 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_156 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_156;

architecture SYN_ASYNCH_FD of FD_156 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_155 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_155;

architecture SYN_ASYNCH_FD of FD_155 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_154 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_154;

architecture SYN_ASYNCH_FD of FD_154 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_153 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_153;

architecture SYN_ASYNCH_FD of FD_153 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_152 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_152;

architecture SYN_ASYNCH_FD of FD_152 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_151 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_151;

architecture SYN_ASYNCH_FD of FD_151 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_150 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_150;

architecture SYN_ASYNCH_FD of FD_150 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_149 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_149;

architecture SYN_ASYNCH_FD of FD_149 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_148 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_148;

architecture SYN_ASYNCH_FD of FD_148 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_147 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_147;

architecture SYN_ASYNCH_FD of FD_147 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_146 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_146;

architecture SYN_ASYNCH_FD of FD_146 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_145 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_145;

architecture SYN_ASYNCH_FD of FD_145 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_144 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_144;

architecture SYN_ASYNCH_FD of FD_144 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_143 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_143;

architecture SYN_ASYNCH_FD of FD_143 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_142 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_142;

architecture SYN_ASYNCH_FD of FD_142 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_141 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_141;

architecture SYN_ASYNCH_FD of FD_141 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_140 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_140;

architecture SYN_ASYNCH_FD of FD_140 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_139 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_139;

architecture SYN_ASYNCH_FD of FD_139 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_138 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_138;

architecture SYN_ASYNCH_FD of FD_138 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_137 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_137;

architecture SYN_ASYNCH_FD of FD_137 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_136 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_136;

architecture SYN_ASYNCH_FD of FD_136 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_135 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_135;

architecture SYN_ASYNCH_FD of FD_135 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_134 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_134;

architecture SYN_ASYNCH_FD of FD_134 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_133 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_133;

architecture SYN_ASYNCH_FD of FD_133 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_132 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_132;

architecture SYN_ASYNCH_FD of FD_132 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_131 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_131;

architecture SYN_ASYNCH_FD of FD_131 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_130 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_130;

architecture SYN_ASYNCH_FD of FD_130 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_129 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_129;

architecture SYN_ASYNCH_FD of FD_129 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U4 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_128 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_128;

architecture SYN_ASYNCH_FD of FD_128 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_127 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_127;

architecture SYN_ASYNCH_FD of FD_127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_126 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_126;

architecture SYN_ASYNCH_FD of FD_126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_125 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_125;

architecture SYN_ASYNCH_FD of FD_125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_124 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_124;

architecture SYN_ASYNCH_FD of FD_124 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_123 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_123;

architecture SYN_ASYNCH_FD of FD_123 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_122 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_122;

architecture SYN_ASYNCH_FD of FD_122 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_121 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_121;

architecture SYN_ASYNCH_FD of FD_121 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_120 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_120;

architecture SYN_ASYNCH_FD of FD_120 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_119 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_119;

architecture SYN_ASYNCH_FD of FD_119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_118 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_118;

architecture SYN_ASYNCH_FD of FD_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_117 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_117;

architecture SYN_ASYNCH_FD of FD_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_116 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_116;

architecture SYN_ASYNCH_FD of FD_116 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_115 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_115;

architecture SYN_ASYNCH_FD of FD_115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_114 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_114;

architecture SYN_ASYNCH_FD of FD_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_113 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_113;

architecture SYN_ASYNCH_FD of FD_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_112 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_112;

architecture SYN_ASYNCH_FD of FD_112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_111 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_111;

architecture SYN_ASYNCH_FD of FD_111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_110 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_110;

architecture SYN_ASYNCH_FD of FD_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_109 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_109;

architecture SYN_ASYNCH_FD of FD_109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_108 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_108;

architecture SYN_ASYNCH_FD of FD_108 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_107 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_107;

architecture SYN_ASYNCH_FD of FD_107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_106 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_106;

architecture SYN_ASYNCH_FD of FD_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_105 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_105;

architecture SYN_ASYNCH_FD of FD_105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_104 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_104;

architecture SYN_ASYNCH_FD of FD_104 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_103 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_103;

architecture SYN_ASYNCH_FD of FD_103 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_102 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_102;

architecture SYN_ASYNCH_FD of FD_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_101 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_101;

architecture SYN_ASYNCH_FD of FD_101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_100 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_100;

architecture SYN_ASYNCH_FD of FD_100 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_99 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_99;

architecture SYN_ASYNCH_FD of FD_99 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_98 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_98;

architecture SYN_ASYNCH_FD of FD_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_97 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_97;

architecture SYN_ASYNCH_FD of FD_97 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_96 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_96;

architecture SYN_ASYNCH_FD of FD_96 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_95 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_95;

architecture SYN_ASYNCH_FD of FD_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_94 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_94;

architecture SYN_ASYNCH_FD of FD_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_93 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_93;

architecture SYN_ASYNCH_FD of FD_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_92 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_92;

architecture SYN_ASYNCH_FD of FD_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_91 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_91;

architecture SYN_ASYNCH_FD of FD_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_90 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_90;

architecture SYN_ASYNCH_FD of FD_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_89 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_89;

architecture SYN_ASYNCH_FD of FD_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_88 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_88;

architecture SYN_ASYNCH_FD of FD_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_87 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_87;

architecture SYN_ASYNCH_FD of FD_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_86 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_86;

architecture SYN_ASYNCH_FD of FD_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_85 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_85;

architecture SYN_ASYNCH_FD of FD_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_84 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_84;

architecture SYN_ASYNCH_FD of FD_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_83 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_83;

architecture SYN_ASYNCH_FD of FD_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_82 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_82;

architecture SYN_ASYNCH_FD of FD_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_81 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_81;

architecture SYN_ASYNCH_FD of FD_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_80 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_80;

architecture SYN_ASYNCH_FD of FD_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_79 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_79;

architecture SYN_ASYNCH_FD of FD_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_78 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_78;

architecture SYN_ASYNCH_FD of FD_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_77 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_77;

architecture SYN_ASYNCH_FD of FD_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_76 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_76;

architecture SYN_ASYNCH_FD of FD_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_75 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_75;

architecture SYN_ASYNCH_FD of FD_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_74 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_74;

architecture SYN_ASYNCH_FD of FD_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_73 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_73;

architecture SYN_ASYNCH_FD of FD_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_72 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_72;

architecture SYN_ASYNCH_FD of FD_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_71 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_71;

architecture SYN_ASYNCH_FD of FD_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_70 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_70;

architecture SYN_ASYNCH_FD of FD_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_69 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_69;

architecture SYN_ASYNCH_FD of FD_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_68 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_68;

architecture SYN_ASYNCH_FD of FD_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_67 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_67;

architecture SYN_ASYNCH_FD of FD_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_66 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_66;

architecture SYN_ASYNCH_FD of FD_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_65 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_65;

architecture SYN_ASYNCH_FD of FD_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_64 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_64;

architecture SYN_ASYNCH_FD of FD_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_63 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_63;

architecture SYN_ASYNCH_FD of FD_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_62 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_62;

architecture SYN_ASYNCH_FD of FD_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_61 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_61;

architecture SYN_ASYNCH_FD of FD_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_60 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_60;

architecture SYN_ASYNCH_FD of FD_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_59 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_59;

architecture SYN_ASYNCH_FD of FD_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_58 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_58;

architecture SYN_ASYNCH_FD of FD_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_57 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_57;

architecture SYN_ASYNCH_FD of FD_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_56 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_56;

architecture SYN_ASYNCH_FD of FD_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_55 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_55;

architecture SYN_ASYNCH_FD of FD_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_54 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_54;

architecture SYN_ASYNCH_FD of FD_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_53 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_53;

architecture SYN_ASYNCH_FD of FD_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_52 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_52;

architecture SYN_ASYNCH_FD of FD_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_51 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_51;

architecture SYN_ASYNCH_FD of FD_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_50 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_50;

architecture SYN_ASYNCH_FD of FD_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_49 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_49;

architecture SYN_ASYNCH_FD of FD_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_48 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_48;

architecture SYN_ASYNCH_FD of FD_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_47 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_47;

architecture SYN_ASYNCH_FD of FD_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_46 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_46;

architecture SYN_ASYNCH_FD of FD_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_45 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_45;

architecture SYN_ASYNCH_FD of FD_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_44 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_44;

architecture SYN_ASYNCH_FD of FD_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_43 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_43;

architecture SYN_ASYNCH_FD of FD_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_42 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_42;

architecture SYN_ASYNCH_FD of FD_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_41 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_41;

architecture SYN_ASYNCH_FD of FD_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_40 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_40;

architecture SYN_ASYNCH_FD of FD_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_39 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_39;

architecture SYN_ASYNCH_FD of FD_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_38 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_38;

architecture SYN_ASYNCH_FD of FD_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_37 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_37;

architecture SYN_ASYNCH_FD of FD_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_36 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_36;

architecture SYN_ASYNCH_FD of FD_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_35 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_35;

architecture SYN_ASYNCH_FD of FD_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_34 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_34;

architecture SYN_ASYNCH_FD of FD_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_33 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_33;

architecture SYN_ASYNCH_FD of FD_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_32 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_32;

architecture SYN_ASYNCH_FD of FD_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_31 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_31;

architecture SYN_ASYNCH_FD of FD_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_30 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_30;

architecture SYN_ASYNCH_FD of FD_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_29 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_29;

architecture SYN_ASYNCH_FD of FD_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_28 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_28;

architecture SYN_ASYNCH_FD of FD_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_27 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_27;

architecture SYN_ASYNCH_FD of FD_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_26 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_26;

architecture SYN_ASYNCH_FD of FD_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_25 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_25;

architecture SYN_ASYNCH_FD of FD_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_24 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_24;

architecture SYN_ASYNCH_FD of FD_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_23 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_23;

architecture SYN_ASYNCH_FD of FD_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_22 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_22;

architecture SYN_ASYNCH_FD of FD_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_21 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_21;

architecture SYN_ASYNCH_FD of FD_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_20 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_20;

architecture SYN_ASYNCH_FD of FD_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_19 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_19;

architecture SYN_ASYNCH_FD of FD_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_18 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_18;

architecture SYN_ASYNCH_FD of FD_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_17 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_17;

architecture SYN_ASYNCH_FD of FD_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_16 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_16;

architecture SYN_ASYNCH_FD of FD_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_15 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_15;

architecture SYN_ASYNCH_FD of FD_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_14 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_14;

architecture SYN_ASYNCH_FD of FD_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_13 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_13;

architecture SYN_ASYNCH_FD of FD_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_12 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_12;

architecture SYN_ASYNCH_FD of FD_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_11 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_11;

architecture SYN_ASYNCH_FD of FD_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_10 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_10;

architecture SYN_ASYNCH_FD of FD_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_9 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_9;

architecture SYN_ASYNCH_FD of FD_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_8 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_8;

architecture SYN_ASYNCH_FD of FD_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_7 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_7;

architecture SYN_ASYNCH_FD of FD_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_6 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_6;

architecture SYN_ASYNCH_FD of FD_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_5 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_5;

architecture SYN_ASYNCH_FD of FD_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_4 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_4;

architecture SYN_ASYNCH_FD of FD_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_3 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_3;

architecture SYN_ASYNCH_FD of FD_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_2 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_2;

architecture SYN_ASYNCH_FD of FD_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_1 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_1;

architecture SYN_ASYNCH_FD of FD_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => ENABLE, A => n6, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n6);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_3;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n33, n66, n67, n68, n69, n70, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n70, Z => n69);
   U2 : INV_X1 port map( A => S, ZN => n70);
   U3 : INV_X1 port map( A => n70, ZN => n68);
   U4 : BUF_X1 port map( A => n69, Z => n33);
   U5 : BUF_X1 port map( A => n69, Z => n67);
   U6 : BUF_X1 port map( A => n69, Z => n66);
   U7 : INV_X1 port map( A => n103, ZN => Y(0));
   U8 : AOI22_X1 port map( A1 => A(0), A2 => n68, B1 => B(0), B2 => n33, ZN => 
                           n103);
   U9 : INV_X1 port map( A => n128, ZN => Y(3));
   U10 : AOI22_X1 port map( A1 => A(3), A2 => n68, B1 => B(3), B2 => n67, ZN =>
                           n128);
   U11 : INV_X1 port map( A => n114, ZN => Y(1));
   U12 : AOI22_X1 port map( A1 => A(1), A2 => n68, B1 => B(1), B2 => n33, ZN =>
                           n114);
   U13 : INV_X1 port map( A => n125, ZN => Y(2));
   U14 : AOI22_X1 port map( A1 => A(2), A2 => S, B1 => B(2), B2 => n66, ZN => 
                           n125);
   U15 : INV_X1 port map( A => n130, ZN => Y(5));
   U16 : AOI22_X1 port map( A1 => A(5), A2 => S, B1 => B(5), B2 => n67, ZN => 
                           n130);
   U17 : INV_X1 port map( A => n132, ZN => Y(7));
   U18 : AOI22_X1 port map( A1 => A(7), A2 => n68, B1 => B(7), B2 => n67, ZN =>
                           n132);
   U19 : INV_X1 port map( A => n129, ZN => Y(4));
   U20 : AOI22_X1 port map( A1 => A(4), A2 => n68, B1 => B(4), B2 => n67, ZN =>
                           n129);
   U21 : INV_X1 port map( A => n131, ZN => Y(6));
   U22 : AOI22_X1 port map( A1 => A(6), A2 => n68, B1 => B(6), B2 => n67, ZN =>
                           n131);
   U23 : INV_X1 port map( A => n134, ZN => Y(9));
   U24 : AOI22_X1 port map( A1 => S, A2 => A(9), B1 => B(9), B2 => n67, ZN => 
                           n134);
   U25 : INV_X1 port map( A => n105, ZN => Y(11));
   U26 : AOI22_X1 port map( A1 => A(11), A2 => n68, B1 => B(11), B2 => n33, ZN 
                           => n105);
   U27 : INV_X1 port map( A => n107, ZN => Y(13));
   U28 : AOI22_X1 port map( A1 => A(13), A2 => n68, B1 => B(13), B2 => n33, ZN 
                           => n107);
   U29 : INV_X1 port map( A => n123, ZN => Y(28));
   U30 : AOI22_X1 port map( A1 => A(28), A2 => n68, B1 => B(28), B2 => n66, ZN 
                           => n123);
   U31 : INV_X1 port map( A => n109, ZN => Y(15));
   U32 : AOI22_X1 port map( A1 => A(15), A2 => n68, B1 => B(15), B2 => n33, ZN 
                           => n109);
   U33 : INV_X1 port map( A => n133, ZN => Y(8));
   U34 : AOI22_X1 port map( A1 => A(8), A2 => S, B1 => B(8), B2 => n67, ZN => 
                           n133);
   U35 : INV_X1 port map( A => n110, ZN => Y(16));
   U36 : AOI22_X1 port map( A1 => A(16), A2 => n68, B1 => B(16), B2 => n33, ZN 
                           => n110);
   U37 : INV_X1 port map( A => n106, ZN => Y(12));
   U38 : AOI22_X1 port map( A1 => A(12), A2 => n68, B1 => B(12), B2 => n33, ZN 
                           => n106);
   U39 : INV_X1 port map( A => n104, ZN => Y(10));
   U40 : AOI22_X1 port map( A1 => A(10), A2 => n68, B1 => B(10), B2 => n33, ZN 
                           => n104);
   U41 : INV_X1 port map( A => n115, ZN => Y(20));
   U42 : AOI22_X1 port map( A1 => A(20), A2 => S, B1 => B(20), B2 => n66, ZN =>
                           n115);
   U43 : INV_X1 port map( A => n108, ZN => Y(14));
   U44 : AOI22_X1 port map( A1 => A(14), A2 => n68, B1 => B(14), B2 => n33, ZN 
                           => n108);
   U45 : INV_X1 port map( A => n111, ZN => Y(17));
   U46 : AOI22_X1 port map( A1 => A(17), A2 => n68, B1 => B(17), B2 => n33, ZN 
                           => n111);
   U47 : INV_X1 port map( A => n113, ZN => Y(19));
   U48 : AOI22_X1 port map( A1 => A(19), A2 => n68, B1 => B(19), B2 => n33, ZN 
                           => n113);
   U49 : INV_X1 port map( A => n119, ZN => Y(24));
   U50 : AOI22_X1 port map( A1 => A(24), A2 => S, B1 => B(24), B2 => n66, ZN =>
                           n119);
   U51 : INV_X1 port map( A => n116, ZN => Y(21));
   U52 : AOI22_X1 port map( A1 => A(21), A2 => S, B1 => B(21), B2 => n66, ZN =>
                           n116);
   U53 : INV_X1 port map( A => n118, ZN => Y(23));
   U54 : AOI22_X1 port map( A1 => A(23), A2 => S, B1 => B(23), B2 => n66, ZN =>
                           n118);
   U55 : INV_X1 port map( A => n112, ZN => Y(18));
   U56 : AOI22_X1 port map( A1 => A(18), A2 => n68, B1 => B(18), B2 => n33, ZN 
                           => n112);
   U57 : INV_X1 port map( A => n117, ZN => Y(22));
   U58 : AOI22_X1 port map( A1 => A(22), A2 => S, B1 => B(22), B2 => n66, ZN =>
                           n117);
   U59 : INV_X1 port map( A => n124, ZN => Y(29));
   U60 : AOI22_X1 port map( A1 => A(29), A2 => S, B1 => B(29), B2 => n66, ZN =>
                           n124);
   U61 : INV_X1 port map( A => n120, ZN => Y(25));
   U62 : AOI22_X1 port map( A1 => A(25), A2 => S, B1 => B(25), B2 => n66, ZN =>
                           n120);
   U63 : INV_X1 port map( A => n122, ZN => Y(27));
   U64 : AOI22_X1 port map( A1 => A(27), A2 => S, B1 => B(27), B2 => n66, ZN =>
                           n122);
   U65 : INV_X1 port map( A => n121, ZN => Y(26));
   U66 : AOI22_X1 port map( A1 => A(26), A2 => S, B1 => B(26), B2 => n66, ZN =>
                           n121);
   U67 : INV_X1 port map( A => n126, ZN => Y(30));
   U68 : AOI22_X1 port map( A1 => A(30), A2 => S, B1 => B(30), B2 => n66, ZN =>
                           n126);
   U69 : INV_X1 port map( A => n127, ZN => Y(31));
   U70 : AOI22_X1 port map( A1 => A(31), A2 => n68, B1 => B(31), B2 => n67, ZN 
                           => n127);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_1;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n33, n66, n67, n68, n69, n70, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n70, Z => n69);
   U2 : INV_X1 port map( A => n70, ZN => n68);
   U3 : BUF_X1 port map( A => n69, Z => n67);
   U4 : BUF_X1 port map( A => n69, Z => n33);
   U5 : BUF_X1 port map( A => n69, Z => n66);
   U6 : INV_X1 port map( A => n128, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n68, B1 => B(3), B2 => n67, ZN => 
                           n128);
   U8 : INV_X1 port map( A => n129, ZN => Y(4));
   U9 : AOI22_X1 port map( A1 => A(4), A2 => n68, B1 => B(4), B2 => n67, ZN => 
                           n129);
   U10 : INV_X1 port map( A => n130, ZN => Y(5));
   U11 : AOI22_X1 port map( A1 => A(5), A2 => n68, B1 => B(5), B2 => n67, ZN =>
                           n130);
   U12 : INV_X1 port map( A => n131, ZN => Y(6));
   U13 : AOI22_X1 port map( A1 => A(6), A2 => n68, B1 => B(6), B2 => n67, ZN =>
                           n131);
   U14 : INV_X1 port map( A => n132, ZN => Y(7));
   U15 : AOI22_X1 port map( A1 => A(7), A2 => n68, B1 => B(7), B2 => n67, ZN =>
                           n132);
   U16 : INV_X1 port map( A => n133, ZN => Y(8));
   U17 : AOI22_X1 port map( A1 => A(8), A2 => n68, B1 => B(8), B2 => n67, ZN =>
                           n133);
   U18 : INV_X1 port map( A => n127, ZN => Y(31));
   U19 : AOI22_X1 port map( A1 => A(31), A2 => S, B1 => B(31), B2 => n67, ZN =>
                           n127);
   U20 : INV_X1 port map( A => S, ZN => n70);
   U21 : INV_X1 port map( A => n103, ZN => Y(0));
   U22 : AOI22_X1 port map( A1 => A(0), A2 => S, B1 => B(0), B2 => n33, ZN => 
                           n103);
   U23 : INV_X1 port map( A => n114, ZN => Y(1));
   U24 : AOI22_X1 port map( A1 => A(1), A2 => S, B1 => B(1), B2 => n33, ZN => 
                           n114);
   U25 : INV_X1 port map( A => n125, ZN => Y(2));
   U26 : AOI22_X1 port map( A1 => A(2), A2 => n68, B1 => B(2), B2 => n66, ZN =>
                           n125);
   U27 : INV_X1 port map( A => n104, ZN => Y(10));
   U28 : AOI22_X1 port map( A1 => A(10), A2 => S, B1 => B(10), B2 => n33, ZN =>
                           n104);
   U29 : INV_X1 port map( A => n105, ZN => Y(11));
   U30 : AOI22_X1 port map( A1 => A(11), A2 => S, B1 => B(11), B2 => n33, ZN =>
                           n105);
   U31 : INV_X1 port map( A => n106, ZN => Y(12));
   U32 : AOI22_X1 port map( A1 => A(12), A2 => S, B1 => B(12), B2 => n33, ZN =>
                           n106);
   U33 : INV_X1 port map( A => n107, ZN => Y(13));
   U34 : AOI22_X1 port map( A1 => A(13), A2 => S, B1 => B(13), B2 => n33, ZN =>
                           n107);
   U35 : INV_X1 port map( A => n108, ZN => Y(14));
   U36 : AOI22_X1 port map( A1 => A(14), A2 => S, B1 => B(14), B2 => n33, ZN =>
                           n108);
   U37 : INV_X1 port map( A => n109, ZN => Y(15));
   U38 : AOI22_X1 port map( A1 => A(15), A2 => S, B1 => B(15), B2 => n33, ZN =>
                           n109);
   U39 : INV_X1 port map( A => n110, ZN => Y(16));
   U40 : AOI22_X1 port map( A1 => A(16), A2 => S, B1 => B(16), B2 => n33, ZN =>
                           n110);
   U41 : INV_X1 port map( A => n111, ZN => Y(17));
   U42 : AOI22_X1 port map( A1 => A(17), A2 => S, B1 => B(17), B2 => n33, ZN =>
                           n111);
   U43 : INV_X1 port map( A => n112, ZN => Y(18));
   U44 : AOI22_X1 port map( A1 => A(18), A2 => S, B1 => B(18), B2 => n33, ZN =>
                           n112);
   U45 : INV_X1 port map( A => n113, ZN => Y(19));
   U46 : AOI22_X1 port map( A1 => A(19), A2 => S, B1 => B(19), B2 => n33, ZN =>
                           n113);
   U47 : INV_X1 port map( A => n115, ZN => Y(20));
   U48 : AOI22_X1 port map( A1 => A(20), A2 => n68, B1 => B(20), B2 => n66, ZN 
                           => n115);
   U49 : INV_X1 port map( A => n116, ZN => Y(21));
   U50 : AOI22_X1 port map( A1 => A(21), A2 => n68, B1 => B(21), B2 => n66, ZN 
                           => n116);
   U51 : INV_X1 port map( A => n117, ZN => Y(22));
   U52 : AOI22_X1 port map( A1 => A(22), A2 => n68, B1 => B(22), B2 => n66, ZN 
                           => n117);
   U53 : INV_X1 port map( A => n118, ZN => Y(23));
   U54 : AOI22_X1 port map( A1 => A(23), A2 => n68, B1 => B(23), B2 => n66, ZN 
                           => n118);
   U55 : INV_X1 port map( A => n119, ZN => Y(24));
   U56 : AOI22_X1 port map( A1 => A(24), A2 => n68, B1 => B(24), B2 => n66, ZN 
                           => n119);
   U57 : INV_X1 port map( A => n120, ZN => Y(25));
   U58 : AOI22_X1 port map( A1 => A(25), A2 => n68, B1 => B(25), B2 => n66, ZN 
                           => n120);
   U59 : INV_X1 port map( A => n121, ZN => Y(26));
   U60 : AOI22_X1 port map( A1 => A(26), A2 => n68, B1 => B(26), B2 => n66, ZN 
                           => n121);
   U61 : INV_X1 port map( A => n122, ZN => Y(27));
   U62 : AOI22_X1 port map( A1 => A(27), A2 => n68, B1 => B(27), B2 => n66, ZN 
                           => n122);
   U63 : INV_X1 port map( A => n123, ZN => Y(28));
   U64 : AOI22_X1 port map( A1 => A(28), A2 => n68, B1 => B(28), B2 => n66, ZN 
                           => n123);
   U65 : INV_X1 port map( A => n124, ZN => Y(29));
   U66 : AOI22_X1 port map( A1 => A(29), A2 => n68, B1 => B(29), B2 => n66, ZN 
                           => n124);
   U67 : INV_X1 port map( A => n126, ZN => Y(30));
   U68 : AOI22_X1 port map( A1 => A(30), A2 => n68, B1 => B(30), B2 => n66, ZN 
                           => n126);
   U69 : INV_X1 port map( A => n134, ZN => Y(9));
   U70 : AOI22_X1 port map( A1 => n68, A2 => A(9), B1 => B(9), B2 => n67, ZN =>
                           n134);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_7 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_7;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_7 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_193
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_194
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_195
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_196
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_197
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_198
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_199
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_200
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_201
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_202
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_203
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_204
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_205
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_206
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_207
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_208
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_209
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_210
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_211
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_212
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_213
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_214
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_215
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_216
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_217
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_218
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_219
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_220
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_221
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_222
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_223
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_224
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_224 port map( D => data_in(0), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(0));
   FF_1 : FD_223 port map( D => data_in(1), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(1));
   FF_2 : FD_222 port map( D => data_in(2), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(2));
   FF_3 : FD_221 port map( D => data_in(3), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(3));
   FF_4 : FD_220 port map( D => data_in(4), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(4));
   FF_5 : FD_219 port map( D => data_in(5), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(5));
   FF_6 : FD_218 port map( D => data_in(6), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(6));
   FF_7 : FD_217 port map( D => data_in(7), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(7));
   FF_8 : FD_216 port map( D => data_in(8), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(8));
   FF_9 : FD_215 port map( D => data_in(9), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(9));
   FF_10 : FD_214 port map( D => data_in(10), CK => CK, RESET => n13, ENABLE =>
                           n9, Q => data_out(10));
   FF_11 : FD_213 port map( D => data_in(11), CK => CK, RESET => n13, ENABLE =>
                           n9, Q => data_out(11));
   FF_12 : FD_212 port map( D => data_in(12), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(12));
   FF_13 : FD_211 port map( D => data_in(13), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(13));
   FF_14 : FD_210 port map( D => data_in(14), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(14));
   FF_15 : FD_209 port map( D => data_in(15), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(15));
   FF_16 : FD_208 port map( D => data_in(16), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(16));
   FF_17 : FD_207 port map( D => data_in(17), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(17));
   FF_18 : FD_206 port map( D => data_in(18), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(18));
   FF_19 : FD_205 port map( D => data_in(19), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(19));
   FF_20 : FD_204 port map( D => data_in(20), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(20));
   FF_21 : FD_203 port map( D => data_in(21), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(21));
   FF_22 : FD_202 port map( D => data_in(22), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(22));
   FF_23 : FD_201 port map( D => data_in(23), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(23));
   FF_24 : FD_200 port map( D => data_in(24), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(24));
   FF_25 : FD_199 port map( D => data_in(25), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(25));
   FF_26 : FD_198 port map( D => data_in(26), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(26));
   FF_27 : FD_197 port map( D => data_in(27), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(27));
   FF_28 : FD_196 port map( D => data_in(28), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(28));
   FF_29 : FD_195 port map( D => data_in(29), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(29));
   FF_30 : FD_194 port map( D => data_in(30), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(30));
   FF_31 : FD_193 port map( D => data_in(31), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(31));
   U1 : BUF_X1 port map( A => n12, Z => n11);
   U2 : BUF_X1 port map( A => ENABLE, Z => n12);
   U3 : BUF_X1 port map( A => RESET, Z => n16);
   U4 : BUF_X2 port map( A => n12, Z => n10);
   U5 : BUF_X2 port map( A => n12, Z => n9);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_6 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_6;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_161
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_162
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_163
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_164
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_165
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_166
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_167
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_168
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_169
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_170
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_171
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_172
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_173
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_174
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_175
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_176
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_177
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_178
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_179
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_180
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_181
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_182
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_183
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_184
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_185
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_186
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_187
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_188
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_189
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_190
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_191
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_192
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12 : std_logic;

begin
   
   FF_0 : FD_192 port map( D => data_in(0), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_191 port map( D => data_in(1), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_190 port map( D => data_in(2), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_189 port map( D => data_in(3), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_188 port map( D => data_in(4), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_187 port map( D => data_in(5), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_186 port map( D => data_in(6), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_185 port map( D => data_in(7), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_184 port map( D => data_in(8), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_183 port map( D => data_in(9), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_182 port map( D => data_in(10), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_181 port map( D => data_in(11), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_180 port map( D => data_in(12), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(12));
   FF_13 : FD_179 port map( D => data_in(13), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(13));
   FF_14 : FD_178 port map( D => data_in(14), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(14));
   FF_15 : FD_177 port map( D => data_in(15), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(15));
   FF_16 : FD_176 port map( D => data_in(16), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(16));
   FF_17 : FD_175 port map( D => data_in(17), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(17));
   FF_18 : FD_174 port map( D => data_in(18), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(18));
   FF_19 : FD_173 port map( D => data_in(19), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(19));
   FF_20 : FD_172 port map( D => data_in(20), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(20));
   FF_21 : FD_171 port map( D => data_in(21), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(21));
   FF_22 : FD_170 port map( D => data_in(22), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(22));
   FF_23 : FD_169 port map( D => data_in(23), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(23));
   FF_24 : FD_168 port map( D => data_in(24), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(24));
   FF_25 : FD_167 port map( D => data_in(25), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(25));
   FF_26 : FD_166 port map( D => data_in(26), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(26));
   FF_27 : FD_165 port map( D => data_in(27), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(27));
   FF_28 : FD_164 port map( D => data_in(28), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(28));
   FF_29 : FD_163 port map( D => data_in(29), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(29));
   FF_30 : FD_162 port map( D => data_in(30), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(30));
   FF_31 : FD_161 port map( D => data_in(31), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => n12, Z => n9);
   U3 : BUF_X1 port map( A => n12, Z => n10);
   U4 : BUF_X1 port map( A => n12, Z => n11);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_10 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_10;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_10 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_289
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_290
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_291
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_292
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_293
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_294
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_295
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_296
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_297
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_298
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_299
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_300
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_301
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_302
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_303
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_304
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_305
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_306
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_307
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_308
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_309
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_310
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_311
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_312
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_313
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_314
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_315
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_316
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_317
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_318
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_319
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_320
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12 : std_logic;

begin
   
   FF_0 : FD_320 port map( D => data_in(0), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_319 port map( D => data_in(1), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_318 port map( D => data_in(2), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_317 port map( D => data_in(3), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_316 port map( D => data_in(4), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_315 port map( D => data_in(5), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_314 port map( D => data_in(6), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_313 port map( D => data_in(7), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_312 port map( D => data_in(8), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_311 port map( D => data_in(9), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_310 port map( D => data_in(10), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_309 port map( D => data_in(11), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_308 port map( D => data_in(12), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(12));
   FF_13 : FD_307 port map( D => data_in(13), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(13));
   FF_14 : FD_306 port map( D => data_in(14), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(14));
   FF_15 : FD_305 port map( D => data_in(15), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(15));
   FF_16 : FD_304 port map( D => data_in(16), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(16));
   FF_17 : FD_303 port map( D => data_in(17), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(17));
   FF_18 : FD_302 port map( D => data_in(18), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(18));
   FF_19 : FD_301 port map( D => data_in(19), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(19));
   FF_20 : FD_300 port map( D => data_in(20), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(20));
   FF_21 : FD_299 port map( D => data_in(21), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(21));
   FF_22 : FD_298 port map( D => data_in(22), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(22));
   FF_23 : FD_297 port map( D => data_in(23), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(23));
   FF_24 : FD_296 port map( D => data_in(24), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(24));
   FF_25 : FD_295 port map( D => data_in(25), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(25));
   FF_26 : FD_294 port map( D => data_in(26), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(26));
   FF_27 : FD_293 port map( D => data_in(27), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(27));
   FF_28 : FD_292 port map( D => data_in(28), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(28));
   FF_29 : FD_291 port map( D => data_in(29), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(29));
   FF_30 : FD_290 port map( D => data_in(30), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(30));
   FF_31 : FD_289 port map( D => data_in(31), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => n12, Z => n9);
   U3 : BUF_X1 port map( A => n12, Z => n10);
   U4 : BUF_X1 port map( A => n12, Z => n11);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_9 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_9;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_9 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_257
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_258
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_259
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_260
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_261
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_262
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_263
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_264
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_265
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_266
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_267
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_268
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_269
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_270
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_271
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_272
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_273
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_274
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_275
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_276
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_277
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_278
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_279
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_280
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_281
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_282
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_283
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_284
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_285
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_286
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_287
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_288
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12 : std_logic;

begin
   
   FF_0 : FD_288 port map( D => data_in(0), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_287 port map( D => data_in(1), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_286 port map( D => data_in(2), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_285 port map( D => data_in(3), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_284 port map( D => data_in(4), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_283 port map( D => data_in(5), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_282 port map( D => data_in(6), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_281 port map( D => data_in(7), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_280 port map( D => data_in(8), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_279 port map( D => data_in(9), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_278 port map( D => data_in(10), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_277 port map( D => data_in(11), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_276 port map( D => data_in(12), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(12));
   FF_13 : FD_275 port map( D => data_in(13), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(13));
   FF_14 : FD_274 port map( D => data_in(14), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(14));
   FF_15 : FD_273 port map( D => data_in(15), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(15));
   FF_16 : FD_272 port map( D => data_in(16), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(16));
   FF_17 : FD_271 port map( D => data_in(17), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(17));
   FF_18 : FD_270 port map( D => data_in(18), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(18));
   FF_19 : FD_269 port map( D => data_in(19), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(19));
   FF_20 : FD_268 port map( D => data_in(20), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(20));
   FF_21 : FD_267 port map( D => data_in(21), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(21));
   FF_22 : FD_266 port map( D => data_in(22), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(22));
   FF_23 : FD_265 port map( D => data_in(23), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(23));
   FF_24 : FD_264 port map( D => data_in(24), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(24));
   FF_25 : FD_263 port map( D => data_in(25), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(25));
   FF_26 : FD_262 port map( D => data_in(26), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(26));
   FF_27 : FD_261 port map( D => data_in(27), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(27));
   FF_28 : FD_260 port map( D => data_in(28), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(28));
   FF_29 : FD_259 port map( D => data_in(29), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(29));
   FF_30 : FD_258 port map( D => data_in(30), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(30));
   FF_31 : FD_257 port map( D => data_in(31), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => n12, Z => n9);
   U3 : BUF_X1 port map( A => n12, Z => n10);
   U4 : BUF_X1 port map( A => n12, Z => n11);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_5 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_5;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_5 is

   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_129
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_130
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_131
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_132
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_133
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_134
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_135
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_136
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_137
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_138
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_139
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_140
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_141
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_142
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_143
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_144
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_145
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_146
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_147
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_148
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_149
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_150
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_151
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_152
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_153
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_154
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_155
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_156
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_157
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_158
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_159
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_160
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_160 port map( D => data_in(0), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(0));
   FF_1 : FD_159 port map( D => data_in(1), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(1));
   FF_2 : FD_158 port map( D => data_in(2), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(2));
   FF_3 : FD_157 port map( D => data_in(3), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(3));
   FF_4 : FD_156 port map( D => data_in(4), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(4));
   FF_5 : FD_155 port map( D => data_in(5), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(5));
   FF_6 : FD_154 port map( D => data_in(6), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(6));
   FF_7 : FD_153 port map( D => data_in(7), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(7));
   FF_8 : FD_152 port map( D => data_in(8), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(8));
   FF_9 : FD_151 port map( D => data_in(9), CK => CK, RESET => n13, ENABLE => 
                           n9, Q => data_out(9));
   FF_10 : FD_150 port map( D => data_in(10), CK => CK, RESET => n13, ENABLE =>
                           n9, Q => data_out(10));
   FF_11 : FD_149 port map( D => data_in(11), CK => CK, RESET => n13, ENABLE =>
                           n9, Q => data_out(11));
   FF_12 : FD_148 port map( D => data_in(12), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(12));
   FF_13 : FD_147 port map( D => data_in(13), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(13));
   FF_14 : FD_146 port map( D => data_in(14), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(14));
   FF_15 : FD_145 port map( D => data_in(15), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(15));
   FF_16 : FD_144 port map( D => data_in(16), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(16));
   FF_17 : FD_143 port map( D => data_in(17), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(17));
   FF_18 : FD_142 port map( D => data_in(18), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(18));
   FF_19 : FD_141 port map( D => data_in(19), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(19));
   FF_20 : FD_140 port map( D => data_in(20), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(20));
   FF_21 : FD_139 port map( D => data_in(21), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(21));
   FF_22 : FD_138 port map( D => data_in(22), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(22));
   FF_23 : FD_137 port map( D => data_in(23), CK => CK, RESET => n14, ENABLE =>
                           n10, Q => data_out(23));
   FF_24 : FD_136 port map( D => data_in(24), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(24));
   FF_25 : FD_135 port map( D => data_in(25), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(25));
   FF_26 : FD_134 port map( D => data_in(26), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(26));
   FF_27 : FD_133 port map( D => data_in(27), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(27));
   FF_28 : FD_132 port map( D => data_in(28), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(28));
   FF_29 : FD_131 port map( D => data_in(29), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(29));
   FF_30 : FD_130 port map( D => data_in(30), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(30));
   FF_31 : FD_129 port map( D => data_in(31), CK => CK, RESET => n15, ENABLE =>
                           n11, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n16);
   U2 : BUF_X1 port map( A => n12, Z => n11);
   U3 : BUF_X1 port map( A => ENABLE, Z => n12);
   U4 : BUF_X1 port map( A => n16, Z => n13);
   U5 : BUF_X1 port map( A => n16, Z => n14);
   U6 : BUF_X1 port map( A => n16, Z => n15);
   U7 : BUF_X2 port map( A => n12, Z => n9);
   U8 : BUF_X2 port map( A => n12, Z => n10);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_4 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_4;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_97
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_98
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_99
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_100
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_101
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_102
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_103
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_104
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_105
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_106
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_107
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_108
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_109
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_110
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_111
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_112
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_113
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_114
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_115
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_116
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_117
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_118
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_119
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_120
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_121
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_122
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_123
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_124
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_125
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_126
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_127
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_128
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12 : std_logic;

begin
   
   FF_0 : FD_128 port map( D => data_in(0), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_127 port map( D => data_in(1), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_126 port map( D => data_in(2), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_125 port map( D => data_in(3), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_124 port map( D => data_in(4), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_123 port map( D => data_in(5), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_122 port map( D => data_in(6), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_121 port map( D => data_in(7), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_120 port map( D => data_in(8), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_119 port map( D => data_in(9), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_118 port map( D => data_in(10), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_117 port map( D => data_in(11), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_116 port map( D => data_in(12), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(12));
   FF_13 : FD_115 port map( D => data_in(13), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(13));
   FF_14 : FD_114 port map( D => data_in(14), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(14));
   FF_15 : FD_113 port map( D => data_in(15), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(15));
   FF_16 : FD_112 port map( D => data_in(16), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(16));
   FF_17 : FD_111 port map( D => data_in(17), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(17));
   FF_18 : FD_110 port map( D => data_in(18), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(18));
   FF_19 : FD_109 port map( D => data_in(19), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(19));
   FF_20 : FD_108 port map( D => data_in(20), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(20));
   FF_21 : FD_107 port map( D => data_in(21), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(21));
   FF_22 : FD_106 port map( D => data_in(22), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(22));
   FF_23 : FD_105 port map( D => data_in(23), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(23));
   FF_24 : FD_104 port map( D => data_in(24), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(24));
   FF_25 : FD_103 port map( D => data_in(25), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(25));
   FF_26 : FD_102 port map( D => data_in(26), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(26));
   FF_27 : FD_101 port map( D => data_in(27), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(27));
   FF_28 : FD_100 port map( D => data_in(28), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(28));
   FF_29 : FD_99 port map( D => data_in(29), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_98 port map( D => data_in(30), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_97 port map( D => data_in(31), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => n12, Z => n9);
   U3 : BUF_X1 port map( A => n12, Z => n10);
   U4 : BUF_X1 port map( A => n12, Z => n11);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_3 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_3;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_65
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_66
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_67
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_68
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_69
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_70
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_71
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_72
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_73
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_74
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_75
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_76
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_77
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_78
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_79
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_80
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_81
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_82
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_83
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_84
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_85
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_86
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_87
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_88
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_89
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_90
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_91
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_92
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_93
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_94
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_95
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_96
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12 : std_logic;

begin
   
   FF_0 : FD_96 port map( D => data_in(0), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_95 port map( D => data_in(1), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_94 port map( D => data_in(2), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_93 port map( D => data_in(3), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_92 port map( D => data_in(4), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_91 port map( D => data_in(5), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_90 port map( D => data_in(6), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_89 port map( D => data_in(7), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_88 port map( D => data_in(8), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_87 port map( D => data_in(9), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_86 port map( D => data_in(10), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_85 port map( D => data_in(11), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_84 port map( D => data_in(12), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_83 port map( D => data_in(13), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_82 port map( D => data_in(14), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_81 port map( D => data_in(15), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_80 port map( D => data_in(16), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_79 port map( D => data_in(17), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_78 port map( D => data_in(18), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_77 port map( D => data_in(19), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_76 port map( D => data_in(20), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_75 port map( D => data_in(21), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_74 port map( D => data_in(22), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_73 port map( D => data_in(23), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_72 port map( D => data_in(24), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_71 port map( D => data_in(25), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_70 port map( D => data_in(26), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_69 port map( D => data_in(27), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_68 port map( D => data_in(28), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_67 port map( D => data_in(29), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_66 port map( D => data_in(30), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_65 port map( D => data_in(31), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => n12, Z => n9);
   U3 : BUF_X1 port map( A => n12, Z => n10);
   U4 : BUF_X1 port map( A => n12, Z => n11);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_2 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_2;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_33
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_34
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_35
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_36
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_37
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_38
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_39
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_40
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_41
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_42
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_43
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_44
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_45
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_46
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_47
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_48
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_49
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_50
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_51
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_52
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_53
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_54
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_55
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_56
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_57
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_58
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_59
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_60
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_61
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_62
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_63
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_64
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12 : std_logic;

begin
   
   FF_0 : FD_64 port map( D => data_in(0), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_63 port map( D => data_in(1), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_62 port map( D => data_in(2), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_61 port map( D => data_in(3), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_60 port map( D => data_in(4), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_59 port map( D => data_in(5), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_58 port map( D => data_in(6), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_57 port map( D => data_in(7), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_56 port map( D => data_in(8), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_55 port map( D => data_in(9), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_54 port map( D => data_in(10), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_53 port map( D => data_in(11), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_52 port map( D => data_in(12), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_51 port map( D => data_in(13), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_50 port map( D => data_in(14), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_49 port map( D => data_in(15), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_48 port map( D => data_in(16), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_47 port map( D => data_in(17), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_46 port map( D => data_in(18), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_45 port map( D => data_in(19), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_44 port map( D => data_in(20), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_43 port map( D => data_in(21), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_42 port map( D => data_in(22), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_41 port map( D => data_in(23), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_40 port map( D => data_in(24), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_39 port map( D => data_in(25), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_38 port map( D => data_in(26), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_37 port map( D => data_in(27), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_36 port map( D => data_in(28), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_35 port map( D => data_in(29), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_34 port map( D => data_in(30), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_33 port map( D => data_in(31), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => n12, Z => n9);
   U3 : BUF_X1 port map( A => n12, Z => n10);
   U4 : BUF_X1 port map( A => n12, Z => n11);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_1 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_1;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_3
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_4
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_5
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_6
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_7
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_8
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_9
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_10
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_11
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_12
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_13
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_14
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_15
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_16
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_17
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_18
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_19
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_20
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_21
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_22
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_23
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_24
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_25
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_26
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_27
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_28
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_29
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_30
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_31
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_32
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12 : std_logic;

begin
   
   FF_0 : FD_32 port map( D => data_in(0), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_31 port map( D => data_in(1), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_30 port map( D => data_in(2), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_29 port map( D => data_in(3), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_28 port map( D => data_in(4), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_27 port map( D => data_in(5), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_26 port map( D => data_in(6), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_25 port map( D => data_in(7), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_24 port map( D => data_in(8), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_23 port map( D => data_in(9), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_22 port map( D => data_in(10), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_21 port map( D => data_in(11), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_20 port map( D => data_in(12), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_19 port map( D => data_in(13), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_18 port map( D => data_in(14), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_17 port map( D => data_in(15), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_16 port map( D => data_in(16), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_15 port map( D => data_in(17), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_14 port map( D => data_in(18), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_13 port map( D => data_in(19), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_12 port map( D => data_in(20), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_11 port map( D => data_in(21), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_10 port map( D => data_in(22), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_9 port map( D => data_in(23), CK => CK, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_8 port map( D => data_in(24), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_7 port map( D => data_in(25), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_6 port map( D => data_in(26), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_5 port map( D => data_in(27), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_4 port map( D => data_in(28), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_3 port map( D => data_in(29), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_2 port map( D => data_in(30), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_1 port map( D => data_in(31), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => n12, Z => n9);
   U3 : BUF_X1 port map( A => n12, Z => n10);
   U4 : BUF_X1 port map( A => n12, Z => n11);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_7;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n13);
   U2 : INV_X1 port map( A => n7, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => S, B1 => B(2), B2 => n13, ZN => n7
                           );
   U4 : INV_X1 port map( A => n6, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => S, A2 => A(3), B1 => B(3), B2 => n13, ZN => n6
                           );
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => S, B1 => B(1), B2 => n13, ZN => n8
                           );
   U8 : INV_X1 port map( A => n9, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => S, B1 => B(0), B2 => n13, ZN => n9
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_0;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n5, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n10, ZN => n5);
   U2 : INV_X1 port map( A => n7, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n10, B1 => B(2), B2 => n5, ZN => 
                           n7);
   U4 : BUF_X1 port map( A => S, Z => n10);
   U5 : INV_X1 port map( A => n6, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => n10, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n6);
   U7 : INV_X1 port map( A => n8, ZN => Y(1));
   U8 : AOI22_X1 port map( A1 => A(1), A2 => n10, B1 => B(1), B2 => n5, ZN => 
                           n8);
   U9 : INV_X1 port map( A => n9, ZN => Y(0));
   U10 : AOI22_X1 port map( A1 => A(0), A2 => n10, B1 => B(0), B2 => n5, ZN => 
                           n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_0;

architecture SYN_BEHAVIORAL of RCA_NBITS4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30 : std_logic;

begin
   
   U25 : XOR2_X1 port map( A => n9, B => n10, Z => S(3));
   U26 : XOR2_X1 port map( A => n23, B => A(3), Z => n10);
   U27 : XOR2_X1 port map( A => n11, B => n12, Z => S(2));
   U28 : XOR2_X1 port map( A => n14, B => n15, Z => S(1));
   U2 : NOR2_X1 port map( A1 => n29, A2 => n26, ZN => n16);
   U3 : INV_X1 port map( A => n20, ZN => n23);
   U4 : AOI21_X1 port map( B1 => n26, B2 => n29, A => n16, ZN => n17);
   U5 : OAI21_X1 port map( B1 => n28, B2 => n23, A => n19, ZN => Co);
   U6 : AOI21_X1 port map( B1 => n16, B2 => A(1), A => n25, ZN => n13);
   U7 : INV_X1 port map( A => n22, ZN => n25);
   U8 : OAI21_X1 port map( B1 => n16, B2 => A(1), A => B(1), ZN => n22);
   U9 : AOI21_X1 port map( B1 => n27, B2 => n13, A => n21, ZN => n20);
   U10 : INV_X1 port map( A => A(2), ZN => n27);
   U11 : AOI21_X1 port map( B1 => n24, B2 => A(2), A => B(2), ZN => n21);
   U12 : INV_X1 port map( A => n13, ZN => n24);
   U13 : INV_X1 port map( A => A(0), ZN => n26);
   U14 : INV_X1 port map( A => B(0), ZN => n29);
   U15 : XNOR2_X1 port map( A => A(2), B => n13, ZN => n11);
   U16 : XNOR2_X1 port map( A => n16, B => A(1), ZN => n15);
   U17 : XNOR2_X1 port map( A => A(0), B => B(0), ZN => n18);
   U18 : OAI21_X1 port map( B1 => n20, B2 => A(3), A => B(3), ZN => n19);
   U19 : INV_X1 port map( A => A(3), ZN => n28);
   U20 : XNOR2_X1 port map( A => n30, B => B(2), ZN => n12);
   U21 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n9);
   U22 : OAI22_X1 port map( A1 => n17, A2 => n30, B1 => Ci, B2 => n18, ZN => 
                           S(0));
   U23 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n14);
   U24 : INV_X1 port map( A => Ci, ZN => n30);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_0 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_0;

architecture SYN_BEHAVIORAL of PG_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);
   U2 : INV_X1 port map( A => n2, ZN => G_ij);
   U3 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_0 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_0;

architecture SYN_BEHAVIORAL of G_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_0 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_0;

architecture SYN_BEHAVIORAL of pg_generator_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_7;

architecture SYN_STRUCTURAL of CarrySelect_7 is

   component MUX21_GENERIC_bits4_7
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1012, n_1013 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1012);
   RCA2 : RCA_NBITS4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1013);
   MUX21_GEN : MUX21_GENERIC_bits4_7 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_0;

architecture SYN_STRUCTURAL of CarrySelect_0 is

   component MUX21_GENERIC_bits4_0
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1014, n_1015 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1014);
   RCA2 : RCA_NBITS4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1015);
   MUX21_GEN : MUX21_GENERIC_bits4_0 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity logic_and_shift_N32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end logic_and_shift_N32_DW01_ash_0;

architecture SYN_mx2 of logic_and_shift_N32_DW01_ash_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal temp_int_SH_4_port, SHMAG_5_port, ML_int_1_31_port, ML_int_1_30_port,
      ML_int_1_29_port, ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, 
      ML_int_1_25_port, ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, 
      ML_int_1_21_port, ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, 
      ML_int_1_17_port, ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, 
      ML_int_1_13_port, ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, 
      ML_int_1_9_port, ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, 
      ML_int_1_5_port, ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, 
      ML_int_1_1_port, ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, 
      ML_int_2_29_port, ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, 
      ML_int_2_25_port, ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, 
      ML_int_2_21_port, ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, 
      ML_int_2_17_port, ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, 
      ML_int_2_13_port, ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, 
      ML_int_2_9_port, ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, 
      ML_int_2_5_port, ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, 
      ML_int_2_1_port, ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, 
      ML_int_3_29_port, ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, 
      ML_int_3_25_port, ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, 
      ML_int_3_21_port, ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, 
      ML_int_3_17_port, ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, 
      ML_int_3_13_port, ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, 
      ML_int_3_9_port, ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, 
      ML_int_3_5_port, ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, 
      ML_int_3_1_port, ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, 
      ML_int_4_29_port, ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, 
      ML_int_4_25_port, ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, 
      ML_int_4_21_port, ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, 
      ML_int_4_17_port, ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, 
      ML_int_4_13_port, ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, 
      ML_int_4_9_port, ML_int_4_8_port, ML_int_5_31_port, ML_int_5_30_port, 
      ML_int_5_29_port, ML_int_5_28_port, ML_int_5_27_port, ML_int_5_26_port, 
      ML_int_5_25_port, ML_int_5_24_port, ML_int_5_23_port, ML_int_5_22_port, 
      ML_int_5_21_port, ML_int_5_20_port, ML_int_5_19_port, ML_int_5_18_port, 
      ML_int_5_17_port, ML_int_5_16_port, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_31_port);
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_30_port);
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_29_port);
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_28_port);
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_27_port);
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_26_port);
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_25_port);
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_24_port);
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => n88, S => 
                           temp_int_SH_4_port, Z => ML_int_5_23_port);
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => n84, S => 
                           temp_int_SH_4_port, Z => ML_int_5_22_port);
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => n86, S => 
                           temp_int_SH_4_port, Z => ML_int_5_21_port);
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => n82, S => 
                           temp_int_SH_4_port, Z => ML_int_5_20_port);
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => n87, S => 
                           temp_int_SH_4_port, Z => ML_int_5_19_port);
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => n83, S => 
                           temp_int_SH_4_port, Z => ML_int_5_18_port);
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => n85, S => 
                           temp_int_SH_4_port, Z => ML_int_5_17_port);
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => n81, S => 
                           temp_int_SH_4_port, Z => ML_int_5_16_port);
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => n80, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => n80, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => n80, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => n80, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => n80, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => n80, Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => n80, Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => n80, Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => n80, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => n80, Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => n80, Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => n80, Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => n79, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => n79, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => n79, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => n79, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => n79, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => n79, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => n79, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => n79, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => n79, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => n79, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           n79, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           n79, Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => n76, Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => n75, Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => n76, Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => n75, Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => n76, Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => n76, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => n76, Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => n76, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => n76, Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => n76, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => n76, Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => n76, Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => n76, Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => n76, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => n76, Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => n76, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => n75, Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => n75, Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => n75, Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => n75, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => n75, Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => n75, Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           n75, Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           n75, Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           n75, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           n75, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           n75, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           n75, Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => n71, Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => n72, Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => n71, Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => n72, Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => n71, Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => n72, Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => n72, Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => n72, Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => n72, Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => n72, Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => n72, Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => n72, Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => n72, Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => n72, Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => n72, Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => n72, Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => n72, Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => n72, Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => n71, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => n71, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => n71, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => n71, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           n71, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           n71, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           n71, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           n71, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           n71, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           n71, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           n71, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           n71, Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => n68, Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => n69, Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => n68, Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => n69, Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => n68, Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => n69, Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => n68, Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => n69, Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => n69, Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => n69, Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => n69, Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => n69, Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => n69, Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => n69, Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => n69, Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => n69, Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => n69, Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => n69, Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => n69, Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => n68, Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => n68, Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => n68, Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => n68, Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => n68, Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => n68, Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => n68, Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => n68, Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => n68, Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => n68, Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => n68, Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => n68, Z => 
                           ML_int_1_1_port);
   U94 : NAND3_X1 port map( A1 => SH(11), A2 => SH(10), A3 => SH(12), ZN => n51
                           );
   U96 : NAND3_X1 port map( A1 => SH(17), A2 => SH(16), A3 => SH(18), ZN => n52
                           );
   U98 : NAND3_X1 port map( A1 => SH(23), A2 => SH(22), A3 => SH(24), ZN => n53
                           );
   U100 : NAND3_X1 port map( A1 => SH(29), A2 => SH(28), A3 => SH(6), ZN => n54
                           );
   U104 : NAND3_X1 port map( A1 => n92, A2 => n93, A3 => n91, ZN => n60);
   U106 : NAND3_X1 port map( A1 => n101, A2 => n102, A3 => n100, ZN => n61);
   U108 : NAND3_X1 port map( A1 => n98, A2 => n99, A3 => n97, ZN => n62);
   U110 : NAND3_X1 port map( A1 => n95, A2 => n96, A3 => n94, ZN => n63);
   U3 : AND2_X1 port map( A1 => n38, A2 => n45, ZN => n64);
   U4 : AND2_X1 port map( A1 => n38, A2 => n42, ZN => n65);
   U5 : AND2_X1 port map( A1 => n38, A2 => n44, ZN => n66);
   U6 : AND2_X1 port map( A1 => n38, A2 => n43, ZN => n67);
   U7 : BUF_X1 port map( A => n64, Z => n70);
   U8 : BUF_X1 port map( A => n66, Z => n73);
   U9 : BUF_X1 port map( A => n67, Z => n77);
   U10 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n89, ZN => B(8));
   U11 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n89, ZN => B(9));
   U12 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n89, ZN => B(10));
   U13 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n89, ZN => B(11));
   U14 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n89, ZN => B(12));
   U15 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n89, ZN => B(13));
   U16 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n89, ZN => B(14));
   U17 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n89, ZN => B(15));
   U18 : INV_X1 port map( A => n28, ZN => n89);
   U19 : NOR2_X1 port map( A1 => n28, A2 => n37, ZN => B(0));
   U20 : NOR2_X1 port map( A1 => n28, A2 => n36, ZN => B(1));
   U21 : NOR2_X1 port map( A1 => n28, A2 => n35, ZN => B(2));
   U22 : NOR2_X1 port map( A1 => n28, A2 => n33, ZN => B(3));
   U23 : NOR2_X1 port map( A1 => n28, A2 => n32, ZN => B(4));
   U24 : NOR2_X1 port map( A1 => n28, A2 => n31, ZN => B(5));
   U25 : NOR2_X1 port map( A1 => n28, A2 => n30, ZN => B(6));
   U26 : NOR2_X1 port map( A1 => n28, A2 => n29, ZN => B(7));
   U27 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => n78, ZN => 
                           ML_int_3_2_port);
   U28 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => n78, ZN => 
                           ML_int_3_3_port);
   U29 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => n78, ZN => 
                           ML_int_3_0_port);
   U30 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => n78, ZN => 
                           ML_int_3_1_port);
   U31 : INV_X1 port map( A => n70, ZN => n68);
   U32 : INV_X1 port map( A => n70, ZN => n69);
   U33 : INV_X1 port map( A => n73, ZN => n71);
   U34 : INV_X1 port map( A => n73, ZN => n72);
   U35 : INV_X1 port map( A => n77, ZN => n76);
   U36 : INV_X1 port map( A => n77, ZN => n75);
   U37 : NAND2_X1 port map( A1 => n34, A2 => n90, ZN => n28);
   U38 : INV_X1 port map( A => temp_int_SH_4_port, ZN => n90);
   U39 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => n65, ZN => n37);
   U40 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => n65, ZN => n36);
   U41 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => n65, ZN => n35);
   U42 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => n65, ZN => n33);
   U43 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => n65, ZN => n32);
   U44 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => n65, ZN => n31);
   U45 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => n65, ZN => n30);
   U46 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => n65, ZN => n29);
   U47 : AND2_X1 port map( A1 => ML_int_5_16_port, A2 => n34, ZN => B(16));
   U48 : INV_X1 port map( A => n37, ZN => n81);
   U49 : AND2_X1 port map( A1 => ML_int_5_17_port, A2 => n34, ZN => B(17));
   U50 : INV_X1 port map( A => n36, ZN => n85);
   U51 : AND2_X1 port map( A1 => ML_int_5_18_port, A2 => n34, ZN => B(18));
   U52 : INV_X1 port map( A => n35, ZN => n83);
   U53 : AND2_X1 port map( A1 => ML_int_5_19_port, A2 => n34, ZN => B(19));
   U54 : INV_X1 port map( A => n33, ZN => n87);
   U55 : AND2_X1 port map( A1 => ML_int_5_20_port, A2 => n34, ZN => B(20));
   U56 : INV_X1 port map( A => n32, ZN => n82);
   U57 : AND2_X1 port map( A1 => ML_int_5_21_port, A2 => n34, ZN => B(21));
   U58 : INV_X1 port map( A => n31, ZN => n86);
   U59 : AND2_X1 port map( A1 => ML_int_5_22_port, A2 => n34, ZN => B(22));
   U60 : INV_X1 port map( A => n30, ZN => n84);
   U61 : AND2_X1 port map( A1 => ML_int_5_23_port, A2 => n34, ZN => B(23));
   U62 : INV_X1 port map( A => n29, ZN => n88);
   U63 : AND2_X1 port map( A1 => ML_int_5_24_port, A2 => n34, ZN => B(24));
   U64 : AND2_X1 port map( A1 => ML_int_5_25_port, A2 => n34, ZN => B(25));
   U65 : AND2_X1 port map( A1 => ML_int_5_26_port, A2 => n34, ZN => B(26));
   U66 : AND2_X1 port map( A1 => ML_int_5_27_port, A2 => n34, ZN => B(27));
   U67 : AND2_X1 port map( A1 => ML_int_5_28_port, A2 => n34, ZN => B(28));
   U68 : AND2_X1 port map( A1 => ML_int_5_29_port, A2 => n34, ZN => B(29));
   U69 : AND2_X1 port map( A1 => ML_int_5_30_port, A2 => n34, ZN => B(30));
   U70 : AND2_X1 port map( A1 => ML_int_5_31_port, A2 => n34, ZN => B(31));
   U71 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => n74, ZN => 
                           ML_int_2_1_port);
   U72 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => n74, ZN => 
                           ML_int_2_0_port);
   U73 : INV_X1 port map( A => n65, ZN => n80);
   U74 : INV_X1 port map( A => n65, ZN => n79);
   U75 : BUF_X1 port map( A => n67, Z => n78);
   U76 : BUF_X1 port map( A => n66, Z => n74);
   U77 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => temp_int_SH_4_port);
   U78 : NAND2_X1 port map( A1 => SH(4), A2 => n40, ZN => n39);
   U79 : NOR4_X1 port map( A1 => n51, A2 => n96, A3 => n94, A4 => n95, ZN => 
                           n50);
   U80 : NOR4_X1 port map( A1 => n60, A2 => SH(28), A3 => SH(6), A4 => SH(29), 
                           ZN => n59);
   U81 : NOR4_X1 port map( A1 => n52, A2 => n99, A3 => n97, A4 => n98, ZN => 
                           n49);
   U82 : NOR4_X1 port map( A1 => n61, A2 => SH(22), A3 => SH(24), A4 => SH(23),
                           ZN => n58);
   U83 : NAND2_X1 port map( A1 => SH(30), A2 => n46, ZN => n40);
   U84 : NAND4_X1 port map( A1 => n47, A2 => n48, A3 => n49, A4 => n50, ZN => 
                           n46);
   U85 : NOR4_X1 port map( A1 => n54, A2 => n93, A3 => n91, A4 => n92, ZN => 
                           n47);
   U86 : NOR4_X1 port map( A1 => n53, A2 => n102, A3 => n100, A4 => n101, ZN =>
                           n48);
   U87 : NAND2_X1 port map( A1 => n55, A2 => n103, ZN => n38);
   U88 : NAND4_X1 port map( A1 => n56, A2 => n57, A3 => n58, A4 => n59, ZN => 
                           n55);
   U89 : NOR4_X1 port map( A1 => n63, A2 => SH(10), A3 => SH(12), A4 => SH(11),
                           ZN => n56);
   U90 : NOR4_X1 port map( A1 => n62, A2 => SH(16), A3 => SH(18), A4 => SH(17),
                           ZN => n57);
   U91 : AND2_X1 port map( A1 => SHMAG_5_port, A2 => n103, ZN => n34);
   U92 : AND2_X1 port map( A1 => n38, A2 => n41, ZN => SHMAG_5_port);
   U93 : NAND2_X1 port map( A1 => SH(5), A2 => n40, ZN => n41);
   U95 : NAND2_X1 port map( A1 => SH(0), A2 => n40, ZN => n45);
   U97 : NAND2_X1 port map( A1 => SH(1), A2 => n40, ZN => n44);
   U99 : NAND2_X1 port map( A1 => SH(2), A2 => n40, ZN => n43);
   U101 : NAND2_X1 port map( A1 => SH(3), A2 => n40, ZN => n42);
   U102 : INV_X1 port map( A => SH(30), ZN => n103);
   U103 : INV_X1 port map( A => SH(26), ZN => n101);
   U105 : INV_X1 port map( A => SH(14), ZN => n95);
   U107 : INV_X1 port map( A => SH(25), ZN => n100);
   U109 : INV_X1 port map( A => SH(13), ZN => n94);
   U111 : INV_X1 port map( A => SH(15), ZN => n96);
   U112 : INV_X1 port map( A => SH(27), ZN => n102);
   U113 : INV_X1 port map( A => SH(8), ZN => n92);
   U114 : INV_X1 port map( A => SH(20), ZN => n98);
   U115 : INV_X1 port map( A => SH(19), ZN => n97);
   U116 : INV_X1 port map( A => SH(7), ZN => n91);
   U117 : INV_X1 port map( A => SH(21), ZN => n99);
   U118 : INV_X1 port map( A => SH(9), ZN => n93);
   U119 : AND2_X1 port map( A1 => A(0), A2 => n64, ZN => ML_int_1_0_port);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity logic_and_shift_N32_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end logic_and_shift_N32_DW_rash_0;

architecture SYN_mx2 of logic_and_shift_N32_DW_rash_0 is

   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247 : std_logic;

begin
   
   U81 : MUX2_X1 port map( A => n193, B => n102, S => SH(4), Z => n94);
   U89 : MUX2_X1 port map( A => n112, B => n214, S => SH(4), Z => n111);
   U113 : MUX2_X1 port map( A => n133, B => n213, S => SH(4), Z => n132);
   U151 : MUX2_X1 port map( A => n125, B => n107, S => SH(2), Z => n120);
   U195 : MUX2_X1 port map( A => n178, B => n210, S => SH(4), Z => n177);
   U3 : NOR2_X1 port map( A1 => n243, A2 => SH(3), ZN => n123);
   U4 : NOR2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n122);
   U5 : NOR2_X1 port map( A1 => n246, A2 => n242, ZN => n67);
   U6 : NOR2_X1 port map( A1 => n91, A2 => n246, ZN => B(20));
   U7 : NOR2_X1 port map( A1 => n88, A2 => n246, ZN => B(21));
   U8 : NOR2_X1 port map( A1 => n82, A2 => n246, ZN => B(22));
   U9 : NOR2_X1 port map( A1 => n141, A2 => n246, ZN => B(16));
   U10 : NOR2_X1 port map( A1 => n134, A2 => n246, ZN => B(17));
   U11 : NOR2_X1 port map( A1 => n113, A2 => n246, ZN => B(18));
   U12 : NOR2_X1 port map( A1 => n72, A2 => n246, ZN => B(24));
   U13 : NOR2_X1 port map( A1 => n63, A2 => n246, ZN => B(25));
   U14 : NOR2_X1 port map( A1 => n121, A2 => n246, ZN => B(26));
   U15 : NOR2_X1 port map( A1 => n220, A2 => n246, ZN => B(23));
   U16 : INV_X1 port map( A => n141, ZN => n210);
   U17 : INV_X1 port map( A => n134, ZN => n213);
   U18 : INV_X1 port map( A => n113, ZN => n214);
   U19 : INV_X1 port map( A => n100, ZN => n237);
   U20 : INV_X1 port map( A => n101, ZN => n239);
   U21 : NAND2_X1 port map( A1 => n122, A2 => n163, ZN => n62);
   U22 : AOI222_X1 port map( A1 => n222, A2 => n123, B1 => n231, B2 => n241, C1
                           => n74, C2 => n122, ZN => n91);
   U23 : AOI222_X1 port map( A1 => n224, A2 => n123, B1 => n233, B2 => n241, C1
                           => n66, C2 => n122, ZN => n88);
   U24 : AOI222_X1 port map( A1 => n227, A2 => n123, B1 => n234, B2 => n241, C1
                           => n127, C2 => n122, ZN => n82);
   U25 : INV_X1 port map( A => n116, ZN => n236);
   U26 : INV_X1 port map( A => n163, ZN => n246);
   U27 : INV_X1 port map( A => n117, ZN => n240);
   U28 : AOI221_X1 port map( B1 => n74, B2 => n123, C1 => n75, C2 => n122, A =>
                           n179, ZN => n141);
   U29 : OAI22_X1 port map( A1 => n104, A2 => n119, B1 => n105, B2 => n129, ZN 
                           => n179);
   U30 : AOI221_X1 port map( B1 => n66, B2 => n123, C1 => n70, C2 => n122, A =>
                           n140, ZN => n134);
   U31 : OAI22_X1 port map( A1 => n104, A2 => n118, B1 => n105, B2 => n128, ZN 
                           => n140);
   U32 : AOI221_X1 port map( B1 => n127, B2 => n123, C1 => n84, C2 => n122, A 
                           => n138, ZN => n113);
   U33 : OAI22_X1 port map( A1 => n104, A2 => n108, B1 => n105, B2 => n139, ZN 
                           => n138);
   U34 : OAI222_X1 port map( A1 => n242, A2 => n76, B1 => n104, B2 => n208, C1 
                           => n105, C2 => n80, ZN => n103);
   U35 : OAI222_X1 port map( A1 => n71, A2 => n105, B1 => n93, B2 => n104, C1 
                           => n90, C2 => n242, ZN => n178);
   U36 : OAI222_X1 port map( A1 => n61, A2 => n105, B1 => n206, B2 => n104, C1 
                           => n87, C2 => n242, ZN => n133);
   U37 : OAI222_X1 port map( A1 => n86, A2 => n105, B1 => n207, B2 => n104, C1 
                           => n81, C2 => n242, ZN => n112);
   U38 : OAI221_X1 port map( B1 => n90, B2 => n62, C1 => n91, C2 => n64, A => 
                           n92, ZN => B(4));
   U39 : AOI222_X1 port map( A1 => n244, A2 => n75, B1 => n67, B2 => n195, C1 
                           => n69, C2 => n204, ZN => n92);
   U40 : INV_X1 port map( A => n71, ZN => n195);
   U41 : OAI221_X1 port map( B1 => n87, B2 => n62, C1 => n88, C2 => n64, A => 
                           n89, ZN => B(5));
   U42 : AOI222_X1 port map( A1 => n244, A2 => n70, B1 => n67, B2 => n197, C1 
                           => n69, C2 => n68, ZN => n89);
   U43 : INV_X1 port map( A => n61, ZN => n197);
   U44 : OAI221_X1 port map( B1 => n81, B2 => n62, C1 => n82, C2 => n64, A => 
                           n83, ZN => B(6));
   U45 : AOI222_X1 port map( A1 => n244, A2 => n84, B1 => n67, B2 => n199, C1 
                           => n69, C2 => n85, ZN => n83);
   U46 : INV_X1 port map( A => n86, ZN => n199);
   U47 : OAI221_X1 port map( B1 => n76, B2 => n62, C1 => n220, C2 => n64, A => 
                           n77, ZN => B(7));
   U48 : AOI222_X1 port map( A1 => n244, A2 => n78, B1 => n67, B2 => n202, C1 
                           => n69, C2 => n79, ZN => n77);
   U49 : INV_X1 port map( A => n80, ZN => n202);
   U50 : OAI221_X1 port map( B1 => n71, B2 => n62, C1 => n72, C2 => n64, A => 
                           n73, ZN => B(8));
   U51 : AOI222_X1 port map( A1 => n244, A2 => n74, B1 => n67, B2 => n204, C1 
                           => n69, C2 => n75, ZN => n73);
   U52 : OAI221_X1 port map( B1 => n61, B2 => n62, C1 => n63, C2 => n64, A => 
                           n65, ZN => B(9));
   U53 : AOI222_X1 port map( A1 => n244, A2 => n66, B1 => n67, B2 => n68, C1 =>
                           n69, C2 => n70, ZN => n65);
   U54 : OAI221_X1 port map( B1 => n86, B2 => n62, C1 => n121, C2 => n64, A => 
                           n159, ZN => B(10));
   U55 : AOI222_X1 port map( A1 => n244, A2 => n127, B1 => n67, B2 => n85, C1 
                           => n69, C2 => n84, ZN => n159);
   U56 : NOR2_X1 port map( A1 => n64, A2 => n245, ZN => n144);
   U57 : OAI221_X1 port map( B1 => n129, B2 => n142, C1 => n93, C2 => n62, A =>
                           n151, ZN => B(12));
   U58 : AOI222_X1 port map( A1 => n69, A2 => n74, B1 => n144, B2 => n231, C1 
                           => n67, C2 => n75, ZN => n151);
   U59 : OAI221_X1 port map( B1 => n128, B2 => n142, C1 => n206, C2 => n62, A 
                           => n146, ZN => B(13));
   U60 : AOI222_X1 port map( A1 => n69, A2 => n66, B1 => n144, B2 => n233, C1 
                           => n67, C2 => n70, ZN => n146);
   U61 : OAI221_X1 port map( B1 => n139, B2 => n142, C1 => n207, C2 => n62, A 
                           => n145, ZN => B(14));
   U62 : AOI222_X1 port map( A1 => n69, A2 => n127, B1 => n144, B2 => n234, C1 
                           => n67, C2 => n84, ZN => n145);
   U63 : OAI221_X1 port map( B1 => n125, B2 => n142, C1 => n208, C2 => n62, A 
                           => n143, ZN => B(15));
   U64 : AOI222_X1 port map( A1 => n69, A2 => n219, B1 => n144, B2 => n235, C1 
                           => n67, C2 => n78, ZN => n143);
   U65 : INV_X1 port map( A => n107, ZN => n235);
   U66 : OAI22_X1 port map( A1 => n100, A2 => n191, B1 => n101, B2 => n192, ZN 
                           => n97);
   U67 : AOI22_X1 port map( A1 => n222, A2 => n122, B1 => n231, B2 => n123, ZN 
                           => n72);
   U68 : AOI22_X1 port map( A1 => n224, A2 => n122, B1 => n233, B2 => n123, ZN 
                           => n63);
   U69 : AOI22_X1 port map( A1 => n227, A2 => n122, B1 => n234, B2 => n123, ZN 
                           => n121);
   U70 : OAI22_X1 port map( A1 => n240, A2 => n189, B1 => n236, B2 => n190, ZN 
                           => n98);
   U71 : INV_X1 port map( A => n142, ZN => n244);
   U72 : INV_X1 port map( A => n123, ZN => n242);
   U73 : AND2_X1 port map( A1 => n161, A2 => n243, ZN => n69);
   U74 : INV_X1 port map( A => n122, ZN => n245);
   U75 : NOR2_X1 port map( A1 => n62, A2 => n107, ZN => B(31));
   U76 : NOR2_X1 port map( A1 => n119, A2 => n62, ZN => B(28));
   U77 : NOR2_X1 port map( A1 => n118, A2 => n62, ZN => B(29));
   U78 : NOR2_X1 port map( A1 => n108, A2 => n62, ZN => B(30));
   U79 : INV_X1 port map( A => n105, ZN => n241);
   U80 : INV_X1 port map( A => n118, ZN => n233);
   U82 : INV_X1 port map( A => n119, ZN => n231);
   U83 : INV_X1 port map( A => n108, ZN => n234);
   U84 : NOR2_X1 port map( A1 => n102, A2 => n246, ZN => B(19));
   U85 : INV_X1 port map( A => n93, ZN => n204);
   U86 : INV_X1 port map( A => n129, ZN => n222);
   U87 : INV_X1 port map( A => n128, ZN => n224);
   U88 : INV_X1 port map( A => n139, ZN => n227);
   U90 : INV_X1 port map( A => n126, ZN => n219);
   U91 : INV_X1 port map( A => n85, ZN => n207);
   U92 : INV_X1 port map( A => n79, ZN => n208);
   U93 : INV_X1 port map( A => n68, ZN => n206);
   U94 : INV_X1 port map( A => n124, ZN => n220);
   U95 : OAI222_X1 port map( A1 => n125, A2 => n242, B1 => n107, B2 => n105, C1
                           => n126, C2 => n245, ZN => n124);
   U96 : NOR2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n117);
   U97 : NOR2_X2 port map( A1 => n238, A2 => SH(1), ZN => n116);
   U98 : AOI222_X1 port map( A1 => n116, A2 => A(30), B1 => n237, B2 => A(31), 
                           C1 => n117, C2 => A(29), ZN => n118);
   U99 : AOI221_X1 port map( B1 => n239, B2 => A(26), C1 => n237, C2 => A(25), 
                           A => n158, ZN => n126);
   U100 : OAI22_X1 port map( A1 => n223, A2 => n236, B1 => n221, B2 => n240, ZN
                           => n158);
   U101 : AOI221_X1 port map( B1 => n239, B2 => A(28), C1 => n237, C2 => A(27),
                           A => n150, ZN => n128);
   U102 : OAI22_X1 port map( A1 => n226, A2 => n236, B1 => n225, B2 => n240, ZN
                           => n150);
   U103 : INV_X1 port map( A => A(26), ZN => n226);
   U104 : AOI221_X1 port map( B1 => n239, B2 => A(29), C1 => n237, C2 => A(28),
                           A => n228, ZN => n139);
   U105 : INV_X1 port map( A => n165, ZN => n228);
   U106 : AOI22_X1 port map( A1 => A(27), A2 => n116, B1 => A(26), B2 => n117, 
                           ZN => n165);
   U107 : AOI221_X1 port map( B1 => n239, B2 => A(27), C1 => n237, C2 => A(26),
                           A => n180, ZN => n129);
   U108 : OAI22_X1 port map( A1 => n225, A2 => n236, B1 => n223, B2 => n240, ZN
                           => n180);
   U109 : AOI221_X1 port map( B1 => n239, B2 => A(13), C1 => n237, C2 => A(12),
                           A => n166, ZN => n86);
   U110 : OAI22_X1 port map( A1 => n201, A2 => n236, B1 => n200, B2 => n240, ZN
                           => n166);
   U111 : INV_X1 port map( A => A(11), ZN => n201);
   U112 : AOI221_X1 port map( B1 => n239, B2 => A(11), C1 => n237, C2 => A(10),
                           A => n186, ZN => n71);
   U114 : OAI22_X1 port map( A1 => n198, A2 => n236, B1 => n196, B2 => n240, ZN
                           => n186);
   U115 : AOI221_X1 port map( B1 => n239, B2 => A(12), C1 => n237, C2 => A(11),
                           A => n136, ZN => n61);
   U116 : OAI22_X1 port map( A1 => n200, A2 => n236, B1 => n198, B2 => n240, ZN
                           => n136);
   U117 : AOI221_X1 port map( B1 => n239, B2 => A(31), C1 => n237, C2 => A(30),
                           A => n232, ZN => n119);
   U118 : INV_X1 port map( A => n181, ZN => n232);
   U119 : AOI22_X1 port map( A1 => A(29), A2 => n116, B1 => A(28), B2 => n117, 
                           ZN => n181);
   U120 : AOI221_X1 port map( B1 => n239, B2 => A(15), C1 => n237, C2 => A(14),
                           A => n205, ZN => n93);
   U121 : INV_X1 port map( A => n185, ZN => n205);
   U122 : AOI22_X1 port map( A1 => A(13), A2 => n116, B1 => A(12), B2 => n117, 
                           ZN => n185);
   U123 : AOI221_X1 port map( B1 => n239, B2 => A(14), C1 => n237, C2 => A(13),
                           A => n203, ZN => n80);
   U124 : INV_X1 port map( A => n157, ZN => n203);
   U125 : AOI22_X1 port map( A1 => A(12), A2 => n116, B1 => A(11), B2 => n117, 
                           ZN => n157);
   U126 : NAND2_X1 port map( A1 => SH(1), A2 => SH(0), ZN => n101);
   U127 : OAI221_X1 port map( B1 => n101, B2 => n216, C1 => n100, C2 => n215, A
                           => n147, ZN => n70);
   U128 : INV_X1 port map( A => A(19), ZN => n215);
   U129 : AOI22_X1 port map( A1 => A(18), A2 => n116, B1 => A(17), B2 => n117, 
                           ZN => n147);
   U130 : OAI221_X1 port map( B1 => n101, B2 => n217, C1 => n100, C2 => n216, A
                           => n160, ZN => n84);
   U131 : AOI22_X1 port map( A1 => A(19), A2 => n116, B1 => A(18), B2 => n117, 
                           ZN => n160);
   U132 : OAI221_X1 port map( B1 => n101, B2 => n218, C1 => n100, C2 => n217, A
                           => n156, ZN => n78);
   U133 : AOI22_X1 port map( A1 => A(20), A2 => n116, B1 => A(19), B2 => n117, 
                           ZN => n156);
   U134 : OAI221_X1 port map( B1 => n236, B2 => n212, C1 => n211, C2 => n240, A
                           => n182, ZN => n75);
   U135 : AOI22_X1 port map( A1 => A(19), A2 => n239, B1 => A(18), B2 => n237, 
                           ZN => n182);
   U136 : OAI221_X1 port map( B1 => n101, B2 => n225, C1 => n100, C2 => n223, A
                           => n164, ZN => n127);
   U137 : AOI22_X1 port map( A1 => A(23), A2 => n116, B1 => A(22), B2 => n117, 
                           ZN => n164);
   U138 : OAI221_X1 port map( B1 => n101, B2 => n221, C1 => n100, C2 => n218, A
                           => n183, ZN => n74);
   U139 : AOI22_X1 port map( A1 => A(21), A2 => n116, B1 => A(20), B2 => n117, 
                           ZN => n183);
   U140 : OAI221_X1 port map( B1 => n101, B2 => n223, C1 => n100, C2 => n221, A
                           => n148, ZN => n66);
   U141 : AOI22_X1 port map( A1 => A(22), A2 => n116, B1 => A(21), B2 => n117, 
                           ZN => n148);
   U142 : AOI221_X1 port map( B1 => n239, B2 => A(30), C1 => n237, C2 => A(29),
                           A => n230, ZN => n125);
   U143 : INV_X1 port map( A => n154, ZN => n230);
   U144 : AOI22_X1 port map( A1 => A(28), A2 => n116, B1 => A(27), B2 => n117, 
                           ZN => n154);
   U145 : NAND2_X1 port map( A1 => SH(1), A2 => n238, ZN => n100);
   U146 : AOI221_X1 port map( B1 => n239, B2 => A(7), C1 => n237, C2 => A(6), A
                           => n184, ZN => n90);
   U147 : OAI22_X1 port map( A1 => n191, A2 => n236, B1 => n190, B2 => n240, ZN
                           => n184);
   U148 : AOI221_X1 port map( B1 => n239, B2 => A(8), C1 => n237, C2 => A(7), A
                           => n135, ZN => n87);
   U149 : OAI22_X1 port map( A1 => n192, A2 => n236, B1 => n191, B2 => n240, ZN
                           => n135);
   U150 : AOI221_X1 port map( B1 => n239, B2 => A(9), C1 => n237, C2 => A(8), A
                           => n114, ZN => n81);
   U152 : OAI22_X1 port map( A1 => n194, A2 => n236, B1 => n192, B2 => n240, ZN
                           => n114);
   U153 : OAI221_X1 port map( B1 => n101, B2 => n211, C1 => n100, C2 => n209, A
                           => n149, ZN => n68);
   U154 : AOI22_X1 port map( A1 => A(14), A2 => n116, B1 => A(13), B2 => n117, 
                           ZN => n149);
   U155 : OAI221_X1 port map( B1 => n101, B2 => n212, C1 => n211, C2 => n100, A
                           => n162, ZN => n85);
   U156 : AOI22_X1 port map( A1 => n116, A2 => A(15), B1 => n117, B2 => A(14), 
                           ZN => n162);
   U157 : OAI221_X1 port map( B1 => n211, B2 => n236, C1 => n209, C2 => n240, A
                           => n155, ZN => n79);
   U158 : AOI22_X1 port map( A1 => A(18), A2 => n239, B1 => A(17), B2 => n237, 
                           ZN => n155);
   U159 : AOI221_X1 port map( B1 => n239, B2 => A(10), C1 => n237, C2 => A(9), 
                           A => n106, ZN => n76);
   U160 : OAI22_X1 port map( A1 => n196, A2 => n236, B1 => n194, B2 => n240, ZN
                           => n106);
   U161 : AOI222_X1 port map( A1 => n78, A2 => n122, B1 => n219, B2 => n123, C1
                           => n229, C2 => SH(3), ZN => n102);
   U162 : INV_X1 port map( A => n120, ZN => n229);
   U163 : NOR4_X1 port map( A1 => n172, A2 => SH(29), A3 => SH(5), A4 => SH(30)
                           , ZN => n171);
   U164 : OR4_X1 port map( A1 => SH(7), A2 => SH(6), A3 => SH(9), A4 => SH(8), 
                           ZN => n172);
   U165 : NAND4_X1 port map( A1 => n168, A2 => n169, A3 => n170, A4 => n171, ZN
                           => n96);
   U166 : NOR4_X1 port map( A1 => n175, A2 => SH(10), A3 => SH(12), A4 => 
                           SH(11), ZN => n168);
   U167 : NOR4_X1 port map( A1 => n174, A2 => SH(16), A3 => SH(18), A4 => 
                           SH(17), ZN => n169);
   U168 : NOR4_X1 port map( A1 => n173, A2 => SH(23), A3 => SH(25), A4 => 
                           SH(24), ZN => n170);
   U169 : NAND2_X1 port map( A1 => SH(3), A2 => n243, ZN => n105);
   U170 : NAND2_X1 port map( A1 => SH(4), A2 => n247, ZN => n64);
   U171 : INV_X1 port map( A => n96, ZN => n247);
   U172 : AOI22_X1 port map( A1 => n117, A2 => A(30), B1 => n116, B2 => A(31), 
                           ZN => n108);
   U173 : NOR2_X1 port map( A1 => n245, A2 => SH(4), ZN => n99);
   U174 : NAND2_X1 port map( A1 => SH(3), A2 => SH(2), ZN => n104);
   U175 : OAI221_X1 port map( B1 => n126, B2 => n142, C1 => n80, C2 => n62, A 
                           => n152, ZN => B(11));
   U176 : AOI221_X1 port map( B1 => n69, B2 => n78, C1 => n67, C2 => n79, A => 
                           n153, ZN => n152);
   U177 : NOR3_X1 port map( A1 => n64, A2 => SH(3), A3 => n120, ZN => n153);
   U178 : NOR2_X1 port map( A1 => n96, A2 => SH(4), ZN => n163);
   U179 : NAND2_X1 port map( A1 => n161, A2 => SH(2), ZN => n142);
   U180 : NOR3_X1 port map( A1 => n246, A2 => SH(3), A3 => n120, ZN => B(27));
   U181 : AOI22_X1 port map( A1 => A(1), A2 => n116, B1 => A(0), B2 => n117, ZN
                           => n187);
   U182 : AOI22_X1 port map( A1 => A(2), A2 => n116, B1 => A(1), B2 => n117, ZN
                           => n137);
   U183 : AOI22_X1 port map( A1 => A(3), A2 => n116, B1 => A(2), B2 => n117, ZN
                           => n115);
   U184 : NAND2_X1 port map( A1 => A(31), A2 => n117, ZN => n107);
   U185 : AOI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => B(3));
   U186 : OAI21_X1 port map( B1 => n97, B2 => n98, A => n99, ZN => n95);
   U187 : INV_X1 port map( A => n103, ZN => n193);
   U188 : NOR2_X1 port map( A1 => n167, A2 => n96, ZN => B(0));
   U189 : AOI21_X1 port map( B1 => n99, B2 => n176, A => n177, ZN => n167);
   U190 : OAI221_X1 port map( B1 => n101, B2 => n189, C1 => n100, C2 => n188, A
                           => n187, ZN => n176);
   U191 : NOR2_X1 port map( A1 => n130, A2 => n96, ZN => B(1));
   U192 : AOI21_X1 port map( B1 => n99, B2 => n131, A => n132, ZN => n130);
   U193 : OAI221_X1 port map( B1 => n101, B2 => n190, C1 => n100, C2 => n189, A
                           => n137, ZN => n131);
   U194 : NOR2_X1 port map( A1 => n109, A2 => n96, ZN => B(2));
   U196 : AOI21_X1 port map( B1 => n99, B2 => n110, A => n111, ZN => n109);
   U197 : OAI221_X1 port map( B1 => n101, B2 => n191, C1 => n100, C2 => n190, A
                           => n115, ZN => n110);
   U198 : INV_X1 port map( A => A(4), ZN => n190);
   U199 : INV_X1 port map( A => A(5), ZN => n191);
   U200 : INV_X1 port map( A => A(24), ZN => n223);
   U201 : INV_X1 port map( A => A(16), ZN => n211);
   U202 : INV_X1 port map( A => SH(2), ZN => n243);
   U203 : INV_X1 port map( A => SH(0), ZN => n238);
   U204 : OR4_X1 port map( A1 => SH(20), A2 => SH(19), A3 => SH(22), A4 => 
                           SH(21), ZN => n174);
   U205 : INV_X1 port map( A => A(3), ZN => n189);
   U206 : INV_X1 port map( A => A(23), ZN => n221);
   U207 : INV_X1 port map( A => A(6), ZN => n192);
   U208 : INV_X1 port map( A => A(25), ZN => n225);
   U209 : INV_X1 port map( A => A(20), ZN => n216);
   U210 : INV_X1 port map( A => A(21), ZN => n217);
   U211 : INV_X1 port map( A => A(22), ZN => n218);
   U212 : INV_X1 port map( A => A(15), ZN => n209);
   U213 : INV_X1 port map( A => A(17), ZN => n212);
   U214 : INV_X1 port map( A => A(10), ZN => n200);
   U215 : INV_X1 port map( A => A(7), ZN => n194);
   U216 : INV_X1 port map( A => A(8), ZN => n196);
   U217 : INV_X1 port map( A => A(9), ZN => n198);
   U218 : AND2_X1 port map( A1 => SH(3), A2 => n163, ZN => n161);
   U219 : INV_X1 port map( A => A(2), ZN => n188);
   U220 : OR3_X1 port map( A1 => SH(28), A2 => SH(27), A3 => SH(26), ZN => n173
                           );
   U221 : OR3_X1 port map( A1 => SH(15), A2 => SH(14), A3 => SH(13), ZN => n175
                           );

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4 is

   port( A, B : in std_logic_vector (32 downto 1);  C0 : in std_logic;  COUT : 
         out std_logic_vector (8 downto 0));

end CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4;

architecture SYN_STRUCTURAL of CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_1
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_2
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_3
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_4
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_1
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_2
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_5
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_6
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_3
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_4
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_5
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_7
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_6
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_7
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_8
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_9
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_10
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_11
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_12
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_8
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_13
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_14
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_15
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_16
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_17
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_18
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_19
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_20
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_21
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_22
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_23
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_24
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_25
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_26
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_0
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_0
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component pg_generator_1
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_2
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_3
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_4
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_5
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_6
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_7
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_8
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_9
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_10
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_11
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_12
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_13
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_14
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_15
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_16
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_17
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_18
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_19
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_20
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_21
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_22
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_23
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_24
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_25
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_26
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_27
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_28
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_29
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_30
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_31
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_0
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   signal COUT_8_port, COUT_7_port, COUT_6_port, COUT_5_port, COUT_4_port, 
      COUT_3_port, COUT_2_port, COUT_1_port, gi_1_port, pi_1_port, 
      gSignal_16_16_port, gSignal_16_15_port, gSignal_16_13_port, 
      gSignal_16_9_port, gSignal_15_15_port, gSignal_14_14_port, 
      gSignal_14_13_port, gSignal_13_13_port, gSignal_12_12_port, 
      gSignal_12_11_port, gSignal_12_9_port, gSignal_11_11_port, 
      gSignal_10_10_port, gSignal_10_9_port, gSignal_9_9_port, gSignal_8_8_port
      , gSignal_8_7_port, gSignal_8_5_port, gSignal_7_7_port, gSignal_6_6_port,
      gSignal_6_5_port, gSignal_5_5_port, gSignal_4_4_port, gSignal_4_3_port, 
      gSignal_3_3_port, gSignal_2_2_port, gSignal_2_1_port, pSignal_16_16_port,
      pSignal_16_15_port, pSignal_16_13_port, pSignal_16_9_port, 
      pSignal_15_15_port, pSignal_14_14_port, pSignal_14_13_port, 
      pSignal_13_13_port, pSignal_12_12_port, pSignal_12_11_port, 
      pSignal_12_9_port, pSignal_11_11_port, pSignal_10_10_port, 
      pSignal_10_9_port, pSignal_9_9_port, pSignal_8_8_port, pSignal_8_7_port, 
      pSignal_8_5_port, pSignal_7_7_port, pSignal_6_6_port, pSignal_6_5_port, 
      pSignal_5_5_port, pSignal_4_4_port, pSignal_4_3_port, pSignal_3_3_port, 
      pSignal_2_2_port, pSignal_32_32_port, pSignal_32_31_port, 
      pSignal_32_29_port, pSignal_32_25_port, pSignal_32_17_port, 
      pSignal_31_31_port, pSignal_30_30_port, pSignal_30_29_port, 
      pSignal_29_29_port, pSignal_28_28_port, pSignal_28_27_port, 
      pSignal_28_25_port, pSignal_28_17_port, pSignal_27_27_port, 
      pSignal_26_26_port, pSignal_26_25_port, pSignal_25_25_port, 
      pSignal_24_24_port, pSignal_24_23_port, pSignal_24_21_port, 
      pSignal_24_17_port, pSignal_23_23_port, pSignal_22_22_port, 
      pSignal_22_21_port, pSignal_21_21_port, pSignal_20_20_port, 
      pSignal_20_19_port, pSignal_20_17_port, pSignal_19_19_port, 
      pSignal_18_18_port, pSignal_18_17_port, pSignal_17_17_port, 
      gSignal_32_32_port, gSignal_32_31_port, gSignal_32_29_port, 
      gSignal_32_25_port, gSignal_32_17_port, gSignal_31_31_port, 
      gSignal_30_30_port, gSignal_30_29_port, gSignal_29_29_port, 
      gSignal_28_28_port, gSignal_28_27_port, gSignal_28_25_port, 
      gSignal_28_17_port, gSignal_27_27_port, gSignal_26_26_port, 
      gSignal_26_25_port, gSignal_25_25_port, gSignal_24_24_port, 
      gSignal_24_23_port, gSignal_24_21_port, gSignal_24_17_port, 
      gSignal_23_23_port, gSignal_22_22_port, gSignal_22_21_port, 
      gSignal_21_21_port, gSignal_20_20_port, gSignal_20_19_port, 
      gSignal_20_17_port, gSignal_19_19_port, gSignal_18_18_port, 
      gSignal_18_17_port, gSignal_17_17_port, n2, n3 : std_logic;

begin
   COUT <= ( COUT_8_port, COUT_7_port, COUT_6_port, COUT_5_port, COUT_4_port, 
      COUT_3_port, COUT_2_port, COUT_1_port, C0 );
   
   pg_inst_1 : pg_generator_0 port map( A => A(1), B => B(1), P => pi_1_port, G
                           => gi_1_port);
   pg_inst_2 : pg_generator_31 port map( A => A(2), B => B(2), P => 
                           pSignal_2_2_port, G => gSignal_2_2_port);
   pg_inst_3 : pg_generator_30 port map( A => A(3), B => B(3), P => 
                           pSignal_3_3_port, G => gSignal_3_3_port);
   pg_inst_4 : pg_generator_29 port map( A => A(4), B => B(4), P => 
                           pSignal_4_4_port, G => gSignal_4_4_port);
   pg_inst_5 : pg_generator_28 port map( A => A(5), B => B(5), P => 
                           pSignal_5_5_port, G => gSignal_5_5_port);
   pg_inst_6 : pg_generator_27 port map( A => A(6), B => B(6), P => 
                           pSignal_6_6_port, G => gSignal_6_6_port);
   pg_inst_7 : pg_generator_26 port map( A => A(7), B => B(7), P => 
                           pSignal_7_7_port, G => gSignal_7_7_port);
   pg_inst_8 : pg_generator_25 port map( A => A(8), B => B(8), P => 
                           pSignal_8_8_port, G => gSignal_8_8_port);
   pg_inst_9 : pg_generator_24 port map( A => A(9), B => B(9), P => 
                           pSignal_9_9_port, G => gSignal_9_9_port);
   pg_inst_10 : pg_generator_23 port map( A => A(10), B => B(10), P => 
                           pSignal_10_10_port, G => gSignal_10_10_port);
   pg_inst_11 : pg_generator_22 port map( A => A(11), B => B(11), P => 
                           pSignal_11_11_port, G => gSignal_11_11_port);
   pg_inst_12 : pg_generator_21 port map( A => A(12), B => B(12), P => 
                           pSignal_12_12_port, G => gSignal_12_12_port);
   pg_inst_13 : pg_generator_20 port map( A => A(13), B => B(13), P => 
                           pSignal_13_13_port, G => gSignal_13_13_port);
   pg_inst_14 : pg_generator_19 port map( A => A(14), B => B(14), P => 
                           pSignal_14_14_port, G => gSignal_14_14_port);
   pg_inst_15 : pg_generator_18 port map( A => A(15), B => B(15), P => 
                           pSignal_15_15_port, G => gSignal_15_15_port);
   pg_inst_16 : pg_generator_17 port map( A => A(16), B => B(16), P => 
                           pSignal_16_16_port, G => gSignal_16_16_port);
   pg_inst_17 : pg_generator_16 port map( A => A(17), B => B(17), P => 
                           pSignal_17_17_port, G => gSignal_17_17_port);
   pg_inst_18 : pg_generator_15 port map( A => A(18), B => B(18), P => 
                           pSignal_18_18_port, G => gSignal_18_18_port);
   pg_inst_19 : pg_generator_14 port map( A => A(19), B => B(19), P => 
                           pSignal_19_19_port, G => gSignal_19_19_port);
   pg_inst_20 : pg_generator_13 port map( A => A(20), B => B(20), P => 
                           pSignal_20_20_port, G => gSignal_20_20_port);
   pg_inst_21 : pg_generator_12 port map( A => A(21), B => B(21), P => 
                           pSignal_21_21_port, G => gSignal_21_21_port);
   pg_inst_22 : pg_generator_11 port map( A => A(22), B => B(22), P => 
                           pSignal_22_22_port, G => gSignal_22_22_port);
   pg_inst_23 : pg_generator_10 port map( A => A(23), B => B(23), P => 
                           pSignal_23_23_port, G => gSignal_23_23_port);
   pg_inst_24 : pg_generator_9 port map( A => A(24), B => B(24), P => 
                           pSignal_24_24_port, G => gSignal_24_24_port);
   pg_inst_25 : pg_generator_8 port map( A => A(25), B => B(25), P => 
                           pSignal_25_25_port, G => gSignal_25_25_port);
   pg_inst_26 : pg_generator_7 port map( A => A(26), B => B(26), P => 
                           pSignal_26_26_port, G => gSignal_26_26_port);
   pg_inst_27 : pg_generator_6 port map( A => A(27), B => B(27), P => 
                           pSignal_27_27_port, G => gSignal_27_27_port);
   pg_inst_28 : pg_generator_5 port map( A => A(28), B => B(28), P => 
                           pSignal_28_28_port, G => gSignal_28_28_port);
   pg_inst_29 : pg_generator_4 port map( A => A(29), B => B(29), P => 
                           pSignal_29_29_port, G => gSignal_29_29_port);
   pg_inst_30 : pg_generator_3 port map( A => A(30), B => B(30), P => 
                           pSignal_30_30_port, G => gSignal_30_30_port);
   pg_inst_31 : pg_generator_2 port map( A => A(31), B => B(31), P => 
                           pSignal_31_31_port, G => gSignal_31_31_port);
   pg_inst_32 : pg_generator_1 port map( A => A(32), B => B(32), P => 
                           pSignal_32_32_port, G => gSignal_32_32_port);
   G1_1_2 : G_0 port map( p_ik => pSignal_2_2_port, g_ik => gSignal_2_2_port, 
                           g_k1j => n3, G_ij => gSignal_2_1_port);
   PG_inst1_1_4 : PG_0 port map( p_ik => pSignal_4_4_port, g_ik => 
                           gSignal_4_4_port, p_k1j => pSignal_3_3_port, g_k1j 
                           => gSignal_3_3_port, P_ij => pSignal_4_3_port, G_ij 
                           => gSignal_4_3_port);
   PG_inst1_1_6 : PG_26 port map( p_ik => pSignal_6_6_port, g_ik => 
                           gSignal_6_6_port, p_k1j => pSignal_5_5_port, g_k1j 
                           => gSignal_5_5_port, P_ij => pSignal_6_5_port, G_ij 
                           => gSignal_6_5_port);
   PG_inst1_1_8 : PG_25 port map( p_ik => pSignal_8_8_port, g_ik => 
                           gSignal_8_8_port, p_k1j => pSignal_7_7_port, g_k1j 
                           => gSignal_7_7_port, P_ij => pSignal_8_7_port, G_ij 
                           => gSignal_8_7_port);
   PG_inst1_1_10 : PG_24 port map( p_ik => pSignal_10_10_port, g_ik => 
                           gSignal_10_10_port, p_k1j => pSignal_9_9_port, g_k1j
                           => gSignal_9_9_port, P_ij => pSignal_10_9_port, G_ij
                           => gSignal_10_9_port);
   PG_inst1_1_12 : PG_23 port map( p_ik => pSignal_12_12_port, g_ik => 
                           gSignal_12_12_port, p_k1j => pSignal_11_11_port, 
                           g_k1j => gSignal_11_11_port, P_ij => 
                           pSignal_12_11_port, G_ij => gSignal_12_11_port);
   PG_inst1_1_14 : PG_22 port map( p_ik => pSignal_14_14_port, g_ik => 
                           gSignal_14_14_port, p_k1j => pSignal_13_13_port, 
                           g_k1j => gSignal_13_13_port, P_ij => 
                           pSignal_14_13_port, G_ij => gSignal_14_13_port);
   PG_inst1_1_16 : PG_21 port map( p_ik => pSignal_16_16_port, g_ik => 
                           gSignal_16_16_port, p_k1j => pSignal_15_15_port, 
                           g_k1j => gSignal_15_15_port, P_ij => 
                           pSignal_16_15_port, G_ij => gSignal_16_15_port);
   PG_inst1_1_18 : PG_20 port map( p_ik => pSignal_18_18_port, g_ik => 
                           gSignal_18_18_port, p_k1j => pSignal_17_17_port, 
                           g_k1j => gSignal_17_17_port, P_ij => 
                           pSignal_18_17_port, G_ij => gSignal_18_17_port);
   PG_inst1_1_20 : PG_19 port map( p_ik => pSignal_20_20_port, g_ik => 
                           gSignal_20_20_port, p_k1j => pSignal_19_19_port, 
                           g_k1j => gSignal_19_19_port, P_ij => 
                           pSignal_20_19_port, G_ij => gSignal_20_19_port);
   PG_inst1_1_22 : PG_18 port map( p_ik => pSignal_22_22_port, g_ik => 
                           gSignal_22_22_port, p_k1j => pSignal_21_21_port, 
                           g_k1j => gSignal_21_21_port, P_ij => 
                           pSignal_22_21_port, G_ij => gSignal_22_21_port);
   PG_inst1_1_24 : PG_17 port map( p_ik => pSignal_24_24_port, g_ik => 
                           gSignal_24_24_port, p_k1j => pSignal_23_23_port, 
                           g_k1j => gSignal_23_23_port, P_ij => 
                           pSignal_24_23_port, G_ij => gSignal_24_23_port);
   PG_inst1_1_26 : PG_16 port map( p_ik => pSignal_26_26_port, g_ik => 
                           gSignal_26_26_port, p_k1j => pSignal_25_25_port, 
                           g_k1j => gSignal_25_25_port, P_ij => 
                           pSignal_26_25_port, G_ij => gSignal_26_25_port);
   PG_inst1_1_28 : PG_15 port map( p_ik => pSignal_28_28_port, g_ik => 
                           gSignal_28_28_port, p_k1j => pSignal_27_27_port, 
                           g_k1j => gSignal_27_27_port, P_ij => 
                           pSignal_28_27_port, G_ij => gSignal_28_27_port);
   PG_inst1_1_30 : PG_14 port map( p_ik => pSignal_30_30_port, g_ik => 
                           gSignal_30_30_port, p_k1j => pSignal_29_29_port, 
                           g_k1j => gSignal_29_29_port, P_ij => 
                           pSignal_30_29_port, G_ij => gSignal_30_29_port);
   PG_inst1_1_32 : PG_13 port map( p_ik => pSignal_32_32_port, g_ik => 
                           gSignal_32_32_port, p_k1j => pSignal_31_31_port, 
                           g_k1j => gSignal_31_31_port, P_ij => 
                           pSignal_32_31_port, G_ij => gSignal_32_31_port);
   G1_2_4 : G_8 port map( p_ik => pSignal_4_3_port, g_ik => gSignal_4_3_port, 
                           g_k1j => gSignal_2_1_port, G_ij => COUT_1_port);
   PG_inst1_2_8 : PG_12 port map( p_ik => pSignal_8_7_port, g_ik => 
                           gSignal_8_7_port, p_k1j => pSignal_6_5_port, g_k1j 
                           => gSignal_6_5_port, P_ij => pSignal_8_5_port, G_ij 
                           => gSignal_8_5_port);
   PG_inst1_2_12 : PG_11 port map( p_ik => pSignal_12_11_port, g_ik => 
                           gSignal_12_11_port, p_k1j => pSignal_10_9_port, 
                           g_k1j => gSignal_10_9_port, P_ij => 
                           pSignal_12_9_port, G_ij => gSignal_12_9_port);
   PG_inst1_2_16 : PG_10 port map( p_ik => pSignal_16_15_port, g_ik => 
                           gSignal_16_15_port, p_k1j => pSignal_14_13_port, 
                           g_k1j => gSignal_14_13_port, P_ij => 
                           pSignal_16_13_port, G_ij => gSignal_16_13_port);
   PG_inst1_2_20 : PG_9 port map( p_ik => pSignal_20_19_port, g_ik => 
                           gSignal_20_19_port, p_k1j => pSignal_18_17_port, 
                           g_k1j => gSignal_18_17_port, P_ij => 
                           pSignal_20_17_port, G_ij => gSignal_20_17_port);
   PG_inst1_2_24 : PG_8 port map( p_ik => pSignal_24_23_port, g_ik => 
                           gSignal_24_23_port, p_k1j => pSignal_22_21_port, 
                           g_k1j => gSignal_22_21_port, P_ij => 
                           pSignal_24_21_port, G_ij => gSignal_24_21_port);
   PG_inst1_2_28 : PG_7 port map( p_ik => pSignal_28_27_port, g_ik => 
                           gSignal_28_27_port, p_k1j => pSignal_26_25_port, 
                           g_k1j => gSignal_26_25_port, P_ij => 
                           pSignal_28_25_port, G_ij => gSignal_28_25_port);
   PG_inst1_2_32 : PG_6 port map( p_ik => pSignal_32_31_port, g_ik => 
                           gSignal_32_31_port, p_k1j => pSignal_30_29_port, 
                           g_k1j => gSignal_30_29_port, P_ij => 
                           pSignal_32_29_port, G_ij => gSignal_32_29_port);
   G_INST2_0_4_8 : G_7 port map( p_ik => pSignal_8_5_port, g_ik => 
                           gSignal_8_5_port, g_k1j => COUT_1_port, G_ij => 
                           COUT_2_port);
   PG_INST2_0_12_16 : PG_5 port map( p_ik => pSignal_16_13_port, g_ik => 
                           gSignal_16_13_port, p_k1j => pSignal_12_9_port, 
                           g_k1j => gSignal_12_9_port, P_ij => 
                           pSignal_16_9_port, G_ij => gSignal_16_9_port);
   PG_INST2_0_20_24 : PG_4 port map( p_ik => pSignal_24_21_port, g_ik => 
                           gSignal_24_21_port, p_k1j => pSignal_20_17_port, 
                           g_k1j => gSignal_20_17_port, P_ij => 
                           pSignal_24_17_port, G_ij => gSignal_24_17_port);
   PG_INST2_0_28_32 : PG_3 port map( p_ik => pSignal_32_29_port, g_ik => 
                           gSignal_32_29_port, p_k1j => pSignal_28_25_port, 
                           g_k1j => gSignal_28_25_port, P_ij => 
                           pSignal_32_25_port, G_ij => gSignal_32_25_port);
   G_INST2_1_8_12 : G_6 port map( p_ik => pSignal_12_9_port, g_ik => 
                           gSignal_12_9_port, g_k1j => COUT_2_port, G_ij => 
                           COUT_3_port);
   G_INST2_1_8_16 : G_5 port map( p_ik => pSignal_16_9_port, g_ik => 
                           gSignal_16_9_port, g_k1j => COUT_2_port, G_ij => 
                           COUT_4_port);
   PG_INST2_1_24_28 : PG_2 port map( p_ik => pSignal_28_25_port, g_ik => 
                           gSignal_28_25_port, p_k1j => pSignal_24_17_port, 
                           g_k1j => gSignal_24_17_port, P_ij => 
                           pSignal_28_17_port, G_ij => gSignal_28_17_port);
   PG_INST2_1_24_32 : PG_1 port map( p_ik => pSignal_32_25_port, g_ik => 
                           gSignal_32_25_port, p_k1j => pSignal_24_17_port, 
                           g_k1j => gSignal_24_17_port, P_ij => 
                           pSignal_32_17_port, G_ij => gSignal_32_17_port);
   G_INST2_2_16_20 : G_4 port map( p_ik => pSignal_20_17_port, g_ik => 
                           gSignal_20_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_5_port);
   G_INST2_2_16_24 : G_3 port map( p_ik => pSignal_24_17_port, g_ik => 
                           gSignal_24_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_6_port);
   G_INST2_2_16_28 : G_2 port map( p_ik => pSignal_28_17_port, g_ik => 
                           gSignal_28_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_7_port);
   G_INST2_2_16_32 : G_1 port map( p_ik => pSignal_32_17_port, g_ik => 
                           gSignal_32_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_8_port);
   U1 : INV_X1 port map( A => n2, ZN => n3);
   U2 : AOI21_X1 port map( B1 => pi_1_port, B2 => C0, A => gi_1_port, ZN => n2)
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (8
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8;

architecture SYN_STRUCTURAL of 
   SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8 is

   component CarrySelect_1
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_2
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_3
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_4
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_5
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_6
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_7
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_0
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   carrySel_0 : CarrySelect_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Cin => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   carrySel_1 : CarrySelect_7 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Cin => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   carrySel_2 : CarrySelect_6 port map( A(3) => A(11), A(2) => A(10), A(1) => 
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Cin => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   carrySel_3 : CarrySelect_5 port map( A(3) => A(15), A(2) => A(14), A(1) => 
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Cin => Ci(3), S(3) => 
                           S(15), S(2) => S(14), S(1) => S(13), S(0) => S(12));
   carrySel_4 : CarrySelect_4 port map( A(3) => A(19), A(2) => A(18), A(1) => 
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Cin => Ci(4), S(3) => 
                           S(19), S(2) => S(18), S(1) => S(17), S(0) => S(16));
   carrySel_5 : CarrySelect_3 port map( A(3) => A(23), A(2) => A(22), A(1) => 
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Cin => Ci(5), S(3) => 
                           S(23), S(2) => S(22), S(1) => S(21), S(0) => S(20));
   carrySel_6 : CarrySelect_2 port map( A(3) => A(27), A(2) => A(26), A(1) => 
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Cin => Ci(6), S(3) => 
                           S(27), S(2) => S(26), S(1) => S(25), S(0) => S(24));
   carrySel_7 : CarrySelect_1 port map( A(3) => A(31), A(2) => A(30), A(1) => 
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Cin => Ci(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_logic_nbits32 is

   port( Cin : in std_logic;  B0 : in std_logic_vector (31 downto 0);  B : out 
         std_logic_vector (31 downto 0));

end xor_logic_nbits32;

architecture SYN_BEHAVIORAL of xor_logic_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n1, B => B0(9), Z => B(9));
   U2 : XOR2_X1 port map( A => n1, B => B0(8), Z => B(8));
   U3 : XOR2_X1 port map( A => n1, B => B0(7), Z => B(7));
   U4 : XOR2_X1 port map( A => n1, B => B0(6), Z => B(6));
   U5 : XOR2_X1 port map( A => n1, B => B0(5), Z => B(5));
   U6 : XOR2_X1 port map( A => n1, B => B0(4), Z => B(4));
   U7 : XOR2_X1 port map( A => n1, B => B0(3), Z => B(3));
   U8 : XOR2_X1 port map( A => n1, B => B0(31), Z => B(31));
   U9 : XOR2_X1 port map( A => n1, B => B0(30), Z => B(30));
   U10 : XOR2_X1 port map( A => n1, B => B0(2), Z => B(2));
   U11 : XOR2_X1 port map( A => n1, B => B0(29), Z => B(29));
   U12 : XOR2_X1 port map( A => n1, B => B0(28), Z => B(28));
   U13 : XOR2_X1 port map( A => n2, B => B0(27), Z => B(27));
   U14 : XOR2_X1 port map( A => n2, B => B0(26), Z => B(26));
   U15 : XOR2_X1 port map( A => n2, B => B0(25), Z => B(25));
   U16 : XOR2_X1 port map( A => n2, B => B0(24), Z => B(24));
   U17 : XOR2_X1 port map( A => n2, B => B0(23), Z => B(23));
   U18 : XOR2_X1 port map( A => n2, B => B0(22), Z => B(22));
   U19 : XOR2_X1 port map( A => n2, B => B0(21), Z => B(21));
   U20 : XOR2_X1 port map( A => n2, B => B0(20), Z => B(20));
   U21 : XOR2_X1 port map( A => n2, B => B0(1), Z => B(1));
   U22 : XOR2_X1 port map( A => n2, B => B0(19), Z => B(19));
   U23 : XOR2_X1 port map( A => n2, B => B0(18), Z => B(18));
   U24 : XOR2_X1 port map( A => n2, B => B0(17), Z => B(17));
   U25 : XOR2_X1 port map( A => n3, B => B0(16), Z => B(16));
   U26 : XOR2_X1 port map( A => n3, B => B0(15), Z => B(15));
   U27 : XOR2_X1 port map( A => n3, B => B0(14), Z => B(14));
   U28 : XOR2_X1 port map( A => n3, B => B0(13), Z => B(13));
   U29 : XOR2_X1 port map( A => n3, B => B0(12), Z => B(12));
   U30 : XOR2_X1 port map( A => n3, B => B0(11), Z => B(11));
   U31 : XOR2_X1 port map( A => n3, B => B0(10), Z => B(10));
   U32 : XOR2_X1 port map( A => n3, B => B0(0), Z => B(0));
   U33 : BUF_X1 port map( A => Cin, Z => n4);
   U34 : BUF_X1 port map( A => n4, Z => n3);
   U35 : BUF_X1 port map( A => n4, Z => n1);
   U36 : BUF_X1 port map( A => n4, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity logic_and_shift_N32 is

   port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
         downto 0));

end logic_and_shift_N32;

architecture SYN_BEHAVIOR of logic_and_shift_N32 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component logic_and_shift_N32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component logic_and_shift_N32_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,
      N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57
      , N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, 
      N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86
      , N87, N88, N89, N90, N91, N92, N190, N191, N192, N193, N194, N195, N196,
      N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, 
      N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, 
      N221, n3, n4, n71_port, n73_port, n74_port, n75_port, n76_port, n77_port,
      n78_port, n80_port, n81_port, n82_port, n83_port, n84_port, n85_port, 
      n86_port, n87_port, n88_port, n89_port, n90_port, n91_port, n92_port, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n207_port, n208_port, n209_port
      , n210_port, n211_port, n212_port, n213_port, n214_port, n215_port, 
      n216_port, n217_port, n218_port, n219_port, n220_port, n221_port, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305 : 
      std_logic;

begin
   
   OUTALU_reg_31_inst : DLH_X1 port map( G => n211_port, D => N221, Q => 
                           OUTALU(31));
   OUTALU_reg_30_inst : DLH_X1 port map( G => n211_port, D => N220, Q => 
                           OUTALU(30));
   OUTALU_reg_29_inst : DLH_X1 port map( G => n209_port, D => N219, Q => 
                           OUTALU(29));
   OUTALU_reg_28_inst : DLH_X1 port map( G => n211_port, D => N218, Q => 
                           OUTALU(28));
   OUTALU_reg_27_inst : DLH_X1 port map( G => n211_port, D => N217, Q => 
                           OUTALU(27));
   OUTALU_reg_26_inst : DLH_X1 port map( G => n211_port, D => N216, Q => 
                           OUTALU(26));
   OUTALU_reg_25_inst : DLH_X1 port map( G => n209_port, D => N215, Q => 
                           OUTALU(25));
   OUTALU_reg_24_inst : DLH_X1 port map( G => n210_port, D => N214, Q => 
                           OUTALU(24));
   OUTALU_reg_23_inst : DLH_X1 port map( G => n210_port, D => N213, Q => 
                           OUTALU(23));
   OUTALU_reg_22_inst : DLH_X1 port map( G => n210_port, D => N212, Q => 
                           OUTALU(22));
   OUTALU_reg_21_inst : DLH_X1 port map( G => n209_port, D => N211, Q => 
                           OUTALU(21));
   OUTALU_reg_20_inst : DLH_X1 port map( G => n210_port, D => N210, Q => 
                           OUTALU(20));
   OUTALU_reg_19_inst : DLH_X1 port map( G => n209_port, D => N209, Q => 
                           OUTALU(19));
   OUTALU_reg_18_inst : DLH_X1 port map( G => n210_port, D => N208, Q => 
                           OUTALU(18));
   OUTALU_reg_17_inst : DLH_X1 port map( G => n209_port, D => N207, Q => 
                           OUTALU(17));
   OUTALU_reg_16_inst : DLH_X1 port map( G => n211_port, D => N206, Q => 
                           OUTALU(16));
   OUTALU_reg_15_inst : DLH_X1 port map( G => n209_port, D => N205, Q => 
                           OUTALU(15));
   OUTALU_reg_14_inst : DLH_X1 port map( G => n210_port, D => N204, Q => 
                           OUTALU(14));
   OUTALU_reg_13_inst : DLH_X1 port map( G => n209_port, D => N203, Q => 
                           OUTALU(13));
   OUTALU_reg_12_inst : DLH_X1 port map( G => n211_port, D => N202, Q => 
                           OUTALU(12));
   OUTALU_reg_11_inst : DLH_X1 port map( G => n209_port, D => N201, Q => 
                           OUTALU(11));
   OUTALU_reg_10_inst : DLH_X1 port map( G => n210_port, D => N200, Q => 
                           OUTALU(10));
   OUTALU_reg_9_inst : DLH_X1 port map( G => n209_port, D => N199, Q => 
                           OUTALU(9));
   OUTALU_reg_8_inst : DLH_X1 port map( G => n210_port, D => N198, Q => 
                           OUTALU(8));
   OUTALU_reg_7_inst : DLH_X1 port map( G => n210_port, D => N197, Q => 
                           OUTALU(7));
   OUTALU_reg_6_inst : DLH_X1 port map( G => n210_port, D => N196, Q => 
                           OUTALU(6));
   OUTALU_reg_5_inst : DLH_X1 port map( G => n209_port, D => N195, Q => 
                           OUTALU(5));
   OUTALU_reg_4_inst : DLH_X1 port map( G => n210_port, D => N194, Q => 
                           OUTALU(4));
   OUTALU_reg_3_inst : DLH_X1 port map( G => n211_port, D => N193, Q => 
                           OUTALU(3));
   OUTALU_reg_2_inst : DLH_X1 port map( G => n211_port, D => N192, Q => 
                           OUTALU(2));
   OUTALU_reg_1_inst : DLH_X1 port map( G => n209_port, D => N191, Q => 
                           OUTALU(1));
   OUTALU_reg_0_inst : DLH_X1 port map( G => n211_port, D => N190, Q => 
                           OUTALU(0));
   n3 <= '0';
   n4 <= '0';
   srl_39 : logic_and_shift_N32_DW_rash_0 port map( A(31) => DATA1(31), A(30) 
                           => DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28)
                           , A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), DATA_TC => n3,
                           SH(30) => DATA2(30), SH(29) => DATA2(29), SH(28) => 
                           DATA2(28), SH(27) => DATA2(27), SH(26) => DATA2(26),
                           SH(25) => DATA2(25), SH(24) => DATA2(24), SH(23) => 
                           DATA2(23), SH(22) => DATA2(22), SH(21) => DATA2(21),
                           SH(20) => DATA2(20), SH(19) => DATA2(19), SH(18) => 
                           DATA2(18), SH(17) => DATA2(17), SH(16) => DATA2(16),
                           SH(15) => DATA2(15), SH(14) => DATA2(14), SH(13) => 
                           DATA2(13), SH(12) => DATA2(12), SH(11) => DATA2(11),
                           SH(10) => DATA2(10), SH(9) => DATA2(9), SH(8) => 
                           DATA2(8), SH(7) => DATA2(7), SH(6) => DATA2(6), 
                           SH(5) => DATA2(5), SH(4) => DATA2(4), SH(3) => 
                           DATA2(3), SH(2) => DATA2(2), SH(1) => DATA2(1), 
                           SH(0) => DATA2(0), SH_TC => n3, B(31) => N92, B(30) 
                           => N91, B(29) => N90, B(28) => N89, B(27) => N88, 
                           B(26) => N87, B(25) => N86, B(24) => N85, B(23) => 
                           N84, B(22) => N83, B(21) => N82, B(20) => N81, B(19)
                           => N80, B(18) => N79, B(17) => N78, B(16) => N77, 
                           B(15) => N76, B(14) => N75, B(13) => N74, B(12) => 
                           N73, B(11) => N72, B(10) => N71, B(9) => N70, B(8) 
                           => N69, B(7) => N68, B(6) => N67, B(5) => N66, B(4) 
                           => N65, B(3) => N64, B(2) => N63, B(1) => N62, B(0) 
                           => N61);
   sll_37 : logic_and_shift_N32_DW01_ash_0 port map( A(31) => DATA1(31), A(30) 
                           => DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28)
                           , A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), DATA_TC => n4,
                           SH(30) => DATA2(30), SH(29) => DATA2(29), SH(28) => 
                           DATA2(28), SH(27) => DATA2(27), SH(26) => DATA2(26),
                           SH(25) => DATA2(25), SH(24) => DATA2(24), SH(23) => 
                           DATA2(23), SH(22) => DATA2(22), SH(21) => DATA2(21),
                           SH(20) => DATA2(20), SH(19) => DATA2(19), SH(18) => 
                           DATA2(18), SH(17) => DATA2(17), SH(16) => DATA2(16),
                           SH(15) => DATA2(15), SH(14) => DATA2(14), SH(13) => 
                           DATA2(13), SH(12) => DATA2(12), SH(11) => DATA2(11),
                           SH(10) => DATA2(10), SH(9) => DATA2(9), SH(8) => 
                           DATA2(8), SH(7) => DATA2(7), SH(6) => DATA2(6), 
                           SH(5) => DATA2(5), SH(4) => DATA2(4), SH(3) => 
                           DATA2(3), SH(2) => DATA2(2), SH(1) => DATA2(1), 
                           SH(0) => DATA2(0), SH_TC => n4, B(31) => N60, B(30) 
                           => N59, B(29) => N58, B(28) => N57, B(27) => N56, 
                           B(26) => N55, B(25) => N54, B(24) => N53, B(23) => 
                           N52, B(22) => N51, B(21) => N50, B(20) => N49, B(19)
                           => N48, B(18) => N47, B(17) => N46, B(16) => N45, 
                           B(15) => N44, B(14) => N43, B(13) => N42, B(12) => 
                           N41, B(11) => N40, B(10) => N39, B(9) => N38, B(8) 
                           => N37, B(7) => N36, B(6) => N35, B(5) => N34, B(4) 
                           => N33, B(3) => N32, B(2) => N31, B(1) => N30, B(0) 
                           => N29);
   U5 : BUF_X1 port map( A => n207_port, Z => n220_port);
   U6 : BUF_X1 port map( A => n208_port, Z => n239);
   U7 : BUF_X1 port map( A => n208_port, Z => n238);
   U8 : BUF_X1 port map( A => n207_port, Z => n219_port);
   U9 : AND2_X1 port map( A1 => n231, A2 => FUNC(3), ZN => n207_port);
   U10 : NOR3_X1 port map( A1 => n305, A2 => FUNC(3), A3 => n304, ZN => 
                           n208_port);
   U11 : BUF_X1 port map( A => n74_port, Z => n228);
   U12 : BUF_X1 port map( A => n73_port, Z => n232);
   U13 : BUF_X1 port map( A => n173, Z => n212_port);
   U14 : BUF_X1 port map( A => n75_port, Z => n221_port);
   U15 : OAI221_X1 port map( B1 => n170, B2 => n240, C1 => n171, C2 => n272, A 
                           => n172, ZN => N190);
   U16 : AOI21_X1 port map( B1 => n235, B2 => n272, A => n218_port, ZN => n170)
                           ;
   U17 : AOI22_X1 port map( A1 => N61, A2 => n224, B1 => N29, B2 => n227, ZN =>
                           n172);
   U18 : AOI221_X1 port map( B1 => n233, B2 => n240, C1 => DATA1(0), C2 => n231
                           , A => n215_port, ZN => n171);
   U19 : OAI221_X1 port map( B1 => n167, B2 => n241, C1 => n168, C2 => n273, A 
                           => n169, ZN => N191);
   U20 : AOI21_X1 port map( B1 => n238, B2 => n273, A => n217_port, ZN => n167)
                           ;
   U21 : AOI22_X1 port map( A1 => N62, A2 => n224, B1 => N30, B2 => n227, ZN =>
                           n169);
   U22 : AOI221_X1 port map( B1 => n233, B2 => n241, C1 => DATA1(1), C2 => n231
                           , A => n215_port, ZN => n168);
   U23 : OAI221_X1 port map( B1 => n164, B2 => n242, C1 => n165, C2 => n274, A 
                           => n166, ZN => N192);
   U24 : AOI21_X1 port map( B1 => n237, B2 => n274, A => n217_port, ZN => n164)
                           ;
   U25 : AOI22_X1 port map( A1 => N63, A2 => n224, B1 => N31, B2 => n227, ZN =>
                           n166);
   U26 : AOI221_X1 port map( B1 => n233, B2 => n242, C1 => DATA1(2), C2 => n231
                           , A => n215_port, ZN => n165);
   U27 : OAI221_X1 port map( B1 => n161, B2 => n243, C1 => n162, C2 => n275, A 
                           => n163, ZN => N193);
   U28 : AOI21_X1 port map( B1 => n237, B2 => n275, A => n217_port, ZN => n161)
                           ;
   U29 : AOI22_X1 port map( A1 => N64, A2 => n224, B1 => N32, B2 => n227, ZN =>
                           n163);
   U30 : AOI221_X1 port map( B1 => n233, B2 => n243, C1 => DATA1(3), C2 => n231
                           , A => n215_port, ZN => n162);
   U31 : OAI221_X1 port map( B1 => n158, B2 => n244, C1 => n159, C2 => n276, A 
                           => n160, ZN => N194);
   U32 : AOI21_X1 port map( B1 => n237, B2 => n276, A => n217_port, ZN => n158)
                           ;
   U33 : AOI22_X1 port map( A1 => N65, A2 => n224, B1 => N33, B2 => n227, ZN =>
                           n160);
   U34 : AOI221_X1 port map( B1 => n233, B2 => n244, C1 => DATA1(4), C2 => n231
                           , A => n215_port, ZN => n159);
   U35 : OAI221_X1 port map( B1 => n155, B2 => n245, C1 => n156, C2 => n277, A 
                           => n157, ZN => N195);
   U36 : AOI21_X1 port map( B1 => n237, B2 => n277, A => n216_port, ZN => n155)
                           ;
   U37 : AOI22_X1 port map( A1 => N66, A2 => n224, B1 => N34, B2 => n227, ZN =>
                           n157);
   U38 : AOI221_X1 port map( B1 => n233, B2 => n245, C1 => DATA1(5), C2 => n231
                           , A => n215_port, ZN => n156);
   U39 : OAI221_X1 port map( B1 => n152, B2 => n246, C1 => n153, C2 => n278, A 
                           => n154, ZN => N196);
   U40 : AOI21_X1 port map( B1 => n237, B2 => n278, A => n216_port, ZN => n152)
                           ;
   U41 : AOI22_X1 port map( A1 => N67, A2 => n224, B1 => N35, B2 => n227, ZN =>
                           n154);
   U42 : AOI221_X1 port map( B1 => n234, B2 => n246, C1 => DATA1(6), C2 => n231
                           , A => n215_port, ZN => n153);
   U43 : OAI221_X1 port map( B1 => n149, B2 => n247, C1 => n150, C2 => n279, A 
                           => n151, ZN => N197);
   U44 : AOI21_X1 port map( B1 => n237, B2 => n279, A => n216_port, ZN => n149)
                           ;
   U45 : AOI22_X1 port map( A1 => N68, A2 => n224, B1 => N36, B2 => n227, ZN =>
                           n151);
   U46 : AOI221_X1 port map( B1 => n233, B2 => n247, C1 => DATA1(7), C2 => n231
                           , A => n214_port, ZN => n150);
   U47 : OAI221_X1 port map( B1 => n146, B2 => n248, C1 => n147, C2 => n280, A 
                           => n148, ZN => N198);
   U48 : AOI21_X1 port map( B1 => n237, B2 => n280, A => n216_port, ZN => n146)
                           ;
   U49 : AOI22_X1 port map( A1 => N69, A2 => n224, B1 => N37, B2 => n227, ZN =>
                           n148);
   U50 : AOI221_X1 port map( B1 => n234, B2 => n248, C1 => DATA1(8), C2 => n230
                           , A => n215_port, ZN => n147);
   U51 : OAI221_X1 port map( B1 => n143, B2 => n249, C1 => n144, C2 => n281, A 
                           => n145, ZN => N199);
   U52 : AOI21_X1 port map( B1 => n237, B2 => n281, A => n216_port, ZN => n143)
                           ;
   U53 : AOI22_X1 port map( A1 => N70, A2 => n223, B1 => N38, B2 => n226, ZN =>
                           n145);
   U54 : AOI221_X1 port map( B1 => n234, B2 => n249, C1 => DATA1(9), C2 => n230
                           , A => n214_port, ZN => n144);
   U55 : OAI221_X1 port map( B1 => n140, B2 => n250, C1 => n141, C2 => n282, A 
                           => n142, ZN => N200);
   U56 : AOI21_X1 port map( B1 => n237, B2 => n282, A => n215_port, ZN => n140)
                           ;
   U57 : AOI22_X1 port map( A1 => N71, A2 => n223, B1 => N39, B2 => n226, ZN =>
                           n142);
   U58 : AOI221_X1 port map( B1 => n234, B2 => n250, C1 => DATA1(10), C2 => 
                           n230, A => n214_port, ZN => n141);
   U59 : OAI221_X1 port map( B1 => n137, B2 => n251, C1 => n138, C2 => n283, A 
                           => n139, ZN => N201);
   U60 : AOI21_X1 port map( B1 => n237, B2 => n283, A => n215_port, ZN => n137)
                           ;
   U61 : AOI22_X1 port map( A1 => N72, A2 => n223, B1 => N40, B2 => n226, ZN =>
                           n139);
   U62 : AOI221_X1 port map( B1 => n233, B2 => n251, C1 => DATA1(11), C2 => 
                           n230, A => n214_port, ZN => n138);
   U63 : OAI221_X1 port map( B1 => n134, B2 => n252, C1 => n135, C2 => n284, A 
                           => n136, ZN => N202);
   U64 : AOI21_X1 port map( B1 => n237, B2 => n284, A => n216_port, ZN => n134)
                           ;
   U65 : AOI22_X1 port map( A1 => N73, A2 => n223, B1 => N41, B2 => n226, ZN =>
                           n136);
   U66 : AOI221_X1 port map( B1 => n234, B2 => n252, C1 => DATA1(12), C2 => 
                           n230, A => n214_port, ZN => n135);
   U67 : OAI221_X1 port map( B1 => n131, B2 => n253, C1 => n132, C2 => n285, A 
                           => n133, ZN => N203);
   U68 : AOI21_X1 port map( B1 => n237, B2 => n285, A => n215_port, ZN => n131)
                           ;
   U69 : AOI22_X1 port map( A1 => N74, A2 => n223, B1 => N42, B2 => n226, ZN =>
                           n133);
   U70 : AOI221_X1 port map( B1 => n234, B2 => n253, C1 => DATA1(13), C2 => 
                           n230, A => n214_port, ZN => n132);
   U71 : OAI221_X1 port map( B1 => n128, B2 => n254, C1 => n129, C2 => n286, A 
                           => n130, ZN => N204);
   U72 : AOI21_X1 port map( B1 => n237, B2 => n286, A => n215_port, ZN => n128)
                           ;
   U73 : AOI22_X1 port map( A1 => N75, A2 => n223, B1 => N43, B2 => n226, ZN =>
                           n130);
   U74 : AOI221_X1 port map( B1 => n235, B2 => n254, C1 => DATA1(14), C2 => 
                           n230, A => n214_port, ZN => n129);
   U75 : OAI221_X1 port map( B1 => n125, B2 => n255, C1 => n126, C2 => n287, A 
                           => n127, ZN => N205);
   U76 : AOI21_X1 port map( B1 => n236, B2 => n287, A => n216_port, ZN => n125)
                           ;
   U77 : AOI22_X1 port map( A1 => N76, A2 => n223, B1 => N44, B2 => n226, ZN =>
                           n127);
   U78 : AOI221_X1 port map( B1 => n235, B2 => n255, C1 => DATA1(15), C2 => 
                           n230, A => n214_port, ZN => n126);
   U79 : OAI221_X1 port map( B1 => n122, B2 => n256, C1 => n123, C2 => n288, A 
                           => n124, ZN => N206);
   U80 : AOI21_X1 port map( B1 => n236, B2 => n288, A => n216_port, ZN => n122)
                           ;
   U81 : AOI22_X1 port map( A1 => N77, A2 => n223, B1 => N45, B2 => n226, ZN =>
                           n124);
   U82 : AOI221_X1 port map( B1 => n234, B2 => n256, C1 => DATA1(16), C2 => 
                           n230, A => n214_port, ZN => n123);
   U83 : OAI221_X1 port map( B1 => n119, B2 => n257, C1 => n120, C2 => n289, A 
                           => n121, ZN => N207);
   U84 : AOI21_X1 port map( B1 => n236, B2 => n289, A => n216_port, ZN => n119)
                           ;
   U85 : AOI22_X1 port map( A1 => N78, A2 => n223, B1 => N46, B2 => n226, ZN =>
                           n121);
   U86 : AOI221_X1 port map( B1 => n235, B2 => n257, C1 => DATA1(17), C2 => 
                           n230, A => n214_port, ZN => n120);
   U87 : OAI221_X1 port map( B1 => n116, B2 => n258, C1 => n117, C2 => n290, A 
                           => n118, ZN => N208);
   U88 : AOI21_X1 port map( B1 => n236, B2 => n290, A => n216_port, ZN => n116)
                           ;
   U89 : AOI22_X1 port map( A1 => N79, A2 => n223, B1 => N47, B2 => n226, ZN =>
                           n118);
   U90 : AOI221_X1 port map( B1 => n235, B2 => n258, C1 => DATA1(18), C2 => 
                           n230, A => n214_port, ZN => n117);
   U91 : OAI221_X1 port map( B1 => n113, B2 => n259, C1 => n114, C2 => n291, A 
                           => n115, ZN => N209);
   U92 : AOI21_X1 port map( B1 => n236, B2 => n291, A => n216_port, ZN => n113)
                           ;
   U93 : AOI22_X1 port map( A1 => N80, A2 => n223, B1 => N48, B2 => n226, ZN =>
                           n115);
   U94 : AOI221_X1 port map( B1 => n235, B2 => n259, C1 => DATA1(19), C2 => 
                           n229, A => n213_port, ZN => n114);
   U95 : OAI221_X1 port map( B1 => n110, B2 => n260, C1 => n111, C2 => n292, A 
                           => n112, ZN => N210);
   U96 : AOI21_X1 port map( B1 => n236, B2 => n292, A => n216_port, ZN => n110)
                           ;
   U97 : AOI22_X1 port map( A1 => N81, A2 => n223, B1 => N49, B2 => n226, ZN =>
                           n112);
   U98 : AOI221_X1 port map( B1 => n235, B2 => n260, C1 => DATA1(20), C2 => 
                           n229, A => n213_port, ZN => n111);
   U99 : OAI221_X1 port map( B1 => n107, B2 => n261, C1 => n108, C2 => n293, A 
                           => n109, ZN => N211);
   U100 : AOI21_X1 port map( B1 => n236, B2 => n293, A => n217_port, ZN => n107
                           );
   U101 : AOI22_X1 port map( A1 => N82, A2 => n222, B1 => N50, B2 => n225, ZN 
                           => n109);
   U102 : AOI221_X1 port map( B1 => n234, B2 => n261, C1 => DATA1(21), C2 => 
                           n229, A => n213_port, ZN => n108);
   U103 : OAI221_X1 port map( B1 => n104, B2 => n262, C1 => n105, C2 => n294, A
                           => n106, ZN => N212);
   U104 : AOI21_X1 port map( B1 => n236, B2 => n294, A => n216_port, ZN => n104
                           );
   U105 : AOI22_X1 port map( A1 => N83, A2 => n222, B1 => N51, B2 => n225, ZN 
                           => n106);
   U106 : AOI221_X1 port map( B1 => n235, B2 => n262, C1 => DATA1(22), C2 => 
                           n229, A => n213_port, ZN => n105);
   U107 : OAI221_X1 port map( B1 => n101, B2 => n263, C1 => n102, C2 => n295, A
                           => n103, ZN => N213);
   U108 : AOI21_X1 port map( B1 => n236, B2 => n295, A => n217_port, ZN => n101
                           );
   U109 : AOI22_X1 port map( A1 => N84, A2 => n222, B1 => N52, B2 => n225, ZN 
                           => n103);
   U110 : AOI221_X1 port map( B1 => n235, B2 => n263, C1 => DATA1(23), C2 => 
                           n229, A => n213_port, ZN => n102);
   U111 : OAI221_X1 port map( B1 => n98, B2 => n264, C1 => n99, C2 => n296, A 
                           => n100, ZN => N214);
   U112 : AOI21_X1 port map( B1 => n236, B2 => n296, A => n217_port, ZN => n98)
                           ;
   U113 : AOI22_X1 port map( A1 => N85, A2 => n222, B1 => N53, B2 => n225, ZN 
                           => n100);
   U114 : AOI221_X1 port map( B1 => n234, B2 => n264, C1 => DATA1(24), C2 => 
                           n230, A => n213_port, ZN => n99);
   U115 : OAI221_X1 port map( B1 => n95, B2 => n265, C1 => n96, C2 => n297, A 
                           => n97, ZN => N215);
   U116 : AOI21_X1 port map( B1 => n235, B2 => n297, A => n217_port, ZN => n95)
                           ;
   U117 : AOI22_X1 port map( A1 => N86, A2 => n222, B1 => N54, B2 => n225, ZN 
                           => n97);
   U118 : AOI221_X1 port map( B1 => n234, B2 => n265, C1 => DATA1(25), C2 => 
                           n229, A => n213_port, ZN => n96);
   U119 : OAI221_X1 port map( B1 => n92_port, B2 => n266, C1 => n93, C2 => n298
                           , A => n94, ZN => N216);
   U120 : AOI21_X1 port map( B1 => n236, B2 => n298, A => n217_port, ZN => 
                           n92_port);
   U121 : AOI22_X1 port map( A1 => N87, A2 => n222, B1 => N55, B2 => n225, ZN 
                           => n94);
   U122 : AOI221_X1 port map( B1 => n234, B2 => n266, C1 => DATA1(26), C2 => 
                           n229, A => n213_port, ZN => n93);
   U123 : OAI221_X1 port map( B1 => n89_port, B2 => n267, C1 => n90_port, C2 =>
                           n299, A => n91_port, ZN => N217);
   U124 : AOI21_X1 port map( B1 => n235, B2 => n299, A => n217_port, ZN => 
                           n89_port);
   U125 : AOI22_X1 port map( A1 => N88, A2 => n222, B1 => N56, B2 => n225, ZN 
                           => n91_port);
   U126 : AOI221_X1 port map( B1 => n234, B2 => n267, C1 => DATA1(27), C2 => 
                           n229, A => n213_port, ZN => n90_port);
   U127 : OAI221_X1 port map( B1 => n86_port, B2 => n268, C1 => n87_port, C2 =>
                           n300, A => n88_port, ZN => N218);
   U128 : AOI21_X1 port map( B1 => n235, B2 => n300, A => n217_port, ZN => 
                           n86_port);
   U129 : AOI22_X1 port map( A1 => N89, A2 => n222, B1 => N57, B2 => n225, ZN 
                           => n88_port);
   U130 : AOI221_X1 port map( B1 => n234, B2 => n268, C1 => DATA1(28), C2 => 
                           n229, A => n213_port, ZN => n87_port);
   U131 : OAI221_X1 port map( B1 => n83_port, B2 => n269, C1 => n84_port, C2 =>
                           n301, A => n85_port, ZN => N219);
   U132 : AOI21_X1 port map( B1 => n236, B2 => n301, A => n217_port, ZN => 
                           n83_port);
   U133 : AOI22_X1 port map( A1 => N90, A2 => n222, B1 => N58, B2 => n225, ZN 
                           => n85_port);
   U134 : AOI221_X1 port map( B1 => n233, B2 => n269, C1 => DATA1(29), C2 => 
                           n229, A => n213_port, ZN => n84_port);
   U135 : OAI221_X1 port map( B1 => n80_port, B2 => n270, C1 => n81_port, C2 =>
                           n302, A => n82_port, ZN => N220);
   U136 : AOI21_X1 port map( B1 => n235, B2 => n302, A => n217_port, ZN => 
                           n80_port);
   U137 : AOI22_X1 port map( A1 => N91, A2 => n222, B1 => N59, B2 => n225, ZN 
                           => n82_port);
   U138 : AOI221_X1 port map( B1 => n233, B2 => n270, C1 => DATA1(30), C2 => 
                           n229, A => n213_port, ZN => n81_port);
   U139 : OAI221_X1 port map( B1 => n76_port, B2 => n271, C1 => n77_port, C2 =>
                           n303, A => n78_port, ZN => N221);
   U140 : AOI21_X1 port map( B1 => n236, B2 => n303, A => n218_port, ZN => 
                           n76_port);
   U141 : AOI22_X1 port map( A1 => N92, A2 => n222, B1 => N60, B2 => n225, ZN 
                           => n78_port);
   U142 : AOI221_X1 port map( B1 => n233, B2 => n271, C1 => DATA1(31), C2 => 
                           n229, A => n214_port, ZN => n77_port);
   U143 : INV_X1 port map( A => DATA2(3), ZN => n275);
   U144 : INV_X1 port map( A => DATA2(1), ZN => n273);
   U145 : INV_X1 port map( A => DATA2(4), ZN => n276);
   U146 : INV_X1 port map( A => DATA1(30), ZN => n270);
   U147 : INV_X1 port map( A => DATA1(14), ZN => n254);
   U148 : INV_X1 port map( A => DATA1(29), ZN => n269);
   U149 : INV_X1 port map( A => DATA2(2), ZN => n274);
   U150 : INV_X1 port map( A => DATA1(11), ZN => n251);
   U151 : INV_X1 port map( A => DATA1(26), ZN => n266);
   U152 : INV_X1 port map( A => DATA1(12), ZN => n252);
   U153 : INV_X1 port map( A => DATA1(13), ZN => n253);
   U154 : INV_X1 port map( A => DATA1(27), ZN => n267);
   U155 : INV_X1 port map( A => DATA1(28), ZN => n268);
   U156 : INV_X1 port map( A => DATA1(19), ZN => n259);
   U157 : INV_X1 port map( A => DATA1(18), ZN => n258);
   U158 : INV_X1 port map( A => DATA1(31), ZN => n271);
   U159 : INV_X1 port map( A => DATA2(0), ZN => n272);
   U160 : INV_X1 port map( A => DATA1(7), ZN => n247);
   U161 : INV_X1 port map( A => DATA1(8), ZN => n248);
   U162 : INV_X1 port map( A => DATA1(9), ZN => n249);
   U163 : INV_X1 port map( A => DATA1(10), ZN => n250);
   U164 : INV_X1 port map( A => DATA1(15), ZN => n255);
   U165 : INV_X1 port map( A => DATA1(2), ZN => n242);
   U166 : INV_X1 port map( A => DATA1(20), ZN => n260);
   U167 : INV_X1 port map( A => DATA1(21), ZN => n261);
   U168 : INV_X1 port map( A => DATA1(22), ZN => n262);
   U169 : INV_X1 port map( A => DATA1(17), ZN => n257);
   U170 : INV_X1 port map( A => DATA1(6), ZN => n246);
   U171 : INV_X1 port map( A => DATA1(25), ZN => n265);
   U172 : INV_X1 port map( A => DATA1(3), ZN => n243);
   U173 : INV_X1 port map( A => DATA1(23), ZN => n263);
   U174 : INV_X1 port map( A => DATA1(1), ZN => n241);
   U175 : INV_X1 port map( A => DATA2(30), ZN => n302);
   U176 : INV_X1 port map( A => DATA1(0), ZN => n240);
   U177 : INV_X1 port map( A => DATA2(11), ZN => n283);
   U178 : INV_X1 port map( A => DATA2(17), ZN => n289);
   U179 : INV_X1 port map( A => DATA2(24), ZN => n296);
   U180 : INV_X1 port map( A => DATA2(12), ZN => n284);
   U181 : INV_X1 port map( A => DATA2(18), ZN => n290);
   U182 : INV_X1 port map( A => DATA2(23), ZN => n295);
   U183 : INV_X1 port map( A => DATA2(29), ZN => n301);
   U184 : INV_X1 port map( A => DATA1(4), ZN => n244);
   U185 : INV_X1 port map( A => DATA1(5), ZN => n245);
   U186 : INV_X1 port map( A => DATA1(16), ZN => n256);
   U187 : INV_X1 port map( A => DATA1(24), ZN => n264);
   U188 : INV_X1 port map( A => DATA2(10), ZN => n282);
   U189 : INV_X1 port map( A => DATA2(16), ZN => n288);
   U190 : INV_X1 port map( A => DATA2(28), ZN => n300);
   U191 : INV_X1 port map( A => DATA2(6), ZN => n278);
   U192 : INV_X1 port map( A => DATA2(22), ZN => n294);
   U193 : INV_X1 port map( A => DATA2(5), ZN => n277);
   U194 : INV_X1 port map( A => DATA2(13), ZN => n285);
   U195 : INV_X1 port map( A => DATA2(25), ZN => n297);
   U196 : INV_X1 port map( A => DATA2(26), ZN => n298);
   U197 : INV_X1 port map( A => DATA2(14), ZN => n286);
   U198 : INV_X1 port map( A => DATA2(27), ZN => n299);
   U199 : INV_X1 port map( A => DATA2(15), ZN => n287);
   U200 : INV_X1 port map( A => DATA2(8), ZN => n280);
   U201 : INV_X1 port map( A => DATA2(21), ZN => n293);
   U202 : INV_X1 port map( A => DATA2(7), ZN => n279);
   U203 : INV_X1 port map( A => DATA2(9), ZN => n281);
   U204 : INV_X1 port map( A => DATA2(19), ZN => n291);
   U205 : INV_X1 port map( A => DATA2(20), ZN => n292);
   U206 : BUF_X1 port map( A => n239, Z => n234);
   U207 : BUF_X1 port map( A => n239, Z => n235);
   U208 : BUF_X1 port map( A => n220_port, Z => n213_port);
   U209 : BUF_X1 port map( A => n220_port, Z => n214_port);
   U210 : BUF_X1 port map( A => n219_port, Z => n216_port);
   U211 : BUF_X1 port map( A => n219_port, Z => n217_port);
   U212 : BUF_X1 port map( A => n238, Z => n237);
   U213 : BUF_X1 port map( A => n238, Z => n236);
   U214 : BUF_X1 port map( A => n220_port, Z => n215_port);
   U215 : BUF_X1 port map( A => n239, Z => n233);
   U216 : BUF_X1 port map( A => n219_port, Z => n218_port);
   U217 : INV_X1 port map( A => DATA2(31), ZN => n303);
   U218 : BUF_X1 port map( A => n232, Z => n230);
   U219 : BUF_X1 port map( A => n232, Z => n229);
   U220 : BUF_X1 port map( A => n221_port, Z => n222);
   U221 : BUF_X1 port map( A => n228, Z => n225);
   U222 : BUF_X1 port map( A => n228, Z => n226);
   U223 : BUF_X1 port map( A => n221_port, Z => n223);
   U224 : BUF_X1 port map( A => n232, Z => n231);
   U225 : BUF_X1 port map( A => n228, Z => n227);
   U226 : BUF_X1 port map( A => n221_port, Z => n224);
   U227 : BUF_X1 port map( A => n212_port, Z => n210_port);
   U228 : BUF_X1 port map( A => n212_port, Z => n209_port);
   U229 : BUF_X1 port map( A => n212_port, Z => n211_port);
   U230 : INV_X1 port map( A => FUNC(2), ZN => n305);
   U231 : INV_X1 port map( A => FUNC(1), ZN => n304);
   U232 : NOR3_X1 port map( A1 => FUNC(2), A2 => FUNC(1), A3 => FUNC(3), ZN => 
                           n74_port);
   U233 : NOR2_X1 port map( A1 => n304, A2 => FUNC(2), ZN => n73_port);
   U234 : NOR2_X1 port map( A1 => FUNC(0), A2 => n71_port, ZN => n173);
   U235 : NOR4_X1 port map( A1 => n233, A2 => n231, A3 => n225, A4 => n222, ZN 
                           => n71_port);
   U236 : AND3_X1 port map( A1 => n305, A2 => n304, A3 => FUNC(3), ZN => 
                           n75_port);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity P4_ADDER_NBITS32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end P4_ADDER_NBITS32;

architecture SYN_STRUCTURAL of P4_ADDER_NBITS32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4
      port( A, B : in std_logic_vector (32 downto 1);  C0 : in std_logic;  COUT
            : out std_logic_vector (8 downto 0));
   end component;
   
   component SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (8 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component xor_logic_nbits32
      port( Cin : in std_logic;  B0 : in std_logic_vector (31 downto 0);  B : 
            out std_logic_vector (31 downto 0));
   end component;
   
   signal Co_port, B_diff_31_port, B_diff_30_port, B_diff_29_port, 
      B_diff_28_port, B_diff_27_port, B_diff_26_port, B_diff_25_port, 
      B_diff_24_port, B_diff_23_port, B_diff_22_port, B_diff_21_port, 
      B_diff_20_port, B_diff_19_port, B_diff_18_port, B_diff_17_port, 
      B_diff_16_port, B_diff_15_port, B_diff_14_port, B_diff_13_port, 
      B_diff_12_port, B_diff_11_port, B_diff_10_port, B_diff_9_port, 
      B_diff_8_port, B_diff_7_port, B_diff_6_port, B_diff_5_port, B_diff_4_port
      , B_diff_3_port, B_diff_2_port, B_diff_1_port, B_diff_0_port, 
      fromCarry_to_adder_7_port, fromCarry_to_adder_6_port, 
      fromCarry_to_adder_5_port, fromCarry_to_adder_4_port, 
      fromCarry_to_adder_3_port, fromCarry_to_adder_2_port, 
      fromCarry_to_adder_1_port, fromCarry_to_adder_0_port, n1 : std_logic;

begin
   Co <= Co_port;
   
   xor_gate : xor_logic_nbits32 port map( Cin => Ci, B0(31) => B(31), B0(30) =>
                           B(30), B0(29) => B(29), B0(28) => B(28), B0(27) => 
                           B(27), B0(26) => B(26), B0(25) => B(25), B0(24) => 
                           B(24), B0(23) => B(23), B0(22) => B(22), B0(21) => 
                           B(21), B0(20) => B(20), B0(19) => B(19), B0(18) => 
                           B(18), B0(17) => B(17), B0(16) => B(16), B0(15) => 
                           B(15), B0(14) => B(14), B0(13) => B(13), B0(12) => 
                           B(12), B0(11) => B(11), B0(10) => B(10), B0(9) => 
                           B(9), B0(8) => B(8), B0(7) => B(7), B0(6) => B(6), 
                           B0(5) => B(5), B0(4) => B(4), B0(3) => B(3), B0(2) 
                           => B(2), B0(1) => B(1), B0(0) => B(0), B(31) => 
                           B_diff_31_port, B(30) => B_diff_30_port, B(29) => 
                           B_diff_29_port, B(28) => B_diff_28_port, B(27) => 
                           B_diff_27_port, B(26) => B_diff_26_port, B(25) => 
                           B_diff_25_port, B(24) => B_diff_24_port, B(23) => 
                           B_diff_23_port, B(22) => B_diff_22_port, B(21) => 
                           B_diff_21_port, B(20) => B_diff_20_port, B(19) => 
                           B_diff_19_port, B(18) => B_diff_18_port, B(17) => 
                           B_diff_17_port, B(16) => B_diff_16_port, B(15) => 
                           B_diff_15_port, B(14) => B_diff_14_port, B(13) => 
                           B_diff_13_port, B(12) => B_diff_12_port, B(11) => 
                           B_diff_11_port, B(10) => B_diff_10_port, B(9) => 
                           B_diff_9_port, B(8) => B_diff_8_port, B(7) => 
                           B_diff_7_port, B(6) => B_diff_6_port, B(5) => 
                           B_diff_5_port, B(4) => B_diff_4_port, B(3) => 
                           B_diff_3_port, B(2) => B_diff_2_port, B(1) => 
                           B_diff_1_port, B(0) => B_diff_0_port);
   SUM_GEN : SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8 port map( A(31)
                           => A(31), A(30) => A(30), A(29) => A(29), A(28) => 
                           A(28), A(27) => A(27), A(26) => A(26), A(25) => 
                           A(25), A(24) => A(24), A(23) => A(23), A(22) => 
                           A(22), A(21) => A(21), A(20) => A(20), A(19) => 
                           A(19), A(18) => A(18), A(17) => A(17), A(16) => 
                           A(16), A(15) => A(15), A(14) => A(14), A(13) => 
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => B_diff_31_port, B(30) => B_diff_30_port, 
                           B(29) => B_diff_29_port, B(28) => B_diff_28_port, 
                           B(27) => B_diff_27_port, B(26) => B_diff_26_port, 
                           B(25) => B_diff_25_port, B(24) => B_diff_24_port, 
                           B(23) => B_diff_23_port, B(22) => B_diff_22_port, 
                           B(21) => B_diff_21_port, B(20) => B_diff_20_port, 
                           B(19) => B_diff_19_port, B(18) => B_diff_18_port, 
                           B(17) => B_diff_17_port, B(16) => B_diff_16_port, 
                           B(15) => B_diff_15_port, B(14) => B_diff_14_port, 
                           B(13) => B_diff_13_port, B(12) => B_diff_12_port, 
                           B(11) => B_diff_11_port, B(10) => B_diff_10_port, 
                           B(9) => B_diff_9_port, B(8) => B_diff_8_port, B(7) 
                           => B_diff_7_port, B(6) => B_diff_6_port, B(5) => 
                           B_diff_5_port, B(4) => B_diff_4_port, B(3) => 
                           B_diff_3_port, B(2) => B_diff_2_port, B(1) => 
                           B_diff_1_port, B(0) => n1, Ci(8) => Co_port, Ci(7) 
                           => fromCarry_to_adder_7_port, Ci(6) => 
                           fromCarry_to_adder_6_port, Ci(5) => 
                           fromCarry_to_adder_5_port, Ci(4) => 
                           fromCarry_to_adder_4_port, Ci(3) => 
                           fromCarry_to_adder_3_port, Ci(2) => 
                           fromCarry_to_adder_2_port, Ci(1) => 
                           fromCarry_to_adder_1_port, Ci(0) => 
                           fromCarry_to_adder_0_port, S(31) => S(31), S(30) => 
                           S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));
   CLA : CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4 port map( A(32) => A(31), A(31)
                           => A(30), A(30) => A(29), A(29) => A(28), A(28) => 
                           A(27), A(27) => A(26), A(26) => A(25), A(25) => 
                           A(24), A(24) => A(23), A(23) => A(22), A(22) => 
                           A(21), A(21) => A(20), A(20) => A(19), A(19) => 
                           A(18), A(18) => A(17), A(17) => A(16), A(16) => 
                           A(15), A(15) => A(14), A(14) => A(13), A(13) => 
                           A(12), A(12) => A(11), A(11) => A(10), A(10) => A(9)
                           , A(9) => A(8), A(8) => A(7), A(7) => A(6), A(6) => 
                           A(5), A(5) => A(4), A(4) => A(3), A(3) => A(2), A(2)
                           => A(1), A(1) => A(0), B(32) => B_diff_31_port, 
                           B(31) => B_diff_30_port, B(30) => B_diff_29_port, 
                           B(29) => B_diff_28_port, B(28) => B_diff_27_port, 
                           B(27) => B_diff_26_port, B(26) => B_diff_25_port, 
                           B(25) => B_diff_24_port, B(24) => B_diff_23_port, 
                           B(23) => B_diff_22_port, B(22) => B_diff_21_port, 
                           B(21) => B_diff_20_port, B(20) => B_diff_19_port, 
                           B(19) => B_diff_18_port, B(18) => B_diff_17_port, 
                           B(17) => B_diff_16_port, B(16) => B_diff_15_port, 
                           B(15) => B_diff_14_port, B(14) => B_diff_13_port, 
                           B(13) => B_diff_12_port, B(12) => B_diff_11_port, 
                           B(11) => B_diff_10_port, B(10) => B_diff_9_port, 
                           B(9) => B_diff_8_port, B(8) => B_diff_7_port, B(7) 
                           => B_diff_6_port, B(6) => B_diff_5_port, B(5) => 
                           B_diff_4_port, B(4) => B_diff_3_port, B(3) => 
                           B_diff_2_port, B(2) => B_diff_1_port, B(1) => n1, C0
                           => Ci, COUT(8) => Co_port, COUT(7) => 
                           fromCarry_to_adder_7_port, COUT(6) => 
                           fromCarry_to_adder_6_port, COUT(5) => 
                           fromCarry_to_adder_5_port, COUT(4) => 
                           fromCarry_to_adder_4_port, COUT(3) => 
                           fromCarry_to_adder_3_port, COUT(2) => 
                           fromCarry_to_adder_2_port, COUT(1) => 
                           fromCarry_to_adder_1_port, COUT(0) => 
                           fromCarry_to_adder_0_port);
   U1 : BUF_X1 port map( A => B_diff_0_port, Z => n1);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ctrl_alu_NBITS32 is

   port( A, B : in std_logic_vector (31 downto 0);  FUNC : in std_logic_vector 
         (0 to 3);  Ap4, Bp4 : out std_logic_vector (31 downto 0);  Cin : out 
         std_logic;  Als, Bls : out std_logic_vector (31 downto 0);  enableComp
         : out std_logic);

end ctrl_alu_NBITS32;

architecture SYN_BEHAVIORAL of ctrl_alu_NBITS32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n70, n71, n72, n73, n74, n75, n77, n78, n79, n80, n81, n82, n83, n84,
      n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99
      , n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n161, n162, n163 : std_logic;

begin
   
   U206 : NAND3_X1 port map( A1 => n161, A2 => n159, A3 => FUNC(2), ZN => n71);
   U3 : NOR2_X1 port map( A1 => n87, A2 => n95, ZN => Ap4(0));
   U4 : NOR2_X1 port map( A1 => n87, A2 => n96, ZN => Ap4(1));
   U5 : NOR2_X1 port map( A1 => n89, A2 => n99, ZN => Ap4(4));
   U6 : NOR2_X1 port map( A1 => n89, A2 => n100, ZN => Ap4(5));
   U7 : NOR2_X1 port map( A1 => n89, A2 => n103, ZN => Ap4(8));
   U8 : NOR2_X1 port map( A1 => n89, A2 => n104, ZN => Ap4(9));
   U9 : NOR2_X1 port map( A1 => n87, A2 => n107, ZN => Ap4(12));
   U10 : NOR2_X1 port map( A1 => n87, A2 => n108, ZN => Ap4(13));
   U11 : NOR2_X1 port map( A1 => n87, A2 => n111, ZN => Ap4(16));
   U12 : NOR2_X1 port map( A1 => n87, A2 => n112, ZN => Ap4(17));
   U13 : NOR2_X1 port map( A1 => n88, A2 => n115, ZN => Ap4(20));
   U14 : NOR2_X1 port map( A1 => n88, A2 => n116, ZN => Ap4(21));
   U15 : NOR2_X1 port map( A1 => n88, A2 => n119, ZN => Ap4(24));
   U16 : NOR2_X1 port map( A1 => n88, A2 => n120, ZN => Ap4(25));
   U17 : NOR2_X1 port map( A1 => n88, A2 => n123, ZN => Ap4(28));
   U18 : NOR2_X1 port map( A1 => n88, A2 => n124, ZN => Ap4(29));
   U19 : NOR2_X1 port map( A1 => n89, A2 => n101, ZN => Ap4(6));
   U20 : NOR2_X1 port map( A1 => n87, A2 => n105, ZN => Ap4(10));
   U21 : NOR2_X1 port map( A1 => n87, A2 => n109, ZN => Ap4(14));
   U22 : NOR2_X1 port map( A1 => n87, A2 => n113, ZN => Ap4(18));
   U23 : NOR2_X1 port map( A1 => n88, A2 => n117, ZN => Ap4(22));
   U24 : NOR2_X1 port map( A1 => n88, A2 => n121, ZN => Ap4(26));
   U25 : NOR2_X1 port map( A1 => n88, A2 => n125, ZN => Ap4(30));
   U26 : NOR2_X1 port map( A1 => n88, A2 => n97, ZN => Ap4(2));
   U27 : NOR2_X1 port map( A1 => n128, A2 => n79, ZN => Bls(1));
   U28 : NOR2_X1 port map( A1 => n131, A2 => n78, ZN => Bls(4));
   U29 : NOR2_X1 port map( A1 => n130, A2 => n78, ZN => Bls(3));
   U30 : NOR2_X1 port map( A1 => n89, A2 => n102, ZN => Ap4(7));
   U31 : NOR2_X1 port map( A1 => n87, A2 => n106, ZN => Ap4(11));
   U32 : NOR2_X1 port map( A1 => n87, A2 => n110, ZN => Ap4(15));
   U33 : NOR2_X1 port map( A1 => n87, A2 => n114, ZN => Ap4(19));
   U34 : NOR2_X1 port map( A1 => n88, A2 => n118, ZN => Ap4(23));
   U35 : NOR2_X1 port map( A1 => n88, A2 => n122, ZN => Ap4(27));
   U36 : NOR2_X1 port map( A1 => n89, A2 => n98, ZN => Ap4(3));
   U37 : BUF_X1 port map( A => n86, Z => n94);
   U38 : BUF_X1 port map( A => n86, Z => n93);
   U39 : BUF_X1 port map( A => n72, Z => n86);
   U40 : BUF_X1 port map( A => n77, Z => n85);
   U41 : BUF_X1 port map( A => n77, Z => n84);
   U42 : BUF_X1 port map( A => n94, Z => n89);
   U43 : BUF_X1 port map( A => n93, Z => n91);
   U44 : BUF_X1 port map( A => n93, Z => n90);
   U45 : BUF_X1 port map( A => n94, Z => n87);
   U46 : BUF_X1 port map( A => n93, Z => n92);
   U47 : BUF_X1 port map( A => n94, Z => n88);
   U48 : BUF_X1 port map( A => n85, Z => n78);
   U49 : BUF_X1 port map( A => n85, Z => n79);
   U50 : BUF_X1 port map( A => n85, Z => n80);
   U51 : BUF_X1 port map( A => n84, Z => n82);
   U52 : BUF_X1 port map( A => n84, Z => n81);
   U53 : BUF_X1 port map( A => n84, Z => n83);
   U54 : INV_X1 port map( A => n70, ZN => enableComp);
   U55 : NOR2_X1 port map( A1 => n89, A2 => n127, ZN => Bp4(0));
   U56 : OAI21_X1 port map( B1 => n163, B2 => n71, A => n70, ZN => Cin);
   U57 : NOR2_X1 port map( A1 => n91, A2 => n130, ZN => Bp4(3));
   U58 : NOR2_X1 port map( A1 => n90, A2 => n128, ZN => Bp4(1));
   U59 : NOR2_X1 port map( A1 => n91, A2 => n129, ZN => Bp4(2));
   U60 : NOR2_X1 port map( A1 => n91, A2 => n132, ZN => Bp4(5));
   U61 : NOR2_X1 port map( A1 => n92, A2 => n134, ZN => Bp4(7));
   U62 : NOR2_X1 port map( A1 => n91, A2 => n131, ZN => Bp4(4));
   U63 : NOR2_X1 port map( A1 => n92, A2 => n133, ZN => Bp4(6));
   U64 : NOR2_X1 port map( A1 => n92, A2 => n136, ZN => Bp4(9));
   U65 : NOR2_X1 port map( A1 => n89, A2 => n138, ZN => Bp4(11));
   U66 : NOR2_X1 port map( A1 => n90, A2 => n140, ZN => Bp4(13));
   U67 : NOR2_X1 port map( A1 => n91, A2 => n155, ZN => Bp4(28));
   U68 : NOR2_X1 port map( A1 => n90, A2 => n142, ZN => Bp4(15));
   U69 : NOR2_X1 port map( A1 => n92, A2 => n135, ZN => Bp4(8));
   U70 : NOR2_X1 port map( A1 => n90, A2 => n143, ZN => Bp4(16));
   U71 : NOR2_X1 port map( A1 => n89, A2 => n139, ZN => Bp4(12));
   U72 : NOR2_X1 port map( A1 => n89, A2 => n137, ZN => Bp4(10));
   U73 : NOR2_X1 port map( A1 => n90, A2 => n141, ZN => Bp4(14));
   U74 : NOR2_X1 port map( A1 => n90, A2 => n147, ZN => Bp4(20));
   U75 : NOR2_X1 port map( A1 => n90, A2 => n144, ZN => Bp4(17));
   U76 : NOR2_X1 port map( A1 => n90, A2 => n146, ZN => Bp4(19));
   U77 : NOR2_X1 port map( A1 => n91, A2 => n151, ZN => Bp4(24));
   U78 : NOR2_X1 port map( A1 => n90, A2 => n148, ZN => Bp4(21));
   U79 : NOR2_X1 port map( A1 => n90, A2 => n150, ZN => Bp4(23));
   U80 : NOR2_X1 port map( A1 => n90, A2 => n145, ZN => Bp4(18));
   U81 : NOR2_X1 port map( A1 => n90, A2 => n149, ZN => Bp4(22));
   U82 : NOR2_X1 port map( A1 => n91, A2 => n156, ZN => Bp4(29));
   U83 : AND2_X1 port map( A1 => n71, A2 => n70, ZN => n72);
   U84 : NOR2_X1 port map( A1 => n91, A2 => n152, ZN => Bp4(25));
   U85 : NOR2_X1 port map( A1 => n91, A2 => n154, ZN => Bp4(27));
   U86 : NOR2_X1 port map( A1 => n91, A2 => n153, ZN => Bp4(26));
   U87 : NOR2_X1 port map( A1 => n91, A2 => n157, ZN => Bp4(30));
   U88 : NOR2_X1 port map( A1 => n91, A2 => n158, ZN => Bp4(31));
   U89 : NOR2_X1 port map( A1 => n89, A2 => n126, ZN => Ap4(31));
   U90 : NOR2_X1 port map( A1 => n81, A2 => n125, ZN => Als(30));
   U91 : NOR2_X1 port map( A1 => n82, A2 => n109, ZN => Als(14));
   U92 : NOR2_X1 port map( A1 => n81, A2 => n124, ZN => Als(29));
   U93 : NOR2_X1 port map( A1 => n83, A2 => n106, ZN => Als(11));
   U94 : NOR2_X1 port map( A1 => n81, A2 => n121, ZN => Als(26));
   U95 : NOR2_X1 port map( A1 => n83, A2 => n107, ZN => Als(12));
   U96 : NOR2_X1 port map( A1 => n82, A2 => n108, ZN => Als(13));
   U97 : NOR2_X1 port map( A1 => n81, A2 => n122, ZN => Als(27));
   U98 : NOR2_X1 port map( A1 => n81, A2 => n123, ZN => Als(28));
   U99 : NOR2_X1 port map( A1 => n129, A2 => n78, ZN => Bls(2));
   U100 : NOR2_X1 port map( A1 => n82, A2 => n114, ZN => Als(19));
   U101 : NOR2_X1 port map( A1 => n82, A2 => n113, ZN => Als(18));
   U102 : NOR2_X1 port map( A1 => n81, A2 => n126, ZN => Als(31));
   U103 : NOR2_X1 port map( A1 => n127, A2 => n80, ZN => Bls(0));
   U104 : NOR2_X1 port map( A1 => n80, A2 => n102, ZN => Als(7));
   U105 : NOR2_X1 port map( A1 => n80, A2 => n103, ZN => Als(8));
   U106 : NOR2_X1 port map( A1 => n80, A2 => n104, ZN => Als(9));
   U107 : NOR2_X1 port map( A1 => n83, A2 => n105, ZN => Als(10));
   U108 : NOR2_X1 port map( A1 => n82, A2 => n110, ZN => Als(15));
   U109 : NOR2_X1 port map( A1 => n81, A2 => n97, ZN => Als(2));
   U110 : NOR2_X1 port map( A1 => n82, A2 => n115, ZN => Als(20));
   U111 : NOR2_X1 port map( A1 => n82, A2 => n116, ZN => Als(21));
   U112 : NOR2_X1 port map( A1 => n82, A2 => n117, ZN => Als(22));
   U113 : NOR2_X1 port map( A1 => n82, A2 => n112, ZN => Als(17));
   U114 : NOR2_X1 port map( A1 => n80, A2 => n101, ZN => Als(6));
   U115 : NOR2_X1 port map( A1 => n81, A2 => n120, ZN => Als(25));
   U116 : NOR2_X1 port map( A1 => n81, A2 => n98, ZN => Als(3));
   U117 : NOR2_X1 port map( A1 => n82, A2 => n118, ZN => Als(23));
   U118 : NOR2_X1 port map( A1 => n82, A2 => n96, ZN => Als(1));
   U119 : NOR2_X1 port map( A1 => n157, A2 => n78, ZN => Bls(30));
   U120 : NOR2_X1 port map( A1 => n83, A2 => n95, ZN => Als(0));
   U121 : NOR2_X1 port map( A1 => n144, A2 => n79, ZN => Bls(17));
   U122 : NOR2_X1 port map( A1 => n138, A2 => n80, ZN => Bls(11));
   U123 : NOR2_X1 port map( A1 => n151, A2 => n79, ZN => Bls(24));
   U124 : NOR2_X1 port map( A1 => n81, A2 => n99, ZN => Als(4));
   U125 : NOR2_X1 port map( A1 => n81, A2 => n100, ZN => Als(5));
   U126 : NOR2_X1 port map( A1 => n82, A2 => n111, ZN => Als(16));
   U127 : NOR2_X1 port map( A1 => n81, A2 => n119, ZN => Als(24));
   U128 : NOR2_X1 port map( A1 => n145, A2 => n79, ZN => Bls(18));
   U129 : NOR2_X1 port map( A1 => n139, A2 => n80, ZN => Bls(12));
   U130 : NOR2_X1 port map( A1 => n156, A2 => n78, ZN => Bls(29));
   U131 : NOR2_X1 port map( A1 => n150, A2 => n79, ZN => Bls(23));
   U132 : NOR2_X1 port map( A1 => n143, A2 => n80, ZN => Bls(16));
   U133 : NOR2_X1 port map( A1 => n137, A2 => n80, ZN => Bls(10));
   U134 : NOR2_X1 port map( A1 => n155, A2 => n78, ZN => Bls(28));
   U135 : NOR2_X1 port map( A1 => n133, A2 => n78, ZN => Bls(6));
   U136 : NOR2_X1 port map( A1 => n149, A2 => n79, ZN => Bls(22));
   U137 : NOR2_X1 port map( A1 => n152, A2 => n79, ZN => Bls(25));
   U138 : NOR2_X1 port map( A1 => n140, A2 => n80, ZN => Bls(13));
   U139 : NOR2_X1 port map( A1 => n153, A2 => n79, ZN => Bls(26));
   U140 : NOR2_X1 port map( A1 => n141, A2 => n80, ZN => Bls(14));
   U141 : NOR2_X1 port map( A1 => n154, A2 => n79, ZN => Bls(27));
   U142 : NOR2_X1 port map( A1 => n142, A2 => n80, ZN => Bls(15));
   U143 : NOR2_X1 port map( A1 => n132, A2 => n78, ZN => Bls(5));
   U144 : NOR2_X1 port map( A1 => n147, A2 => n79, ZN => Bls(20));
   U145 : NOR2_X1 port map( A1 => n134, A2 => n78, ZN => Bls(7));
   U146 : NOR2_X1 port map( A1 => n146, A2 => n79, ZN => Bls(19));
   U147 : NOR2_X1 port map( A1 => n136, A2 => n78, ZN => Bls(9));
   U148 : NOR2_X1 port map( A1 => n148, A2 => n79, ZN => Bls(21));
   U149 : NOR2_X1 port map( A1 => n135, A2 => n78, ZN => Bls(8));
   U150 : NOR2_X1 port map( A1 => n158, A2 => n78, ZN => Bls(31));
   U151 : INV_X1 port map( A => A(0), ZN => n95);
   U152 : OAI221_X1 port map( B1 => FUNC(0), B2 => FUNC(2), C1 => FUNC(1), C2 
                           => n162, A => n74, ZN => n70);
   U153 : INV_X1 port map( A => FUNC(2), ZN => n162);
   U154 : OAI21_X1 port map( B1 => FUNC(0), B2 => n163, A => FUNC(1), ZN => n74
                           );
   U155 : INV_X1 port map( A => FUNC(3), ZN => n163);
   U156 : INV_X1 port map( A => A(1), ZN => n96);
   U157 : INV_X1 port map( A => A(3), ZN => n98);
   U158 : INV_X1 port map( A => A(5), ZN => n100);
   U159 : INV_X1 port map( A => A(2), ZN => n97);
   U160 : INV_X1 port map( A => A(7), ZN => n102);
   U161 : INV_X1 port map( A => B(0), ZN => n127);
   U162 : INV_X1 port map( A => A(9), ZN => n104);
   U163 : INV_X1 port map( A => FUNC(1), ZN => n161);
   U164 : INV_X1 port map( A => B(3), ZN => n130);
   U165 : INV_X1 port map( A => A(6), ZN => n101);
   U166 : INV_X1 port map( A => A(13), ZN => n108);
   U167 : INV_X1 port map( A => FUNC(0), ZN => n159);
   U168 : INV_X1 port map( A => B(1), ZN => n128);
   U169 : INV_X1 port map( A => A(11), ZN => n106);
   U170 : INV_X1 port map( A => A(15), ZN => n110);
   U171 : INV_X1 port map( A => A(4), ZN => n99);
   U172 : INV_X1 port map( A => B(2), ZN => n129);
   U173 : INV_X1 port map( A => B(5), ZN => n132);
   U174 : INV_X1 port map( A => A(28), ZN => n123);
   U175 : INV_X1 port map( A => A(10), ZN => n105);
   U176 : INV_X1 port map( A => B(7), ZN => n134);
   U177 : INV_X1 port map( A => A(17), ZN => n112);
   U178 : INV_X1 port map( A => A(16), ZN => n111);
   U179 : INV_X1 port map( A => A(12), ZN => n107);
   U180 : INV_X1 port map( A => A(14), ZN => n109);
   U181 : INV_X1 port map( A => A(21), ZN => n116);
   U182 : INV_X1 port map( A => A(8), ZN => n103);
   U183 : INV_X1 port map( A => A(19), ZN => n114);
   U184 : INV_X1 port map( A => B(4), ZN => n131);
   U185 : INV_X1 port map( A => B(6), ZN => n133);
   U186 : INV_X1 port map( A => A(20), ZN => n115);
   U187 : INV_X1 port map( A => A(23), ZN => n118);
   U188 : INV_X1 port map( A => B(9), ZN => n136);
   U189 : INV_X1 port map( A => B(11), ZN => n138);
   U190 : INV_X1 port map( A => A(24), ZN => n119);
   U191 : INV_X1 port map( A => B(13), ZN => n140);
   U192 : INV_X1 port map( A => B(28), ZN => n155);
   U193 : INV_X1 port map( A => A(18), ZN => n113);
   U194 : INV_X1 port map( A => B(15), ZN => n142);
   U195 : INV_X1 port map( A => B(8), ZN => n135);
   U196 : INV_X1 port map( A => B(16), ZN => n143);
   U197 : INV_X1 port map( A => B(12), ZN => n139);
   U198 : INV_X1 port map( A => A(22), ZN => n117);
   U199 : INV_X1 port map( A => B(10), ZN => n137);
   U200 : INV_X1 port map( A => B(20), ZN => n147);
   U201 : INV_X1 port map( A => B(14), ZN => n141);
   U202 : INV_X1 port map( A => B(17), ZN => n144);
   U203 : INV_X1 port map( A => A(29), ZN => n124);
   U204 : INV_X1 port map( A => B(19), ZN => n146);
   U205 : INV_X1 port map( A => A(25), ZN => n120);
   U207 : INV_X1 port map( A => B(24), ZN => n151);
   U208 : INV_X1 port map( A => B(21), ZN => n148);
   U209 : INV_X1 port map( A => B(23), ZN => n150);
   U210 : INV_X1 port map( A => A(27), ZN => n122);
   U211 : INV_X1 port map( A => B(18), ZN => n145);
   U212 : INV_X1 port map( A => B(22), ZN => n149);
   U213 : INV_X1 port map( A => A(26), ZN => n121);
   U214 : INV_X1 port map( A => B(29), ZN => n156);
   U215 : INV_X1 port map( A => B(25), ZN => n152);
   U216 : INV_X1 port map( A => B(27), ZN => n154);
   U217 : INV_X1 port map( A => B(26), ZN => n153);
   U218 : INV_X1 port map( A => A(30), ZN => n125);
   U219 : INV_X1 port map( A => B(30), ZN => n157);
   U220 : INV_X1 port map( A => A(31), ZN => n126);
   U221 : INV_X1 port map( A => B(31), ZN => n158);
   U222 : BUF_X1 port map( A => n73, Z => n77);
   U223 : NAND2_X1 port map( A1 => n159, A2 => n75, ZN => n73);
   U224 : OAI21_X1 port map( B1 => FUNC(3), B2 => n161, A => FUNC(2), ZN => n75
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity comparator_bits32 is

   port( Cout, EN : in std_logic;  func : in std_logic_vector (0 to 3);  sum : 
         in std_logic_vector (31 downto 0);  set : out std_logic_vector (31 
         downto 0));

end comparator_bits32;

architecture SYN_BEHAVIORAL of comparator_bits32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, set_0_port, n5, n6, n7, n8, n9, n10, n13, n14, n15, 
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26 : std_logic;

begin
   set <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, set_0_port 
      );
   
   X_Logic0_port <= '0';
   U20 : OAI33_X1 port map( A1 => n6, A2 => n7, A3 => n23, B1 => n8, B2 => n25,
                           B3 => n24, ZN => n5);
   U21 : NAND3_X1 port map( A1 => n9, A2 => n23, A3 => func(3), ZN => n8);
   U22 : XOR2_X1 port map( A => n10, B => Cout, Z => n7);
   U2 : NOR4_X1 port map( A1 => sum(9), A2 => sum(8), A3 => sum(7), A4 => 
                           sum(6), ZN => n20);
   U3 : OR2_X1 port map( A1 => n21, A2 => n22, ZN => n9);
   U4 : NAND4_X1 port map( A1 => n17, A2 => n18, A3 => n19, A4 => n20, ZN => 
                           n21);
   U5 : NAND4_X1 port map( A1 => n13, A2 => n14, A3 => n15, A4 => n16, ZN => 
                           n22);
   U6 : NOR4_X1 port map( A1 => sum(1), A2 => sum(19), A3 => sum(18), A4 => 
                           sum(17), ZN => n15);
   U7 : NOR4_X1 port map( A1 => sum(23), A2 => sum(22), A3 => sum(21), A4 => 
                           sum(20), ZN => n16);
   U8 : NAND2_X1 port map( A1 => n26, A2 => n9, ZN => n10);
   U9 : AND2_X1 port map( A1 => EN, A2 => n5, ZN => set_0_port);
   U10 : NAND2_X1 port map( A1 => n25, A2 => n24, ZN => n6);
   U11 : NOR4_X1 port map( A1 => sum(5), A2 => sum(4), A3 => sum(3), A4 => 
                           sum(31), ZN => n19);
   U12 : NOR4_X1 port map( A1 => sum(30), A2 => sum(2), A3 => sum(29), A4 => 
                           sum(28), ZN => n18);
   U13 : NOR4_X1 port map( A1 => sum(27), A2 => sum(26), A3 => sum(25), A4 => 
                           sum(24), ZN => n17);
   U14 : NOR4_X1 port map( A1 => sum(16), A2 => sum(15), A3 => sum(14), A4 => 
                           sum(13), ZN => n14);
   U15 : NOR4_X1 port map( A1 => sum(12), A2 => sum(11), A3 => sum(10), A4 => 
                           sum(0), ZN => n13);
   U16 : INV_X1 port map( A => func(3), ZN => n26);
   U17 : INV_X1 port map( A => func(1), ZN => n24);
   U18 : INV_X1 port map( A => func(2), ZN => n25);
   U19 : INV_X1 port map( A => func(0), ZN => n23);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity outputSelect_nbits32 is

   port( FUNC : in std_logic_vector (0 to 3);  p4_out, LS_OUT, comp_out : in 
         std_logic_vector (31 downto 0);  outputSel : out std_logic_vector (31 
         downto 0));

end outputSelect_nbits32;

architecture SYN_BEHAVIORAL of outputSelect_nbits32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n120, n121, n122 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => n38, Z => n83);
   U3 : BUF_X1 port map( A => n39, Z => n76);
   U4 : BUF_X1 port map( A => n37, Z => n87);
   U5 : BUF_X1 port map( A => n83, Z => n81);
   U6 : BUF_X1 port map( A => n87, Z => n85);
   U7 : BUF_X1 port map( A => n87, Z => n86);
   U8 : BUF_X1 port map( A => n87, Z => n84);
   U9 : BUF_X1 port map( A => n76, Z => n79);
   U10 : BUF_X1 port map( A => n76, Z => n78);
   U11 : BUF_X1 port map( A => n76, Z => n77);
   U12 : BUF_X1 port map( A => n83, Z => n80);
   U13 : BUF_X1 port map( A => n83, Z => n82);
   U14 : INV_X1 port map( A => n55, ZN => outputSel(0));
   U15 : AOI222_X1 port map( A1 => p4_out(0), A2 => n85, B1 => comp_out(0), B2 
                           => n81, C1 => LS_OUT(0), C2 => n78, ZN => n55);
   U16 : INV_X1 port map( A => n65, ZN => outputSel(20));
   U17 : AOI222_X1 port map( A1 => p4_out(20), A2 => n84, B1 => comp_out(20), 
                           B2 => n80, C1 => LS_OUT(20), C2 => n77, ZN => n65);
   U18 : INV_X1 port map( A => n67, ZN => outputSel(24));
   U19 : AOI222_X1 port map( A1 => p4_out(24), A2 => n84, B1 => comp_out(24), 
                           B2 => n80, C1 => LS_OUT(24), C2 => n77, ZN => n67);
   U20 : INV_X1 port map( A => n69, ZN => outputSel(28));
   U21 : AOI222_X1 port map( A1 => p4_out(28), A2 => n84, B1 => comp_out(28), 
                           B2 => n80, C1 => LS_OUT(28), C2 => n77, ZN => n69);
   U22 : INV_X1 port map( A => n68, ZN => outputSel(31));
   U23 : AOI222_X1 port map( A1 => p4_out(31), A2 => n84, B1 => comp_out(31), 
                           B2 => n80, C1 => LS_OUT(31), C2 => n77, ZN => n68);
   U24 : INV_X1 port map( A => n47, ZN => outputSel(21));
   U25 : AOI222_X1 port map( A1 => p4_out(21), A2 => n85, B1 => comp_out(21), 
                           B2 => n81, C1 => LS_OUT(21), C2 => n78, ZN => n47);
   U26 : INV_X1 port map( A => n49, ZN => outputSel(25));
   U27 : AOI222_X1 port map( A1 => p4_out(25), A2 => n85, B1 => comp_out(25), 
                           B2 => n81, C1 => LS_OUT(25), C2 => n78, ZN => n49);
   U28 : INV_X1 port map( A => n51, ZN => outputSel(29));
   U29 : AOI222_X1 port map( A1 => p4_out(29), A2 => n85, B1 => comp_out(29), 
                           B2 => n81, C1 => LS_OUT(29), C2 => n78, ZN => n51);
   U30 : INV_X1 port map( A => n48, ZN => outputSel(22));
   U31 : AOI222_X1 port map( A1 => p4_out(22), A2 => n85, B1 => comp_out(22), 
                           B2 => n81, C1 => LS_OUT(22), C2 => n78, ZN => n48);
   U32 : INV_X1 port map( A => n50, ZN => outputSel(26));
   U33 : AOI222_X1 port map( A1 => p4_out(26), A2 => n85, B1 => comp_out(26), 
                           B2 => n81, C1 => LS_OUT(26), C2 => n78, ZN => n50);
   U34 : INV_X1 port map( A => n64, ZN => outputSel(23));
   U35 : AOI222_X1 port map( A1 => p4_out(23), A2 => n84, B1 => comp_out(23), 
                           B2 => n80, C1 => LS_OUT(23), C2 => n77, ZN => n64);
   U36 : INV_X1 port map( A => n66, ZN => outputSel(27));
   U37 : AOI222_X1 port map( A1 => p4_out(27), A2 => n84, B1 => comp_out(27), 
                           B2 => n80, C1 => LS_OUT(27), C2 => n77, ZN => n66);
   U38 : INV_X1 port map( A => n52, ZN => outputSel(30));
   U39 : AOI222_X1 port map( A1 => p4_out(30), A2 => n85, B1 => comp_out(30), 
                           B2 => n81, C1 => LS_OUT(30), C2 => n78, ZN => n52);
   U40 : INV_X1 port map( A => n45, ZN => outputSel(17));
   U41 : AOI222_X1 port map( A1 => p4_out(17), A2 => n86, B1 => comp_out(17), 
                           B2 => n82, C1 => LS_OUT(17), C2 => n79, ZN => n45);
   U42 : INV_X1 port map( A => n46, ZN => outputSel(18));
   U43 : AOI222_X1 port map( A1 => p4_out(18), A2 => n86, B1 => comp_out(18), 
                           B2 => n82, C1 => LS_OUT(18), C2 => n79, ZN => n46);
   U44 : INV_X1 port map( A => n62, ZN => outputSel(19));
   U45 : AOI222_X1 port map( A1 => p4_out(19), A2 => n84, B1 => comp_out(19), 
                           B2 => n80, C1 => LS_OUT(19), C2 => n77, ZN => n62);
   U46 : INV_X1 port map( A => n63, ZN => outputSel(16));
   U47 : AOI222_X1 port map( A1 => p4_out(16), A2 => n84, B1 => comp_out(16), 
                           B2 => n80, C1 => LS_OUT(16), C2 => n77, ZN => n63);
   U48 : INV_X1 port map( A => n60, ZN => outputSel(15));
   U49 : AOI222_X1 port map( A1 => p4_out(15), A2 => n84, B1 => comp_out(15), 
                           B2 => n80, C1 => LS_OUT(15), C2 => n77, ZN => n60);
   U50 : INV_X1 port map( A => n56, ZN => outputSel(7));
   U51 : AOI222_X1 port map( A1 => p4_out(7), A2 => n85, B1 => comp_out(7), B2 
                           => n81, C1 => LS_OUT(7), C2 => n78, ZN => n56);
   U52 : INV_X1 port map( A => n43, ZN => outputSel(13));
   U53 : AOI222_X1 port map( A1 => p4_out(13), A2 => n86, B1 => comp_out(13), 
                           B2 => n82, C1 => LS_OUT(13), C2 => n79, ZN => n43);
   U54 : INV_X1 port map( A => n58, ZN => outputSel(11));
   U55 : AOI222_X1 port map( A1 => p4_out(11), A2 => n85, B1 => comp_out(11), 
                           B2 => n81, C1 => LS_OUT(11), C2 => n78, ZN => n58);
   U56 : INV_X1 port map( A => n44, ZN => outputSel(14));
   U57 : AOI222_X1 port map( A1 => p4_out(14), A2 => n86, B1 => comp_out(14), 
                           B2 => n82, C1 => LS_OUT(14), C2 => n79, ZN => n44);
   U58 : INV_X1 port map( A => n61, ZN => outputSel(12));
   U59 : AOI222_X1 port map( A1 => p4_out(12), A2 => n84, B1 => comp_out(12), 
                           B2 => n80, C1 => LS_OUT(12), C2 => n77, ZN => n61);
   U60 : INV_X1 port map( A => n53, ZN => outputSel(3));
   U61 : AOI222_X1 port map( A1 => p4_out(3), A2 => n85, B1 => comp_out(3), B2 
                           => n81, C1 => LS_OUT(3), C2 => n78, ZN => n53);
   U62 : INV_X1 port map( A => n42, ZN => outputSel(10));
   U63 : AOI222_X1 port map( A1 => p4_out(10), A2 => n86, B1 => comp_out(10), 
                           B2 => n82, C1 => LS_OUT(10), C2 => n79, ZN => n42);
   U64 : INV_X1 port map( A => n59, ZN => outputSel(8));
   U65 : AOI222_X1 port map( A1 => p4_out(8), A2 => n84, B1 => comp_out(8), B2 
                           => n80, C1 => LS_OUT(8), C2 => n77, ZN => n59);
   U66 : INV_X1 port map( A => n41, ZN => outputSel(9));
   U67 : AOI222_X1 port map( A1 => p4_out(9), A2 => n86, B1 => comp_out(9), B2 
                           => n82, C1 => LS_OUT(9), C2 => n79, ZN => n41);
   U68 : INV_X1 port map( A => n40, ZN => outputSel(6));
   U69 : AOI222_X1 port map( A1 => p4_out(6), A2 => n86, B1 => comp_out(6), B2 
                           => n82, C1 => LS_OUT(6), C2 => n79, ZN => n40);
   U70 : INV_X1 port map( A => n70, ZN => outputSel(2));
   U71 : AOI222_X1 port map( A1 => p4_out(2), A2 => n84, B1 => comp_out(2), B2 
                           => n80, C1 => LS_OUT(2), C2 => n77, ZN => n70);
   U72 : INV_X1 port map( A => n57, ZN => outputSel(4));
   U73 : AOI222_X1 port map( A1 => p4_out(4), A2 => n85, B1 => comp_out(4), B2 
                           => n81, C1 => LS_OUT(4), C2 => n78, ZN => n57);
   U74 : INV_X1 port map( A => n36, ZN => outputSel(5));
   U75 : AOI222_X1 port map( A1 => p4_out(5), A2 => n86, B1 => comp_out(5), B2 
                           => n82, C1 => LS_OUT(5), C2 => n79, ZN => n36);
   U76 : INV_X1 port map( A => n54, ZN => outputSel(1));
   U77 : AOI222_X1 port map( A1 => p4_out(1), A2 => n85, B1 => comp_out(1), B2 
                           => n81, C1 => LS_OUT(1), C2 => n78, ZN => n54);
   U78 : INV_X1 port map( A => FUNC(2), ZN => n122);
   U79 : AOI221_X1 port map( B1 => n120, B2 => n122, C1 => n121, C2 => FUNC(2),
                           A => n72, ZN => n38);
   U80 : AOI21_X1 port map( B1 => n120, B2 => FUNC(3), A => n121, ZN => n72);
   U81 : INV_X1 port map( A => FUNC(1), ZN => n121);
   U82 : INV_X1 port map( A => FUNC(0), ZN => n120);
   U83 : NOR3_X1 port map( A1 => FUNC(1), A2 => FUNC(0), A3 => n122, ZN => n37)
                           ;
   U84 : AND2_X1 port map( A1 => n71, A2 => n120, ZN => n39);
   U85 : OAI21_X1 port map( B1 => FUNC(3), B2 => n121, A => FUNC(2), ZN => n71)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_352 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_352;

architecture SYN_ASYNCH_FD of FD_352 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   Q_reg : SDFFR_X1 port map( D => n6, SI => n7, SE => n5, CK => CK, RN => n2, 
                           Q => Q, QN => n4);
   U2 : OAI21_X1 port map( B1 => n4, B2 => ENABLE, A => n3, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D, A2 => ENABLE, ZN => n3);
   U4 : INV_X1 port map( A => n1, ZN => n5);
   n6 <= '1';
   n7 <= '0';
   U7 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_2;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n33, n66, n67, n68, n69, n70 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n70, Z => n69);
   U2 : INV_X1 port map( A => n70, ZN => n68);
   U3 : BUF_X1 port map( A => n69, Z => n33);
   U4 : BUF_X1 port map( A => n69, Z => n67);
   U5 : BUF_X1 port map( A => n69, Z => n66);
   U6 : INV_X1 port map( A => n42, ZN => Y(30));
   U7 : AOI22_X1 port map( A1 => A(30), A2 => n68, B1 => B(30), B2 => n66, ZN 
                           => n42);
   U8 : INV_X1 port map( A => n44, ZN => Y(29));
   U9 : AOI22_X1 port map( A1 => A(29), A2 => n68, B1 => B(29), B2 => n66, ZN 
                           => n44);
   U10 : INV_X1 port map( A => n45, ZN => Y(28));
   U11 : AOI22_X1 port map( A1 => A(28), A2 => n68, B1 => B(28), B2 => n66, ZN 
                           => n45);
   U12 : INV_X1 port map( A => n46, ZN => Y(27));
   U13 : AOI22_X1 port map( A1 => A(27), A2 => n68, B1 => B(27), B2 => n66, ZN 
                           => n46);
   U14 : INV_X1 port map( A => n47, ZN => Y(26));
   U15 : AOI22_X1 port map( A1 => A(26), A2 => S, B1 => B(26), B2 => n66, ZN =>
                           n47);
   U16 : INV_X1 port map( A => n48, ZN => Y(25));
   U17 : AOI22_X1 port map( A1 => A(25), A2 => S, B1 => B(25), B2 => n66, ZN =>
                           n48);
   U18 : INV_X1 port map( A => n49, ZN => Y(24));
   U19 : AOI22_X1 port map( A1 => A(24), A2 => S, B1 => B(24), B2 => n66, ZN =>
                           n49);
   U20 : INV_X1 port map( A => n50, ZN => Y(23));
   U21 : AOI22_X1 port map( A1 => A(23), A2 => S, B1 => B(23), B2 => n66, ZN =>
                           n50);
   U22 : INV_X1 port map( A => n51, ZN => Y(22));
   U23 : AOI22_X1 port map( A1 => A(22), A2 => S, B1 => B(22), B2 => n66, ZN =>
                           n51);
   U24 : INV_X1 port map( A => n52, ZN => Y(21));
   U25 : AOI22_X1 port map( A1 => A(21), A2 => S, B1 => B(21), B2 => n66, ZN =>
                           n52);
   U26 : INV_X1 port map( A => n53, ZN => Y(20));
   U27 : AOI22_X1 port map( A1 => A(20), A2 => S, B1 => B(20), B2 => n66, ZN =>
                           n53);
   U28 : INV_X1 port map( A => n55, ZN => Y(19));
   U29 : AOI22_X1 port map( A1 => A(19), A2 => n68, B1 => B(19), B2 => n33, ZN 
                           => n55);
   U30 : INV_X1 port map( A => n56, ZN => Y(18));
   U31 : AOI22_X1 port map( A1 => A(18), A2 => n68, B1 => B(18), B2 => n33, ZN 
                           => n56);
   U32 : INV_X1 port map( A => n57, ZN => Y(17));
   U33 : AOI22_X1 port map( A1 => A(17), A2 => n68, B1 => B(17), B2 => n33, ZN 
                           => n57);
   U34 : INV_X1 port map( A => n58, ZN => Y(16));
   U35 : AOI22_X1 port map( A1 => A(16), A2 => n68, B1 => B(16), B2 => n33, ZN 
                           => n58);
   U36 : INV_X1 port map( A => n59, ZN => Y(15));
   U37 : AOI22_X1 port map( A1 => A(15), A2 => n68, B1 => B(15), B2 => n33, ZN 
                           => n59);
   U38 : INV_X1 port map( A => n60, ZN => Y(14));
   U39 : AOI22_X1 port map( A1 => A(14), A2 => n68, B1 => B(14), B2 => n33, ZN 
                           => n60);
   U40 : INV_X1 port map( A => n61, ZN => Y(13));
   U41 : AOI22_X1 port map( A1 => A(13), A2 => n68, B1 => B(13), B2 => n33, ZN 
                           => n61);
   U42 : AOI22_X1 port map( A1 => A(0), A2 => n68, B1 => B(0), B2 => n33, ZN =>
                           n65);
   U43 : INV_X1 port map( A => n65, ZN => Y(0));
   U44 : INV_X1 port map( A => S, ZN => n70);
   U45 : INV_X1 port map( A => n62, ZN => Y(12));
   U46 : AOI22_X1 port map( A1 => A(12), A2 => n68, B1 => B(12), B2 => n33, ZN 
                           => n62);
   U47 : INV_X1 port map( A => n40, ZN => Y(3));
   U48 : AOI22_X1 port map( A1 => A(3), A2 => S, B1 => B(3), B2 => n67, ZN => 
                           n40);
   U49 : INV_X1 port map( A => n39, ZN => Y(4));
   U50 : AOI22_X1 port map( A1 => A(4), A2 => S, B1 => B(4), B2 => n67, ZN => 
                           n39);
   U51 : INV_X1 port map( A => n38, ZN => Y(5));
   U52 : AOI22_X1 port map( A1 => A(5), A2 => S, B1 => B(5), B2 => n67, ZN => 
                           n38);
   U53 : INV_X1 port map( A => n37, ZN => Y(6));
   U54 : AOI22_X1 port map( A1 => A(6), A2 => S, B1 => B(6), B2 => n67, ZN => 
                           n37);
   U55 : INV_X1 port map( A => n36, ZN => Y(7));
   U56 : AOI22_X1 port map( A1 => A(7), A2 => S, B1 => B(7), B2 => n67, ZN => 
                           n36);
   U57 : INV_X1 port map( A => n35, ZN => Y(8));
   U58 : AOI22_X1 port map( A1 => A(8), A2 => S, B1 => B(8), B2 => n67, ZN => 
                           n35);
   U59 : INV_X1 port map( A => n54, ZN => Y(1));
   U60 : AOI22_X1 port map( A1 => A(1), A2 => n68, B1 => B(1), B2 => n33, ZN =>
                           n54);
   U61 : INV_X1 port map( A => n43, ZN => Y(2));
   U62 : AOI22_X1 port map( A1 => A(2), A2 => S, B1 => B(2), B2 => n66, ZN => 
                           n43);
   U63 : INV_X1 port map( A => n64, ZN => Y(10));
   U64 : AOI22_X1 port map( A1 => A(10), A2 => n68, B1 => B(10), B2 => n33, ZN 
                           => n64);
   U65 : INV_X1 port map( A => n63, ZN => Y(11));
   U66 : AOI22_X1 port map( A1 => A(11), A2 => n68, B1 => B(11), B2 => n33, ZN 
                           => n63);
   U67 : INV_X1 port map( A => n34, ZN => Y(9));
   U68 : AOI22_X1 port map( A1 => S, A2 => A(9), B1 => B(9), B2 => n67, ZN => 
                           n34);
   U69 : AOI22_X1 port map( A1 => A(31), A2 => S, B1 => B(31), B2 => n67, ZN =>
                           n41);
   U70 : INV_X1 port map( A => n41, ZN => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21;

architecture SYN_BEHAVIORAL of MUX21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Y);
   U2 : AOI22_X1 port map( A1 => S, A2 => A, B1 => B, B2 => n4, ZN => n3);
   U3 : INV_X1 port map( A => S, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_0 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_0;

architecture SYN_ASYNCH_FD of FD_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n3, n4, n1, n2 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CK, RN => n3, Q => Q, QN => n2);
   U2 : OAI21_X1 port map( B1 => n2, B2 => ENABLE, A => n1, ZN => n4);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D, ZN => n1);
   U4 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n3);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity XNOR_logic is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR_logic;

architecture SYN_BEHAVIORAL of XNOR_logic is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity alu_nbits32 is

   port( FUNC : in std_logic_vector (0 to 3);  A, B : in std_logic_vector (31 
         downto 0);  OUTALU : out std_logic_vector (31 downto 0));

end alu_nbits32;

architecture SYN_STRUCTURAL of alu_nbits32 is

   component logic_and_shift_N32
      port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4_ADDER_NBITS32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component ctrl_alu_NBITS32
      port( A, B : in std_logic_vector (31 downto 0);  FUNC : in 
            std_logic_vector (0 to 3);  Ap4, Bp4 : out std_logic_vector (31 
            downto 0);  Cin : out std_logic;  Als, Bls : out std_logic_vector 
            (31 downto 0);  enableComp : out std_logic);
   end component;
   
   component comparator_bits32
      port( Cout, EN : in std_logic;  func : in std_logic_vector (0 to 3);  sum
            : in std_logic_vector (31 downto 0);  set : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component outputSelect_nbits32
      port( FUNC : in std_logic_vector (0 to 3);  p4_out, LS_OUT, comp_out : in
            std_logic_vector (31 downto 0);  outputSel : out std_logic_vector 
            (31 downto 0));
   end component;
   
   signal p4_outsig_31_port, p4_outsig_30_port, p4_outsig_29_port, 
      p4_outsig_28_port, p4_outsig_27_port, p4_outsig_26_port, 
      p4_outsig_25_port, p4_outsig_24_port, p4_outsig_23_port, 
      p4_outsig_22_port, p4_outsig_21_port, p4_outsig_20_port, 
      p4_outsig_19_port, p4_outsig_18_port, p4_outsig_17_port, 
      p4_outsig_16_port, p4_outsig_15_port, p4_outsig_14_port, 
      p4_outsig_13_port, p4_outsig_12_port, p4_outsig_11_port, 
      p4_outsig_10_port, p4_outsig_9_port, p4_outsig_8_port, p4_outsig_7_port, 
      p4_outsig_6_port, p4_outsig_5_port, p4_outsig_4_port, p4_outsig_3_port, 
      p4_outsig_2_port, p4_outsig_1_port, p4_outsig_0_port, LS_OUTsig_31_port, 
      LS_OUTsig_30_port, LS_OUTsig_29_port, LS_OUTsig_28_port, 
      LS_OUTsig_27_port, LS_OUTsig_26_port, LS_OUTsig_25_port, 
      LS_OUTsig_24_port, LS_OUTsig_23_port, LS_OUTsig_22_port, 
      LS_OUTsig_21_port, LS_OUTsig_20_port, LS_OUTsig_19_port, 
      LS_OUTsig_18_port, LS_OUTsig_17_port, LS_OUTsig_16_port, 
      LS_OUTsig_15_port, LS_OUTsig_14_port, LS_OUTsig_13_port, 
      LS_OUTsig_12_port, LS_OUTsig_11_port, LS_OUTsig_10_port, LS_OUTsig_9_port
      , LS_OUTsig_8_port, LS_OUTsig_7_port, LS_OUTsig_6_port, LS_OUTsig_5_port,
      LS_OUTsig_4_port, LS_OUTsig_3_port, LS_OUTsig_2_port, LS_OUTsig_1_port, 
      LS_OUTsig_0_port, comp_outsig_31_port, comp_outsig_30_port, 
      comp_outsig_29_port, comp_outsig_28_port, comp_outsig_27_port, 
      comp_outsig_26_port, comp_outsig_25_port, comp_outsig_24_port, 
      comp_outsig_23_port, comp_outsig_22_port, comp_outsig_21_port, 
      comp_outsig_20_port, comp_outsig_19_port, comp_outsig_18_port, 
      comp_outsig_17_port, comp_outsig_16_port, comp_outsig_15_port, 
      comp_outsig_14_port, comp_outsig_13_port, comp_outsig_12_port, 
      comp_outsig_11_port, comp_outsig_10_port, comp_outsig_9_port, 
      comp_outsig_8_port, comp_outsig_7_port, comp_outsig_6_port, 
      comp_outsig_5_port, comp_outsig_4_port, comp_outsig_3_port, 
      comp_outsig_2_port, comp_outsig_1_port, comp_outsig_0_port, p4_comp_Co, 
      enable_Comp, p4_ctrl_A_31_port, p4_ctrl_A_30_port, p4_ctrl_A_29_port, 
      p4_ctrl_A_28_port, p4_ctrl_A_27_port, p4_ctrl_A_26_port, 
      p4_ctrl_A_25_port, p4_ctrl_A_24_port, p4_ctrl_A_23_port, 
      p4_ctrl_A_22_port, p4_ctrl_A_21_port, p4_ctrl_A_20_port, 
      p4_ctrl_A_19_port, p4_ctrl_A_18_port, p4_ctrl_A_17_port, 
      p4_ctrl_A_16_port, p4_ctrl_A_15_port, p4_ctrl_A_14_port, 
      p4_ctrl_A_13_port, p4_ctrl_A_12_port, p4_ctrl_A_11_port, 
      p4_ctrl_A_10_port, p4_ctrl_A_9_port, p4_ctrl_A_8_port, p4_ctrl_A_7_port, 
      p4_ctrl_A_6_port, p4_ctrl_A_5_port, p4_ctrl_A_4_port, p4_ctrl_A_3_port, 
      p4_ctrl_A_2_port, p4_ctrl_A_1_port, p4_ctrl_A_0_port, p4_ctrl_B_31_port, 
      p4_ctrl_B_30_port, p4_ctrl_B_29_port, p4_ctrl_B_28_port, 
      p4_ctrl_B_27_port, p4_ctrl_B_26_port, p4_ctrl_B_25_port, 
      p4_ctrl_B_24_port, p4_ctrl_B_23_port, p4_ctrl_B_22_port, 
      p4_ctrl_B_21_port, p4_ctrl_B_20_port, p4_ctrl_B_19_port, 
      p4_ctrl_B_18_port, p4_ctrl_B_17_port, p4_ctrl_B_16_port, 
      p4_ctrl_B_15_port, p4_ctrl_B_14_port, p4_ctrl_B_13_port, 
      p4_ctrl_B_12_port, p4_ctrl_B_11_port, p4_ctrl_B_10_port, p4_ctrl_B_9_port
      , p4_ctrl_B_8_port, p4_ctrl_B_7_port, p4_ctrl_B_6_port, p4_ctrl_B_5_port,
      p4_ctrl_B_4_port, p4_ctrl_B_3_port, p4_ctrl_B_2_port, p4_ctrl_B_1_port, 
      p4_ctrl_B_0_port, p4_ctrl_Cin, ctrl_LS_A_31_port, ctrl_LS_A_30_port, 
      ctrl_LS_A_29_port, ctrl_LS_A_28_port, ctrl_LS_A_27_port, 
      ctrl_LS_A_26_port, ctrl_LS_A_25_port, ctrl_LS_A_24_port, 
      ctrl_LS_A_23_port, ctrl_LS_A_22_port, ctrl_LS_A_21_port, 
      ctrl_LS_A_20_port, ctrl_LS_A_19_port, ctrl_LS_A_18_port, 
      ctrl_LS_A_17_port, ctrl_LS_A_16_port, ctrl_LS_A_15_port, 
      ctrl_LS_A_14_port, ctrl_LS_A_13_port, ctrl_LS_A_12_port, 
      ctrl_LS_A_11_port, ctrl_LS_A_10_port, ctrl_LS_A_9_port, ctrl_LS_A_8_port,
      ctrl_LS_A_7_port, ctrl_LS_A_6_port, ctrl_LS_A_5_port, ctrl_LS_A_4_port, 
      ctrl_LS_A_3_port, ctrl_LS_A_2_port, ctrl_LS_A_1_port, ctrl_LS_A_0_port, 
      ctrl_LS_B_31_port, ctrl_LS_B_30_port, ctrl_LS_B_29_port, 
      ctrl_LS_B_28_port, ctrl_LS_B_27_port, ctrl_LS_B_26_port, 
      ctrl_LS_B_25_port, ctrl_LS_B_24_port, ctrl_LS_B_23_port, 
      ctrl_LS_B_22_port, ctrl_LS_B_21_port, ctrl_LS_B_20_port, 
      ctrl_LS_B_19_port, ctrl_LS_B_18_port, ctrl_LS_B_17_port, 
      ctrl_LS_B_16_port, ctrl_LS_B_15_port, ctrl_LS_B_14_port, 
      ctrl_LS_B_13_port, ctrl_LS_B_12_port, ctrl_LS_B_11_port, 
      ctrl_LS_B_10_port, ctrl_LS_B_9_port, ctrl_LS_B_8_port, ctrl_LS_B_7_port, 
      ctrl_LS_B_6_port, ctrl_LS_B_5_port, ctrl_LS_B_4_port, ctrl_LS_B_3_port, 
      ctrl_LS_B_2_port, ctrl_LS_B_1_port, ctrl_LS_B_0_port, n_1020, n_1021, 
      n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, 
      n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, 
      n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, 
      n_1049, n_1050 : std_logic;

begin
   
   comp_outsig_1_port <= '0';
   comp_outsig_2_port <= '0';
   comp_outsig_3_port <= '0';
   comp_outsig_4_port <= '0';
   comp_outsig_5_port <= '0';
   comp_outsig_6_port <= '0';
   comp_outsig_7_port <= '0';
   comp_outsig_8_port <= '0';
   comp_outsig_9_port <= '0';
   comp_outsig_10_port <= '0';
   comp_outsig_11_port <= '0';
   comp_outsig_12_port <= '0';
   comp_outsig_13_port <= '0';
   comp_outsig_14_port <= '0';
   comp_outsig_15_port <= '0';
   comp_outsig_16_port <= '0';
   comp_outsig_17_port <= '0';
   comp_outsig_18_port <= '0';
   comp_outsig_19_port <= '0';
   comp_outsig_20_port <= '0';
   comp_outsig_21_port <= '0';
   comp_outsig_22_port <= '0';
   comp_outsig_23_port <= '0';
   comp_outsig_24_port <= '0';
   comp_outsig_25_port <= '0';
   comp_outsig_26_port <= '0';
   comp_outsig_27_port <= '0';
   comp_outsig_28_port <= '0';
   comp_outsig_29_port <= '0';
   comp_outsig_30_port <= '0';
   comp_outsig_31_port <= '0';
   SELOUT : outputSelect_nbits32 port map( FUNC(0) => FUNC(0), FUNC(1) => 
                           FUNC(1), FUNC(2) => FUNC(2), FUNC(3) => FUNC(3), 
                           p4_out(31) => p4_outsig_31_port, p4_out(30) => 
                           p4_outsig_30_port, p4_out(29) => p4_outsig_29_port, 
                           p4_out(28) => p4_outsig_28_port, p4_out(27) => 
                           p4_outsig_27_port, p4_out(26) => p4_outsig_26_port, 
                           p4_out(25) => p4_outsig_25_port, p4_out(24) => 
                           p4_outsig_24_port, p4_out(23) => p4_outsig_23_port, 
                           p4_out(22) => p4_outsig_22_port, p4_out(21) => 
                           p4_outsig_21_port, p4_out(20) => p4_outsig_20_port, 
                           p4_out(19) => p4_outsig_19_port, p4_out(18) => 
                           p4_outsig_18_port, p4_out(17) => p4_outsig_17_port, 
                           p4_out(16) => p4_outsig_16_port, p4_out(15) => 
                           p4_outsig_15_port, p4_out(14) => p4_outsig_14_port, 
                           p4_out(13) => p4_outsig_13_port, p4_out(12) => 
                           p4_outsig_12_port, p4_out(11) => p4_outsig_11_port, 
                           p4_out(10) => p4_outsig_10_port, p4_out(9) => 
                           p4_outsig_9_port, p4_out(8) => p4_outsig_8_port, 
                           p4_out(7) => p4_outsig_7_port, p4_out(6) => 
                           p4_outsig_6_port, p4_out(5) => p4_outsig_5_port, 
                           p4_out(4) => p4_outsig_4_port, p4_out(3) => 
                           p4_outsig_3_port, p4_out(2) => p4_outsig_2_port, 
                           p4_out(1) => p4_outsig_1_port, p4_out(0) => 
                           p4_outsig_0_port, LS_OUT(31) => LS_OUTsig_31_port, 
                           LS_OUT(30) => LS_OUTsig_30_port, LS_OUT(29) => 
                           LS_OUTsig_29_port, LS_OUT(28) => LS_OUTsig_28_port, 
                           LS_OUT(27) => LS_OUTsig_27_port, LS_OUT(26) => 
                           LS_OUTsig_26_port, LS_OUT(25) => LS_OUTsig_25_port, 
                           LS_OUT(24) => LS_OUTsig_24_port, LS_OUT(23) => 
                           LS_OUTsig_23_port, LS_OUT(22) => LS_OUTsig_22_port, 
                           LS_OUT(21) => LS_OUTsig_21_port, LS_OUT(20) => 
                           LS_OUTsig_20_port, LS_OUT(19) => LS_OUTsig_19_port, 
                           LS_OUT(18) => LS_OUTsig_18_port, LS_OUT(17) => 
                           LS_OUTsig_17_port, LS_OUT(16) => LS_OUTsig_16_port, 
                           LS_OUT(15) => LS_OUTsig_15_port, LS_OUT(14) => 
                           LS_OUTsig_14_port, LS_OUT(13) => LS_OUTsig_13_port, 
                           LS_OUT(12) => LS_OUTsig_12_port, LS_OUT(11) => 
                           LS_OUTsig_11_port, LS_OUT(10) => LS_OUTsig_10_port, 
                           LS_OUT(9) => LS_OUTsig_9_port, LS_OUT(8) => 
                           LS_OUTsig_8_port, LS_OUT(7) => LS_OUTsig_7_port, 
                           LS_OUT(6) => LS_OUTsig_6_port, LS_OUT(5) => 
                           LS_OUTsig_5_port, LS_OUT(4) => LS_OUTsig_4_port, 
                           LS_OUT(3) => LS_OUTsig_3_port, LS_OUT(2) => 
                           LS_OUTsig_2_port, LS_OUT(1) => LS_OUTsig_1_port, 
                           LS_OUT(0) => LS_OUTsig_0_port, comp_out(31) => 
                           comp_outsig_31_port, comp_out(30) => 
                           comp_outsig_30_port, comp_out(29) => 
                           comp_outsig_29_port, comp_out(28) => 
                           comp_outsig_28_port, comp_out(27) => 
                           comp_outsig_27_port, comp_out(26) => 
                           comp_outsig_26_port, comp_out(25) => 
                           comp_outsig_25_port, comp_out(24) => 
                           comp_outsig_24_port, comp_out(23) => 
                           comp_outsig_23_port, comp_out(22) => 
                           comp_outsig_22_port, comp_out(21) => 
                           comp_outsig_21_port, comp_out(20) => 
                           comp_outsig_20_port, comp_out(19) => 
                           comp_outsig_19_port, comp_out(18) => 
                           comp_outsig_18_port, comp_out(17) => 
                           comp_outsig_17_port, comp_out(16) => 
                           comp_outsig_16_port, comp_out(15) => 
                           comp_outsig_15_port, comp_out(14) => 
                           comp_outsig_14_port, comp_out(13) => 
                           comp_outsig_13_port, comp_out(12) => 
                           comp_outsig_12_port, comp_out(11) => 
                           comp_outsig_11_port, comp_out(10) => 
                           comp_outsig_10_port, comp_out(9) => 
                           comp_outsig_9_port, comp_out(8) => 
                           comp_outsig_8_port, comp_out(7) => 
                           comp_outsig_7_port, comp_out(6) => 
                           comp_outsig_6_port, comp_out(5) => 
                           comp_outsig_5_port, comp_out(4) => 
                           comp_outsig_4_port, comp_out(3) => 
                           comp_outsig_3_port, comp_out(2) => 
                           comp_outsig_2_port, comp_out(1) => 
                           comp_outsig_1_port, comp_out(0) => 
                           comp_outsig_0_port, outputSel(31) => OUTALU(31), 
                           outputSel(30) => OUTALU(30), outputSel(29) => 
                           OUTALU(29), outputSel(28) => OUTALU(28), 
                           outputSel(27) => OUTALU(27), outputSel(26) => 
                           OUTALU(26), outputSel(25) => OUTALU(25), 
                           outputSel(24) => OUTALU(24), outputSel(23) => 
                           OUTALU(23), outputSel(22) => OUTALU(22), 
                           outputSel(21) => OUTALU(21), outputSel(20) => 
                           OUTALU(20), outputSel(19) => OUTALU(19), 
                           outputSel(18) => OUTALU(18), outputSel(17) => 
                           OUTALU(17), outputSel(16) => OUTALU(16), 
                           outputSel(15) => OUTALU(15), outputSel(14) => 
                           OUTALU(14), outputSel(13) => OUTALU(13), 
                           outputSel(12) => OUTALU(12), outputSel(11) => 
                           OUTALU(11), outputSel(10) => OUTALU(10), 
                           outputSel(9) => OUTALU(9), outputSel(8) => OUTALU(8)
                           , outputSel(7) => OUTALU(7), outputSel(6) => 
                           OUTALU(6), outputSel(5) => OUTALU(5), outputSel(4) 
                           => OUTALU(4), outputSel(3) => OUTALU(3), 
                           outputSel(2) => OUTALU(2), outputSel(1) => OUTALU(1)
                           , outputSel(0) => OUTALU(0));
   COMP : comparator_bits32 port map( Cout => p4_comp_Co, EN => enable_Comp, 
                           func(0) => FUNC(0), func(1) => FUNC(1), func(2) => 
                           FUNC(2), func(3) => FUNC(3), sum(31) => 
                           p4_outsig_31_port, sum(30) => p4_outsig_30_port, 
                           sum(29) => p4_outsig_29_port, sum(28) => 
                           p4_outsig_28_port, sum(27) => p4_outsig_27_port, 
                           sum(26) => p4_outsig_26_port, sum(25) => 
                           p4_outsig_25_port, sum(24) => p4_outsig_24_port, 
                           sum(23) => p4_outsig_23_port, sum(22) => 
                           p4_outsig_22_port, sum(21) => p4_outsig_21_port, 
                           sum(20) => p4_outsig_20_port, sum(19) => 
                           p4_outsig_19_port, sum(18) => p4_outsig_18_port, 
                           sum(17) => p4_outsig_17_port, sum(16) => 
                           p4_outsig_16_port, sum(15) => p4_outsig_15_port, 
                           sum(14) => p4_outsig_14_port, sum(13) => 
                           p4_outsig_13_port, sum(12) => p4_outsig_12_port, 
                           sum(11) => p4_outsig_11_port, sum(10) => 
                           p4_outsig_10_port, sum(9) => p4_outsig_9_port, 
                           sum(8) => p4_outsig_8_port, sum(7) => 
                           p4_outsig_7_port, sum(6) => p4_outsig_6_port, sum(5)
                           => p4_outsig_5_port, sum(4) => p4_outsig_4_port, 
                           sum(3) => p4_outsig_3_port, sum(2) => 
                           p4_outsig_2_port, sum(1) => p4_outsig_1_port, sum(0)
                           => p4_outsig_0_port, set(31) => n_1020, set(30) => 
                           n_1021, set(29) => n_1022, set(28) => n_1023, 
                           set(27) => n_1024, set(26) => n_1025, set(25) => 
                           n_1026, set(24) => n_1027, set(23) => n_1028, 
                           set(22) => n_1029, set(21) => n_1030, set(20) => 
                           n_1031, set(19) => n_1032, set(18) => n_1033, 
                           set(17) => n_1034, set(16) => n_1035, set(15) => 
                           n_1036, set(14) => n_1037, set(13) => n_1038, 
                           set(12) => n_1039, set(11) => n_1040, set(10) => 
                           n_1041, set(9) => n_1042, set(8) => n_1043, set(7) 
                           => n_1044, set(6) => n_1045, set(5) => n_1046, 
                           set(4) => n_1047, set(3) => n_1048, set(2) => n_1049
                           , set(1) => n_1050, set(0) => comp_outsig_0_port);
   CTRLALU : ctrl_alu_NBITS32 port map( A(31) => A(31), A(30) => A(30), A(29) 
                           => A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), FUNC(0) => FUNC(0), FUNC(1) => FUNC(1), 
                           FUNC(2) => FUNC(2), FUNC(3) => FUNC(3), Ap4(31) => 
                           p4_ctrl_A_31_port, Ap4(30) => p4_ctrl_A_30_port, 
                           Ap4(29) => p4_ctrl_A_29_port, Ap4(28) => 
                           p4_ctrl_A_28_port, Ap4(27) => p4_ctrl_A_27_port, 
                           Ap4(26) => p4_ctrl_A_26_port, Ap4(25) => 
                           p4_ctrl_A_25_port, Ap4(24) => p4_ctrl_A_24_port, 
                           Ap4(23) => p4_ctrl_A_23_port, Ap4(22) => 
                           p4_ctrl_A_22_port, Ap4(21) => p4_ctrl_A_21_port, 
                           Ap4(20) => p4_ctrl_A_20_port, Ap4(19) => 
                           p4_ctrl_A_19_port, Ap4(18) => p4_ctrl_A_18_port, 
                           Ap4(17) => p4_ctrl_A_17_port, Ap4(16) => 
                           p4_ctrl_A_16_port, Ap4(15) => p4_ctrl_A_15_port, 
                           Ap4(14) => p4_ctrl_A_14_port, Ap4(13) => 
                           p4_ctrl_A_13_port, Ap4(12) => p4_ctrl_A_12_port, 
                           Ap4(11) => p4_ctrl_A_11_port, Ap4(10) => 
                           p4_ctrl_A_10_port, Ap4(9) => p4_ctrl_A_9_port, 
                           Ap4(8) => p4_ctrl_A_8_port, Ap4(7) => 
                           p4_ctrl_A_7_port, Ap4(6) => p4_ctrl_A_6_port, Ap4(5)
                           => p4_ctrl_A_5_port, Ap4(4) => p4_ctrl_A_4_port, 
                           Ap4(3) => p4_ctrl_A_3_port, Ap4(2) => 
                           p4_ctrl_A_2_port, Ap4(1) => p4_ctrl_A_1_port, Ap4(0)
                           => p4_ctrl_A_0_port, Bp4(31) => p4_ctrl_B_31_port, 
                           Bp4(30) => p4_ctrl_B_30_port, Bp4(29) => 
                           p4_ctrl_B_29_port, Bp4(28) => p4_ctrl_B_28_port, 
                           Bp4(27) => p4_ctrl_B_27_port, Bp4(26) => 
                           p4_ctrl_B_26_port, Bp4(25) => p4_ctrl_B_25_port, 
                           Bp4(24) => p4_ctrl_B_24_port, Bp4(23) => 
                           p4_ctrl_B_23_port, Bp4(22) => p4_ctrl_B_22_port, 
                           Bp4(21) => p4_ctrl_B_21_port, Bp4(20) => 
                           p4_ctrl_B_20_port, Bp4(19) => p4_ctrl_B_19_port, 
                           Bp4(18) => p4_ctrl_B_18_port, Bp4(17) => 
                           p4_ctrl_B_17_port, Bp4(16) => p4_ctrl_B_16_port, 
                           Bp4(15) => p4_ctrl_B_15_port, Bp4(14) => 
                           p4_ctrl_B_14_port, Bp4(13) => p4_ctrl_B_13_port, 
                           Bp4(12) => p4_ctrl_B_12_port, Bp4(11) => 
                           p4_ctrl_B_11_port, Bp4(10) => p4_ctrl_B_10_port, 
                           Bp4(9) => p4_ctrl_B_9_port, Bp4(8) => 
                           p4_ctrl_B_8_port, Bp4(7) => p4_ctrl_B_7_port, Bp4(6)
                           => p4_ctrl_B_6_port, Bp4(5) => p4_ctrl_B_5_port, 
                           Bp4(4) => p4_ctrl_B_4_port, Bp4(3) => 
                           p4_ctrl_B_3_port, Bp4(2) => p4_ctrl_B_2_port, Bp4(1)
                           => p4_ctrl_B_1_port, Bp4(0) => p4_ctrl_B_0_port, Cin
                           => p4_ctrl_Cin, Als(31) => ctrl_LS_A_31_port, 
                           Als(30) => ctrl_LS_A_30_port, Als(29) => 
                           ctrl_LS_A_29_port, Als(28) => ctrl_LS_A_28_port, 
                           Als(27) => ctrl_LS_A_27_port, Als(26) => 
                           ctrl_LS_A_26_port, Als(25) => ctrl_LS_A_25_port, 
                           Als(24) => ctrl_LS_A_24_port, Als(23) => 
                           ctrl_LS_A_23_port, Als(22) => ctrl_LS_A_22_port, 
                           Als(21) => ctrl_LS_A_21_port, Als(20) => 
                           ctrl_LS_A_20_port, Als(19) => ctrl_LS_A_19_port, 
                           Als(18) => ctrl_LS_A_18_port, Als(17) => 
                           ctrl_LS_A_17_port, Als(16) => ctrl_LS_A_16_port, 
                           Als(15) => ctrl_LS_A_15_port, Als(14) => 
                           ctrl_LS_A_14_port, Als(13) => ctrl_LS_A_13_port, 
                           Als(12) => ctrl_LS_A_12_port, Als(11) => 
                           ctrl_LS_A_11_port, Als(10) => ctrl_LS_A_10_port, 
                           Als(9) => ctrl_LS_A_9_port, Als(8) => 
                           ctrl_LS_A_8_port, Als(7) => ctrl_LS_A_7_port, Als(6)
                           => ctrl_LS_A_6_port, Als(5) => ctrl_LS_A_5_port, 
                           Als(4) => ctrl_LS_A_4_port, Als(3) => 
                           ctrl_LS_A_3_port, Als(2) => ctrl_LS_A_2_port, Als(1)
                           => ctrl_LS_A_1_port, Als(0) => ctrl_LS_A_0_port, 
                           Bls(31) => ctrl_LS_B_31_port, Bls(30) => 
                           ctrl_LS_B_30_port, Bls(29) => ctrl_LS_B_29_port, 
                           Bls(28) => ctrl_LS_B_28_port, Bls(27) => 
                           ctrl_LS_B_27_port, Bls(26) => ctrl_LS_B_26_port, 
                           Bls(25) => ctrl_LS_B_25_port, Bls(24) => 
                           ctrl_LS_B_24_port, Bls(23) => ctrl_LS_B_23_port, 
                           Bls(22) => ctrl_LS_B_22_port, Bls(21) => 
                           ctrl_LS_B_21_port, Bls(20) => ctrl_LS_B_20_port, 
                           Bls(19) => ctrl_LS_B_19_port, Bls(18) => 
                           ctrl_LS_B_18_port, Bls(17) => ctrl_LS_B_17_port, 
                           Bls(16) => ctrl_LS_B_16_port, Bls(15) => 
                           ctrl_LS_B_15_port, Bls(14) => ctrl_LS_B_14_port, 
                           Bls(13) => ctrl_LS_B_13_port, Bls(12) => 
                           ctrl_LS_B_12_port, Bls(11) => ctrl_LS_B_11_port, 
                           Bls(10) => ctrl_LS_B_10_port, Bls(9) => 
                           ctrl_LS_B_9_port, Bls(8) => ctrl_LS_B_8_port, Bls(7)
                           => ctrl_LS_B_7_port, Bls(6) => ctrl_LS_B_6_port, 
                           Bls(5) => ctrl_LS_B_5_port, Bls(4) => 
                           ctrl_LS_B_4_port, Bls(3) => ctrl_LS_B_3_port, Bls(2)
                           => ctrl_LS_B_2_port, Bls(1) => ctrl_LS_B_1_port, 
                           Bls(0) => ctrl_LS_B_0_port, enableComp => 
                           enable_Comp);
   ADDER_SUB : P4_ADDER_NBITS32 port map( A(31) => p4_ctrl_A_31_port, A(30) => 
                           p4_ctrl_A_30_port, A(29) => p4_ctrl_A_29_port, A(28)
                           => p4_ctrl_A_28_port, A(27) => p4_ctrl_A_27_port, 
                           A(26) => p4_ctrl_A_26_port, A(25) => 
                           p4_ctrl_A_25_port, A(24) => p4_ctrl_A_24_port, A(23)
                           => p4_ctrl_A_23_port, A(22) => p4_ctrl_A_22_port, 
                           A(21) => p4_ctrl_A_21_port, A(20) => 
                           p4_ctrl_A_20_port, A(19) => p4_ctrl_A_19_port, A(18)
                           => p4_ctrl_A_18_port, A(17) => p4_ctrl_A_17_port, 
                           A(16) => p4_ctrl_A_16_port, A(15) => 
                           p4_ctrl_A_15_port, A(14) => p4_ctrl_A_14_port, A(13)
                           => p4_ctrl_A_13_port, A(12) => p4_ctrl_A_12_port, 
                           A(11) => p4_ctrl_A_11_port, A(10) => 
                           p4_ctrl_A_10_port, A(9) => p4_ctrl_A_9_port, A(8) =>
                           p4_ctrl_A_8_port, A(7) => p4_ctrl_A_7_port, A(6) => 
                           p4_ctrl_A_6_port, A(5) => p4_ctrl_A_5_port, A(4) => 
                           p4_ctrl_A_4_port, A(3) => p4_ctrl_A_3_port, A(2) => 
                           p4_ctrl_A_2_port, A(1) => p4_ctrl_A_1_port, A(0) => 
                           p4_ctrl_A_0_port, B(31) => p4_ctrl_B_31_port, B(30) 
                           => p4_ctrl_B_30_port, B(29) => p4_ctrl_B_29_port, 
                           B(28) => p4_ctrl_B_28_port, B(27) => 
                           p4_ctrl_B_27_port, B(26) => p4_ctrl_B_26_port, B(25)
                           => p4_ctrl_B_25_port, B(24) => p4_ctrl_B_24_port, 
                           B(23) => p4_ctrl_B_23_port, B(22) => 
                           p4_ctrl_B_22_port, B(21) => p4_ctrl_B_21_port, B(20)
                           => p4_ctrl_B_20_port, B(19) => p4_ctrl_B_19_port, 
                           B(18) => p4_ctrl_B_18_port, B(17) => 
                           p4_ctrl_B_17_port, B(16) => p4_ctrl_B_16_port, B(15)
                           => p4_ctrl_B_15_port, B(14) => p4_ctrl_B_14_port, 
                           B(13) => p4_ctrl_B_13_port, B(12) => 
                           p4_ctrl_B_12_port, B(11) => p4_ctrl_B_11_port, B(10)
                           => p4_ctrl_B_10_port, B(9) => p4_ctrl_B_9_port, B(8)
                           => p4_ctrl_B_8_port, B(7) => p4_ctrl_B_7_port, B(6) 
                           => p4_ctrl_B_6_port, B(5) => p4_ctrl_B_5_port, B(4) 
                           => p4_ctrl_B_4_port, B(3) => p4_ctrl_B_3_port, B(2) 
                           => p4_ctrl_B_2_port, B(1) => p4_ctrl_B_1_port, B(0) 
                           => p4_ctrl_B_0_port, Ci => p4_ctrl_Cin, S(31) => 
                           p4_outsig_31_port, S(30) => p4_outsig_30_port, S(29)
                           => p4_outsig_29_port, S(28) => p4_outsig_28_port, 
                           S(27) => p4_outsig_27_port, S(26) => 
                           p4_outsig_26_port, S(25) => p4_outsig_25_port, S(24)
                           => p4_outsig_24_port, S(23) => p4_outsig_23_port, 
                           S(22) => p4_outsig_22_port, S(21) => 
                           p4_outsig_21_port, S(20) => p4_outsig_20_port, S(19)
                           => p4_outsig_19_port, S(18) => p4_outsig_18_port, 
                           S(17) => p4_outsig_17_port, S(16) => 
                           p4_outsig_16_port, S(15) => p4_outsig_15_port, S(14)
                           => p4_outsig_14_port, S(13) => p4_outsig_13_port, 
                           S(12) => p4_outsig_12_port, S(11) => 
                           p4_outsig_11_port, S(10) => p4_outsig_10_port, S(9) 
                           => p4_outsig_9_port, S(8) => p4_outsig_8_port, S(7) 
                           => p4_outsig_7_port, S(6) => p4_outsig_6_port, S(5) 
                           => p4_outsig_5_port, S(4) => p4_outsig_4_port, S(3) 
                           => p4_outsig_3_port, S(2) => p4_outsig_2_port, S(1) 
                           => p4_outsig_1_port, S(0) => p4_outsig_0_port, Co =>
                           p4_comp_Co);
   LOGIC_SHIFT : logic_and_shift_N32 port map( FUNC(0) => FUNC(0), FUNC(1) => 
                           FUNC(1), FUNC(2) => FUNC(2), FUNC(3) => FUNC(3), 
                           DATA1(31) => ctrl_LS_A_31_port, DATA1(30) => 
                           ctrl_LS_A_30_port, DATA1(29) => ctrl_LS_A_29_port, 
                           DATA1(28) => ctrl_LS_A_28_port, DATA1(27) => 
                           ctrl_LS_A_27_port, DATA1(26) => ctrl_LS_A_26_port, 
                           DATA1(25) => ctrl_LS_A_25_port, DATA1(24) => 
                           ctrl_LS_A_24_port, DATA1(23) => ctrl_LS_A_23_port, 
                           DATA1(22) => ctrl_LS_A_22_port, DATA1(21) => 
                           ctrl_LS_A_21_port, DATA1(20) => ctrl_LS_A_20_port, 
                           DATA1(19) => ctrl_LS_A_19_port, DATA1(18) => 
                           ctrl_LS_A_18_port, DATA1(17) => ctrl_LS_A_17_port, 
                           DATA1(16) => ctrl_LS_A_16_port, DATA1(15) => 
                           ctrl_LS_A_15_port, DATA1(14) => ctrl_LS_A_14_port, 
                           DATA1(13) => ctrl_LS_A_13_port, DATA1(12) => 
                           ctrl_LS_A_12_port, DATA1(11) => ctrl_LS_A_11_port, 
                           DATA1(10) => ctrl_LS_A_10_port, DATA1(9) => 
                           ctrl_LS_A_9_port, DATA1(8) => ctrl_LS_A_8_port, 
                           DATA1(7) => ctrl_LS_A_7_port, DATA1(6) => 
                           ctrl_LS_A_6_port, DATA1(5) => ctrl_LS_A_5_port, 
                           DATA1(4) => ctrl_LS_A_4_port, DATA1(3) => 
                           ctrl_LS_A_3_port, DATA1(2) => ctrl_LS_A_2_port, 
                           DATA1(1) => ctrl_LS_A_1_port, DATA1(0) => 
                           ctrl_LS_A_0_port, DATA2(31) => ctrl_LS_B_31_port, 
                           DATA2(30) => ctrl_LS_B_30_port, DATA2(29) => 
                           ctrl_LS_B_29_port, DATA2(28) => ctrl_LS_B_28_port, 
                           DATA2(27) => ctrl_LS_B_27_port, DATA2(26) => 
                           ctrl_LS_B_26_port, DATA2(25) => ctrl_LS_B_25_port, 
                           DATA2(24) => ctrl_LS_B_24_port, DATA2(23) => 
                           ctrl_LS_B_23_port, DATA2(22) => ctrl_LS_B_22_port, 
                           DATA2(21) => ctrl_LS_B_21_port, DATA2(20) => 
                           ctrl_LS_B_20_port, DATA2(19) => ctrl_LS_B_19_port, 
                           DATA2(18) => ctrl_LS_B_18_port, DATA2(17) => 
                           ctrl_LS_B_17_port, DATA2(16) => ctrl_LS_B_16_port, 
                           DATA2(15) => ctrl_LS_B_15_port, DATA2(14) => 
                           ctrl_LS_B_14_port, DATA2(13) => ctrl_LS_B_13_port, 
                           DATA2(12) => ctrl_LS_B_12_port, DATA2(11) => 
                           ctrl_LS_B_11_port, DATA2(10) => ctrl_LS_B_10_port, 
                           DATA2(9) => ctrl_LS_B_9_port, DATA2(8) => 
                           ctrl_LS_B_8_port, DATA2(7) => ctrl_LS_B_7_port, 
                           DATA2(6) => ctrl_LS_B_6_port, DATA2(5) => 
                           ctrl_LS_B_5_port, DATA2(4) => ctrl_LS_B_4_port, 
                           DATA2(3) => ctrl_LS_B_3_port, DATA2(2) => 
                           ctrl_LS_B_2_port, DATA2(1) => ctrl_LS_B_1_port, 
                           DATA2(0) => ctrl_LS_B_0_port, OUTALU(31) => 
                           LS_OUTsig_31_port, OUTALU(30) => LS_OUTsig_30_port, 
                           OUTALU(29) => LS_OUTsig_29_port, OUTALU(28) => 
                           LS_OUTsig_28_port, OUTALU(27) => LS_OUTsig_27_port, 
                           OUTALU(26) => LS_OUTsig_26_port, OUTALU(25) => 
                           LS_OUTsig_25_port, OUTALU(24) => LS_OUTsig_24_port, 
                           OUTALU(23) => LS_OUTsig_23_port, OUTALU(22) => 
                           LS_OUTsig_22_port, OUTALU(21) => LS_OUTsig_21_port, 
                           OUTALU(20) => LS_OUTsig_20_port, OUTALU(19) => 
                           LS_OUTsig_19_port, OUTALU(18) => LS_OUTsig_18_port, 
                           OUTALU(17) => LS_OUTsig_17_port, OUTALU(16) => 
                           LS_OUTsig_16_port, OUTALU(15) => LS_OUTsig_15_port, 
                           OUTALU(14) => LS_OUTsig_14_port, OUTALU(13) => 
                           LS_OUTsig_13_port, OUTALU(12) => LS_OUTsig_12_port, 
                           OUTALU(11) => LS_OUTsig_11_port, OUTALU(10) => 
                           LS_OUTsig_10_port, OUTALU(9) => LS_OUTsig_9_port, 
                           OUTALU(8) => LS_OUTsig_8_port, OUTALU(7) => 
                           LS_OUTsig_7_port, OUTALU(6) => LS_OUTsig_6_port, 
                           OUTALU(5) => LS_OUTsig_5_port, OUTALU(4) => 
                           LS_OUTsig_4_port, OUTALU(3) => LS_OUTsig_3_port, 
                           OUTALU(2) => LS_OUTsig_2_port, OUTALU(1) => 
                           LS_OUTsig_1_port, OUTALU(0) => LS_OUTsig_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_0;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n33, n66, n67, n68, n69, n70 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n70, Z => n69);
   U2 : INV_X1 port map( A => S, ZN => n70);
   U3 : INV_X1 port map( A => n70, ZN => n68);
   U4 : BUF_X1 port map( A => n69, Z => n33);
   U5 : BUF_X1 port map( A => n69, Z => n67);
   U6 : BUF_X1 port map( A => n69, Z => n66);
   U7 : INV_X1 port map( A => n65, ZN => Y(0));
   U8 : AOI22_X1 port map( A1 => A(0), A2 => S, B1 => B(0), B2 => n33, ZN => 
                           n65);
   U9 : INV_X1 port map( A => n54, ZN => Y(1));
   U10 : AOI22_X1 port map( A1 => A(1), A2 => n68, B1 => B(1), B2 => n33, ZN =>
                           n54);
   U11 : INV_X1 port map( A => n40, ZN => Y(3));
   U12 : AOI22_X1 port map( A1 => A(3), A2 => n68, B1 => B(3), B2 => n67, ZN =>
                           n40);
   U13 : INV_X1 port map( A => n38, ZN => Y(5));
   U14 : AOI22_X1 port map( A1 => A(5), A2 => n68, B1 => B(5), B2 => n67, ZN =>
                           n38);
   U15 : INV_X1 port map( A => n43, ZN => Y(2));
   U16 : AOI22_X1 port map( A1 => A(2), A2 => n68, B1 => B(2), B2 => n66, ZN =>
                           n43);
   U17 : INV_X1 port map( A => n36, ZN => Y(7));
   U18 : AOI22_X1 port map( A1 => A(7), A2 => n68, B1 => B(7), B2 => n67, ZN =>
                           n36);
   U19 : INV_X1 port map( A => n34, ZN => Y(9));
   U20 : AOI22_X1 port map( A1 => n68, A2 => A(9), B1 => B(9), B2 => n67, ZN =>
                           n34);
   U21 : INV_X1 port map( A => n37, ZN => Y(6));
   U22 : AOI22_X1 port map( A1 => A(6), A2 => n68, B1 => B(6), B2 => n67, ZN =>
                           n37);
   U23 : INV_X1 port map( A => n61, ZN => Y(13));
   U24 : AOI22_X1 port map( A1 => A(13), A2 => S, B1 => B(13), B2 => n33, ZN =>
                           n61);
   U25 : INV_X1 port map( A => n63, ZN => Y(11));
   U26 : AOI22_X1 port map( A1 => A(11), A2 => S, B1 => B(11), B2 => n33, ZN =>
                           n63);
   U27 : INV_X1 port map( A => n59, ZN => Y(15));
   U28 : AOI22_X1 port map( A1 => A(15), A2 => S, B1 => B(15), B2 => n33, ZN =>
                           n59);
   U29 : INV_X1 port map( A => n39, ZN => Y(4));
   U30 : AOI22_X1 port map( A1 => A(4), A2 => n68, B1 => B(4), B2 => n67, ZN =>
                           n39);
   U31 : INV_X1 port map( A => n45, ZN => Y(28));
   U32 : AOI22_X1 port map( A1 => A(28), A2 => n68, B1 => B(28), B2 => n66, ZN 
                           => n45);
   U33 : INV_X1 port map( A => n64, ZN => Y(10));
   U34 : AOI22_X1 port map( A1 => A(10), A2 => S, B1 => B(10), B2 => n33, ZN =>
                           n64);
   U35 : INV_X1 port map( A => n57, ZN => Y(17));
   U36 : AOI22_X1 port map( A1 => A(17), A2 => S, B1 => B(17), B2 => n33, ZN =>
                           n57);
   U37 : INV_X1 port map( A => n58, ZN => Y(16));
   U38 : AOI22_X1 port map( A1 => A(16), A2 => S, B1 => B(16), B2 => n33, ZN =>
                           n58);
   U39 : INV_X1 port map( A => n62, ZN => Y(12));
   U40 : AOI22_X1 port map( A1 => A(12), A2 => S, B1 => B(12), B2 => n33, ZN =>
                           n62);
   U41 : INV_X1 port map( A => n60, ZN => Y(14));
   U42 : AOI22_X1 port map( A1 => A(14), A2 => S, B1 => B(14), B2 => n33, ZN =>
                           n60);
   U43 : INV_X1 port map( A => n52, ZN => Y(21));
   U44 : AOI22_X1 port map( A1 => A(21), A2 => n68, B1 => B(21), B2 => n66, ZN 
                           => n52);
   U45 : INV_X1 port map( A => n35, ZN => Y(8));
   U46 : AOI22_X1 port map( A1 => A(8), A2 => n68, B1 => B(8), B2 => n67, ZN =>
                           n35);
   U47 : INV_X1 port map( A => n55, ZN => Y(19));
   U48 : AOI22_X1 port map( A1 => A(19), A2 => S, B1 => B(19), B2 => n33, ZN =>
                           n55);
   U49 : INV_X1 port map( A => n53, ZN => Y(20));
   U50 : AOI22_X1 port map( A1 => A(20), A2 => n68, B1 => B(20), B2 => n66, ZN 
                           => n53);
   U51 : INV_X1 port map( A => n50, ZN => Y(23));
   U52 : AOI22_X1 port map( A1 => A(23), A2 => n68, B1 => B(23), B2 => n66, ZN 
                           => n50);
   U53 : INV_X1 port map( A => n49, ZN => Y(24));
   U54 : AOI22_X1 port map( A1 => A(24), A2 => n68, B1 => B(24), B2 => n66, ZN 
                           => n49);
   U55 : INV_X1 port map( A => n56, ZN => Y(18));
   U56 : AOI22_X1 port map( A1 => A(18), A2 => S, B1 => B(18), B2 => n33, ZN =>
                           n56);
   U57 : INV_X1 port map( A => n51, ZN => Y(22));
   U58 : AOI22_X1 port map( A1 => A(22), A2 => n68, B1 => B(22), B2 => n66, ZN 
                           => n51);
   U59 : INV_X1 port map( A => n44, ZN => Y(29));
   U60 : AOI22_X1 port map( A1 => A(29), A2 => n68, B1 => B(29), B2 => n66, ZN 
                           => n44);
   U61 : INV_X1 port map( A => n48, ZN => Y(25));
   U62 : AOI22_X1 port map( A1 => A(25), A2 => S, B1 => B(25), B2 => n66, ZN =>
                           n48);
   U63 : INV_X1 port map( A => n46, ZN => Y(27));
   U64 : AOI22_X1 port map( A1 => A(27), A2 => n68, B1 => B(27), B2 => n66, ZN 
                           => n46);
   U65 : INV_X1 port map( A => n47, ZN => Y(26));
   U66 : AOI22_X1 port map( A1 => A(26), A2 => n68, B1 => B(26), B2 => n66, ZN 
                           => n47);
   U67 : INV_X1 port map( A => n42, ZN => Y(30));
   U68 : AOI22_X1 port map( A1 => A(30), A2 => S, B1 => B(30), B2 => n66, ZN =>
                           n42);
   U69 : INV_X1 port map( A => n41, ZN => Y(31));
   U70 : AOI22_X1 port map( A1 => A(31), A2 => n68, B1 => B(31), B2 => n67, ZN 
                           => n41);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ZERO_DEC_bits32 is

   port( data : in std_logic_vector (31 downto 0);  zero_detect : out std_logic
         );

end ZERO_DEC_bits32;

architecture SYN_BEHAVIORAL of ZERO_DEC_bits32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1 : NOR4_X1 port map( A1 => data(23), A2 => data(22), A3 => data(21), A4 =>
                           data(20), ZN => n6);
   U2 : NAND4_X1 port map( A1 => n3, A2 => n4, A3 => n5, A4 => n6, ZN => n2);
   U3 : NOR4_X1 port map( A1 => data(12), A2 => data(11), A3 => data(10), A4 =>
                           data(0), ZN => n3);
   U4 : NOR4_X1 port map( A1 => data(16), A2 => data(15), A3 => data(14), A4 =>
                           data(13), ZN => n4);
   U5 : NOR4_X1 port map( A1 => data(1), A2 => data(19), A3 => data(18), A4 => 
                           data(17), ZN => n5);
   U6 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => zero_detect);
   U7 : NOR4_X1 port map( A1 => data(9), A2 => data(8), A3 => data(7), A4 => 
                           data(6), ZN => n10);
   U8 : NAND4_X1 port map( A1 => n7, A2 => n8, A3 => n9, A4 => n10, ZN => n1);
   U9 : NOR4_X1 port map( A1 => data(27), A2 => data(26), A3 => data(25), A4 =>
                           data(24), ZN => n7);
   U10 : NOR4_X1 port map( A1 => data(30), A2 => data(2), A3 => data(29), A4 =>
                           data(28), ZN => n8);
   U11 : NOR4_X1 port map( A1 => data(5), A2 => data(4), A3 => data(3), A4 => 
                           data(31), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity REGISTER_FILE_NBITS32_NREGISTERS32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end REGISTER_FILE_NBITS32_NREGISTERS32;

architecture SYN_BEHAVIORAL of REGISTER_FILE_NBITS32_NREGISTERS32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
      n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
      n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
      n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
      n2323, n2324, n2325, n2326, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, 
      n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, 
      n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, 
      n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
      n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, 
      n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, 
      n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, 
      n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
      n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, 
      n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, 
      n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, 
      n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, 
      n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, 
      n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, 
      n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
      n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, 
      n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
      n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
      n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, 
      n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, 
      n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, 
      n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, 
      n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, 
      n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
      n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, 
      n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, 
      n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, 
      n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
      n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
      n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, 
      n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, 
      n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
      n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, 
      n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, 
      n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
      n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
      n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, 
      n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, 
      n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, 
      n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, 
      n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, 
      n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, 
      n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, 
      n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
      n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, 
      n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, 
      n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, 
      n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, 
      n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, 
      n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, 
      n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, 
      n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, 
      n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, 
      n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, 
      n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, 
      n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, 
      n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, 
      n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, 
      n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, 
      n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, 
      n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, 
      n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, 
      n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, 
      n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, 
      n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, 
      n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, 
      n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, 
      n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, 
      n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, 
      n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, 
      n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, 
      n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, 
      n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, 
      n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, 
      n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, 
      n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, 
      n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, 
      n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, 
      n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, 
      n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, 
      n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, 
      n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, 
      n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, 
      n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, 
      n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, 
      n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, 
      n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, 
      n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, 
      n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, 
      n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, 
      n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, 
      n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, 
      n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, 
      n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, 
      n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, 
      n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, 
      n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, 
      n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, 
      n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, 
      n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, 
      n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, 
      n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, 
      n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, 
      n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, 
      n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, 
      n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, 
      n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, 
      n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, 
      n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, 
      n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, 
      n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, 
      n4157, n4158, n4159, n4160, n4161, n4162, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
      n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
      n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
      n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, 
      n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, 
      n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
      n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, 
      n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, 
      n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, 
      n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
      n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, 
      n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, 
      n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
      n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, 
      n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, 
      n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
      n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, 
      n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, 
      n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, 
      n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
      n1301, n1302, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, 
      n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, 
      n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, 
      n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, 
      n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, 
      n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, 
      n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, 
      n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, 
      n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, 
      n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, 
      n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, 
      n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, 
      n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, 
      n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, 
      n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, 
      n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, 
      n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
      n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, 
      n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, 
      n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, 
      n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, 
      n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
      n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, 
      n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, 
      n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, 
      n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, 
      n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, 
      n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, 
      n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, 
      n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, 
      n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, 
      n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, 
      n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, 
      n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, 
      n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, 
      n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, 
      n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, 
      n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, 
      n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, 
      n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, 
      n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, 
      n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, 
      n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, 
      n2755, n2756, n2757, n2758, n2759, n2760, n4163, n4164, n4165, n4166, 
      n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, 
      n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, 
      n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, 
      n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, 
      n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, 
      n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, 
      n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, 
      n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, 
      n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, 
      n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, 
      n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, 
      n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, 
      n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, 
      n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, 
      n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, 
      n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, 
      n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, 
      n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, 
      n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, 
      n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, 
      n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, 
      n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, 
      n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, 
      n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, 
      n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, 
      n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, 
      n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, 
      n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, 
      n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, 
      n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, 
      n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, 
      n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, 
      n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, 
      n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, 
      n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, 
      n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, 
      n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, 
      n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, 
      n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, 
      n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, 
      n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, 
      n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, 
      n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, 
      n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, 
      n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, 
      n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, 
      n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, 
      n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, 
      n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, 
      n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, 
      n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, 
      n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, 
      n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, 
      n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, 
      n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, 
      n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, 
      n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, 
      n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, 
      n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, 
      n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, 
      n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, 
      n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, 
      n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, 
      n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, 
      n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, 
      n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, 
      n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, 
      n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, 
      n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, 
      n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, 
      n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, 
      n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, 
      n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, 
      n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, 
      n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, 
      n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, 
      n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, 
      n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, 
      n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, 
      n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, 
      n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, 
      n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, 
      n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, 
      n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, 
      n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, 
      n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, 
      n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, 
      n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, 
      n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, 
      n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, 
      n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, 
      n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, 
      n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, 
      n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, 
      n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, 
      n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, 
      n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, 
      n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, 
      n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, 
      n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, 
      n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, 
      n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, 
      n5187, n5188, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, 
      n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, 
      n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, 
      n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, 
      n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, 
      n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, 
      n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, 
      n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, 
      n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, 
      n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, 
      n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, 
      n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, 
      n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, 
      n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, 
      n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, 
      n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, 
      n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, 
      n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, 
      n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, 
      n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, 
      n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, 
      n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, 
      n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, 
      n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, 
      n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, 
      n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, 
      n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, 
      n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, 
      n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, 
      n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, 
      n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, 
      n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, 
      n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, 
      n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, 
      n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, 
      n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, 
      n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, 
      n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, 
      n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, 
      n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, 
      n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, 
      n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, 
      n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, 
      n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, 
      n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, 
      n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, 
      n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, 
      n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, 
      n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, 
      n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, 
      n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, 
      n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, 
      n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, 
      n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, 
      n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, 
      n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, 
      n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, 
      n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, 
      n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, 
      n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, 
      n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, 
      n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, 
      n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, 
      n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, 
      n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, 
      n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, 
      n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, 
      n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, 
      n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, 
      n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, 
      n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, 
      n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, 
      n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, 
      n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, 
      n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, 
      n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, 
      n_1751, n_1752, n_1753, n_1754 : std_logic;

begin
   
   OUT2_reg_31_inst : DFF_X1 port map( D => n4130, CK => CLK, Q => OUT2(31), QN
                           => n3074);
   OUT2_reg_30_inst : DFF_X1 port map( D => n4129, CK => CLK, Q => OUT2(30), QN
                           => n3073);
   OUT2_reg_29_inst : DFF_X1 port map( D => n4128, CK => CLK, Q => OUT2(29), QN
                           => n3072);
   OUT2_reg_28_inst : DFF_X1 port map( D => n4127, CK => CLK, Q => OUT2(28), QN
                           => n3071);
   OUT2_reg_27_inst : DFF_X1 port map( D => n4126, CK => CLK, Q => OUT2(27), QN
                           => n3070);
   OUT2_reg_26_inst : DFF_X1 port map( D => n4125, CK => CLK, Q => OUT2(26), QN
                           => n3069);
   OUT2_reg_25_inst : DFF_X1 port map( D => n4124, CK => CLK, Q => OUT2(25), QN
                           => n3068);
   OUT2_reg_24_inst : DFF_X1 port map( D => n4123, CK => CLK, Q => OUT2(24), QN
                           => n3067);
   OUT2_reg_23_inst : DFF_X1 port map( D => n4122, CK => CLK, Q => OUT2(23), QN
                           => n3066);
   OUT2_reg_22_inst : DFF_X1 port map( D => n4121, CK => CLK, Q => OUT2(22), QN
                           => n3065);
   OUT2_reg_21_inst : DFF_X1 port map( D => n4120, CK => CLK, Q => OUT2(21), QN
                           => n3064);
   OUT2_reg_20_inst : DFF_X1 port map( D => n4119, CK => CLK, Q => OUT2(20), QN
                           => n3063);
   OUT2_reg_19_inst : DFF_X1 port map( D => n4118, CK => CLK, Q => OUT2(19), QN
                           => n3062);
   OUT2_reg_18_inst : DFF_X1 port map( D => n4117, CK => CLK, Q => OUT2(18), QN
                           => n3061);
   OUT2_reg_17_inst : DFF_X1 port map( D => n4116, CK => CLK, Q => OUT2(17), QN
                           => n3060);
   OUT2_reg_16_inst : DFF_X1 port map( D => n4115, CK => CLK, Q => OUT2(16), QN
                           => n3059);
   OUT2_reg_15_inst : DFF_X1 port map( D => n4114, CK => CLK, Q => OUT2(15), QN
                           => n3058);
   OUT2_reg_14_inst : DFF_X1 port map( D => n4113, CK => CLK, Q => OUT2(14), QN
                           => n3057);
   OUT2_reg_13_inst : DFF_X1 port map( D => n4112, CK => CLK, Q => OUT2(13), QN
                           => n3056);
   OUT2_reg_12_inst : DFF_X1 port map( D => n4111, CK => CLK, Q => OUT2(12), QN
                           => n3055);
   OUT2_reg_11_inst : DFF_X1 port map( D => n4110, CK => CLK, Q => OUT2(11), QN
                           => n3054);
   OUT2_reg_10_inst : DFF_X1 port map( D => n4109, CK => CLK, Q => OUT2(10), QN
                           => n3053);
   OUT2_reg_9_inst : DFF_X1 port map( D => n4108, CK => CLK, Q => OUT2(9), QN 
                           => n3052);
   OUT2_reg_8_inst : DFF_X1 port map( D => n4107, CK => CLK, Q => OUT2(8), QN 
                           => n3051);
   OUT2_reg_7_inst : DFF_X1 port map( D => n4106, CK => CLK, Q => OUT2(7), QN 
                           => n3050);
   OUT2_reg_6_inst : DFF_X1 port map( D => n4105, CK => CLK, Q => OUT2(6), QN 
                           => n3049);
   OUT2_reg_5_inst : DFF_X1 port map( D => n4104, CK => CLK, Q => OUT2(5), QN 
                           => n3048);
   OUT2_reg_4_inst : DFF_X1 port map( D => n4103, CK => CLK, Q => OUT2(4), QN 
                           => n3047);
   OUT2_reg_3_inst : DFF_X1 port map( D => n4102, CK => CLK, Q => OUT2(3), QN 
                           => n3046);
   OUT2_reg_2_inst : DFF_X1 port map( D => n4101, CK => CLK, Q => OUT2(2), QN 
                           => n3045);
   OUT2_reg_1_inst : DFF_X1 port map( D => n4100, CK => CLK, Q => OUT2(1), QN 
                           => n3044);
   OUT2_reg_0_inst : DFF_X1 port map( D => n4099, CK => CLK, Q => OUT2(0), QN 
                           => n3043);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2326, CK => CLK, Q => 
                           n_1051, QN => n4098);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2325, CK => CLK, Q => 
                           n_1052, QN => n4097);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2324, CK => CLK, Q => 
                           n_1053, QN => n4096);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2323, CK => CLK, Q => 
                           n_1054, QN => n4095);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2322, CK => CLK, Q => 
                           n_1055, QN => n4094);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2321, CK => CLK, Q => 
                           n_1056, QN => n4093);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2320, CK => CLK, Q => 
                           n_1057, QN => n4092);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2319, CK => CLK, Q => 
                           n_1058, QN => n4091);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2318, CK => CLK, Q => 
                           n_1059, QN => n4090);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2317, CK => CLK, Q => 
                           n_1060, QN => n4089);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2316, CK => CLK, Q => 
                           n_1061, QN => n4088);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2315, CK => CLK, Q => 
                           n_1062, QN => n4087);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2314, CK => CLK, Q => 
                           n_1063, QN => n4086);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2313, CK => CLK, Q => 
                           n_1064, QN => n4085);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2312, CK => CLK, Q => 
                           n_1065, QN => n4084);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2311, CK => CLK, Q => 
                           n_1066, QN => n4083);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2310, CK => CLK, Q => 
                           n_1067, QN => n4082);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2309, CK => CLK, Q => 
                           n_1068, QN => n4081);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2308, CK => CLK, Q => 
                           n_1069, QN => n4080);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2307, CK => CLK, Q => 
                           n_1070, QN => n4079);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2306, CK => CLK, Q => 
                           n_1071, QN => n4078);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2305, CK => CLK, Q => 
                           n_1072, QN => n4077);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2304, CK => CLK, Q => n_1073
                           , QN => n4076);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2303, CK => CLK, Q => n_1074
                           , QN => n4075);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2302, CK => CLK, Q => n_1075
                           , QN => n4074);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2301, CK => CLK, Q => n_1076
                           , QN => n4073);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2300, CK => CLK, Q => n_1077
                           , QN => n4072);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2299, CK => CLK, Q => n_1078
                           , QN => n4071);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2298, CK => CLK, Q => n_1079
                           , QN => n4070);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2297, CK => CLK, Q => n_1080
                           , QN => n4069);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2296, CK => CLK, Q => n_1081
                           , QN => n4068);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2295, CK => CLK, Q => n_1082
                           , QN => n4067);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2294, CK => CLK, Q => 
                           n_1083, QN => n4066);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2293, CK => CLK, Q => 
                           n_1084, QN => n4065);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2292, CK => CLK, Q => 
                           n_1085, QN => n4064);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2291, CK => CLK, Q => 
                           n_1086, QN => n4063);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2290, CK => CLK, Q => 
                           n_1087, QN => n4062);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2289, CK => CLK, Q => 
                           n_1088, QN => n4061);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2288, CK => CLK, Q => 
                           n_1089, QN => n4060);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2287, CK => CLK, Q => 
                           n_1090, QN => n4059);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2286, CK => CLK, Q => 
                           n_1091, QN => n4058);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2285, CK => CLK, Q => 
                           n_1092, QN => n4057);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2284, CK => CLK, Q => 
                           n_1093, QN => n4056);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2283, CK => CLK, Q => 
                           n_1094, QN => n4055);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2282, CK => CLK, Q => 
                           n_1095, QN => n4054);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2281, CK => CLK, Q => 
                           n_1096, QN => n4053);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2280, CK => CLK, Q => 
                           n_1097, QN => n4052);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2279, CK => CLK, Q => 
                           n_1098, QN => n4051);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2278, CK => CLK, Q => 
                           n_1099, QN => n4050);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2277, CK => CLK, Q => 
                           n_1100, QN => n4049);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2276, CK => CLK, Q => 
                           n_1101, QN => n4048);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2275, CK => CLK, Q => 
                           n_1102, QN => n4047);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2274, CK => CLK, Q => 
                           n_1103, QN => n4046);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2273, CK => CLK, Q => 
                           n_1104, QN => n4045);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2272, CK => CLK, Q => n_1105
                           , QN => n4044);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2271, CK => CLK, Q => n_1106
                           , QN => n4043);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2270, CK => CLK, Q => n_1107
                           , QN => n4042);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2269, CK => CLK, Q => n_1108
                           , QN => n4041);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2268, CK => CLK, Q => n_1109
                           , QN => n4040);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2267, CK => CLK, Q => n_1110
                           , QN => n4039);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2266, CK => CLK, Q => n_1111
                           , QN => n4038);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2265, CK => CLK, Q => n_1112
                           , QN => n4037);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2264, CK => CLK, Q => n_1113
                           , QN => n4036);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2263, CK => CLK, Q => n_1114
                           , QN => n4035);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2262, CK => CLK, Q => 
                           n_1115, QN => n4034);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2261, CK => CLK, Q => 
                           n_1116, QN => n4033);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2260, CK => CLK, Q => 
                           n_1117, QN => n4032);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2259, CK => CLK, Q => 
                           n_1118, QN => n4031);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2258, CK => CLK, Q => 
                           n_1119, QN => n4030);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2257, CK => CLK, Q => 
                           n_1120, QN => n4029);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2256, CK => CLK, Q => 
                           n_1121, QN => n4028);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2255, CK => CLK, Q => 
                           n_1122, QN => n4027);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2254, CK => CLK, Q => 
                           n_1123, QN => n4026);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2253, CK => CLK, Q => 
                           n_1124, QN => n4025);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2252, CK => CLK, Q => 
                           n_1125, QN => n4024);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2251, CK => CLK, Q => 
                           n_1126, QN => n4023);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2250, CK => CLK, Q => 
                           n_1127, QN => n4022);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2249, CK => CLK, Q => 
                           n_1128, QN => n4021);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2248, CK => CLK, Q => 
                           n_1129, QN => n4020);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2247, CK => CLK, Q => 
                           n_1130, QN => n4019);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2246, CK => CLK, Q => 
                           n_1131, QN => n4018);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2245, CK => CLK, Q => 
                           n_1132, QN => n4017);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2244, CK => CLK, Q => 
                           n_1133, QN => n4016);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2243, CK => CLK, Q => 
                           n_1134, QN => n4015);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2242, CK => CLK, Q => 
                           n_1135, QN => n4014);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2241, CK => CLK, Q => 
                           n_1136, QN => n4013);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2240, CK => CLK, Q => n_1137
                           , QN => n4012);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2239, CK => CLK, Q => n_1138
                           , QN => n4011);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2238, CK => CLK, Q => n_1139
                           , QN => n4010);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2237, CK => CLK, Q => n_1140
                           , QN => n4009);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2236, CK => CLK, Q => n_1141
                           , QN => n4008);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2235, CK => CLK, Q => n_1142
                           , QN => n4007);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2234, CK => CLK, Q => n_1143
                           , QN => n4006);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2233, CK => CLK, Q => n_1144
                           , QN => n4005);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2232, CK => CLK, Q => n_1145
                           , QN => n4004);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2231, CK => CLK, Q => n_1146
                           , QN => n4003);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2230, CK => CLK, Q => 
                           n_1147, QN => n4002);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2229, CK => CLK, Q => 
                           n_1148, QN => n4001);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2228, CK => CLK, Q => 
                           n_1149, QN => n4000);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2227, CK => CLK, Q => 
                           n_1150, QN => n3999);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2226, CK => CLK, Q => 
                           n_1151, QN => n3998);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2225, CK => CLK, Q => 
                           n_1152, QN => n3997);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2224, CK => CLK, Q => 
                           n_1153, QN => n3996);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2223, CK => CLK, Q => 
                           n_1154, QN => n3995);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2222, CK => CLK, Q => 
                           n_1155, QN => n3994);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2221, CK => CLK, Q => 
                           n_1156, QN => n3993);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2220, CK => CLK, Q => 
                           n_1157, QN => n3992);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2219, CK => CLK, Q => 
                           n_1158, QN => n3991);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2218, CK => CLK, Q => 
                           n_1159, QN => n3990);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2217, CK => CLK, Q => 
                           n_1160, QN => n3989);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2216, CK => CLK, Q => 
                           n_1161, QN => n3988);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2215, CK => CLK, Q => 
                           n_1162, QN => n3987);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2214, CK => CLK, Q => 
                           n_1163, QN => n3986);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2213, CK => CLK, Q => 
                           n_1164, QN => n3985);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2212, CK => CLK, Q => 
                           n_1165, QN => n3984);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2211, CK => CLK, Q => 
                           n_1166, QN => n3983);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2210, CK => CLK, Q => 
                           n_1167, QN => n3982);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2209, CK => CLK, Q => 
                           n_1168, QN => n3981);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2208, CK => CLK, Q => n_1169
                           , QN => n3980);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2207, CK => CLK, Q => n_1170
                           , QN => n3979);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2206, CK => CLK, Q => n_1171
                           , QN => n3978);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2205, CK => CLK, Q => n_1172
                           , QN => n3977);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2204, CK => CLK, Q => n_1173
                           , QN => n3976);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2203, CK => CLK, Q => n_1174
                           , QN => n3975);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2202, CK => CLK, Q => n_1175
                           , QN => n3974);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2201, CK => CLK, Q => n_1176
                           , QN => n3973);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2200, CK => CLK, Q => n_1177
                           , QN => n3972);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2199, CK => CLK, Q => n_1178
                           , QN => n3971);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2198, CK => CLK, Q => 
                           n_1179, QN => n3970);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2197, CK => CLK, Q => 
                           n_1180, QN => n3969);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2196, CK => CLK, Q => 
                           n_1181, QN => n3968);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2195, CK => CLK, Q => 
                           n_1182, QN => n3967);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2194, CK => CLK, Q => 
                           n_1183, QN => n3966);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2193, CK => CLK, Q => 
                           n_1184, QN => n3965);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2192, CK => CLK, Q => 
                           n_1185, QN => n3964);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2191, CK => CLK, Q => 
                           n_1186, QN => n3963);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2190, CK => CLK, Q => 
                           n_1187, QN => n3962);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2189, CK => CLK, Q => 
                           n_1188, QN => n3961);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2188, CK => CLK, Q => 
                           n_1189, QN => n3960);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2187, CK => CLK, Q => 
                           n_1190, QN => n3959);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2186, CK => CLK, Q => 
                           n_1191, QN => n3958);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2185, CK => CLK, Q => 
                           n_1192, QN => n3957);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2184, CK => CLK, Q => 
                           n_1193, QN => n3956);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2183, CK => CLK, Q => 
                           n_1194, QN => n3955);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2182, CK => CLK, Q => 
                           n_1195, QN => n3954);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2181, CK => CLK, Q => 
                           n_1196, QN => n3953);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2180, CK => CLK, Q => 
                           n_1197, QN => n3952);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2179, CK => CLK, Q => 
                           n_1198, QN => n3951);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2178, CK => CLK, Q => 
                           n_1199, QN => n3950);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2177, CK => CLK, Q => 
                           n_1200, QN => n3949);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2176, CK => CLK, Q => n_1201
                           , QN => n3948);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2175, CK => CLK, Q => n_1202
                           , QN => n3947);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2174, CK => CLK, Q => n_1203
                           , QN => n3946);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2173, CK => CLK, Q => n_1204
                           , QN => n3945);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2172, CK => CLK, Q => n_1205
                           , QN => n3944);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2171, CK => CLK, Q => n_1206
                           , QN => n3943);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2170, CK => CLK, Q => n_1207
                           , QN => n3942);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2169, CK => CLK, Q => n_1208
                           , QN => n3941);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2168, CK => CLK, Q => n_1209
                           , QN => n3940);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2167, CK => CLK, Q => n_1210
                           , QN => n3939);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           n_1211, QN => n3938);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           n_1212, QN => n3937);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           n_1213, QN => n3936);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           n_1214, QN => n3935);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           n_1215, QN => n3934);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           n_1216, QN => n3933);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           n_1217, QN => n3932);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           n_1218, QN => n3931);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           n_1219, QN => n3930);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           n_1220, QN => n3929);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           n_1221, QN => n3928);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           n_1222, QN => n3927);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           n_1223, QN => n3926);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => 
                           n_1224, QN => n3925);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => 
                           n_1225, QN => n3924);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => 
                           n_1226, QN => n3923);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => 
                           n_1227, QN => n3922);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => 
                           n_1228, QN => n3921);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => 
                           n_1229, QN => n3920);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => 
                           n_1230, QN => n3919);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => 
                           n_1231, QN => n3918);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => 
                           n_1232, QN => n3917);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => n_1233
                           , QN => n3916);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => n_1234
                           , QN => n3915);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => n_1235
                           , QN => n3914);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => n_1236
                           , QN => n3913);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => n_1237
                           , QN => n3912);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => n_1238
                           , QN => n3911);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => n_1239
                           , QN => n3910);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => n_1240
                           , QN => n3909);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => n_1241
                           , QN => n3908);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => n_1242
                           , QN => n3907);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => 
                           n_1243, QN => n3906);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => 
                           n_1244, QN => n3905);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => 
                           n_1245, QN => n3904);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => 
                           n_1246, QN => n3903);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => 
                           n_1247, QN => n3902);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => 
                           n_1248, QN => n3901);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => 
                           n_1249, QN => n3900);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => 
                           n_1250, QN => n3899);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           n_1251, QN => n3898);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           n_1252, QN => n3897);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           n_1253, QN => n3896);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           n_1254, QN => n3895);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           n_1255, QN => n3894);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => 
                           n_1256, QN => n3893);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => 
                           n_1257, QN => n3892);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => 
                           n_1258, QN => n3891);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => 
                           n_1259, QN => n3890);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => 
                           n_1260, QN => n3889);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => 
                           n_1261, QN => n3888);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => 
                           n_1262, QN => n3887);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => 
                           n_1263, QN => n3886);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => 
                           n_1264, QN => n3885);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => n_1265
                           , QN => n3884);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => n_1266
                           , QN => n3883);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => n_1267
                           , QN => n3882);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => n_1268
                           , QN => n3881);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => n_1269
                           , QN => n3880);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => n_1270
                           , QN => n3879);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => n_1271
                           , QN => n3878);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => n_1272
                           , QN => n3877);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => n_1273
                           , QN => n3876);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => n_1274
                           , QN => n3875);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           n_1275, QN => n3874);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           n_1276, QN => n3873);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           n_1277, QN => n3872);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           n_1278, QN => n3871);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           n_1279, QN => n3870);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           n_1280, QN => n3869);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           n_1281, QN => n3868);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           n_1282, QN => n3867);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           n_1283, QN => n3866);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           n_1284, QN => n3865);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           n_1285, QN => n3864);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           n_1286, QN => n3863);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           n_1287, QN => n3862);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => 
                           n_1288, QN => n3861);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           n_1289, QN => n3860);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => 
                           n_1290, QN => n3859);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => 
                           n_1291, QN => n3858);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => 
                           n_1292, QN => n3857);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => 
                           n_1293, QN => n3856);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => 
                           n_1294, QN => n3855);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => 
                           n_1295, QN => n3854);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => 
                           n_1296, QN => n3853);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => n_1297
                           , QN => n3852);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => n_1298
                           , QN => n3851);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => n_1299
                           , QN => n3850);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => n_1300
                           , QN => n3849);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => n_1301
                           , QN => n3848);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => n_1302
                           , QN => n3847);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => n_1303
                           , QN => n3846);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => n_1304
                           , QN => n3845);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => n_1305
                           , QN => n3844);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => n_1306
                           , QN => n3843);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           n_1307, QN => n3842);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           n_1308, QN => n3841);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           n_1309, QN => n3840);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           n_1310, QN => n3839);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           n_1311, QN => n3838);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           n_1312, QN => n3837);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           n_1313, QN => n3836);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           n_1314, QN => n3835);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           n_1315, QN => n3834);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           n_1316, QN => n3833);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           n_1317, QN => n3832);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           n_1318, QN => n3831);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           n_1319, QN => n3830);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           n_1320, QN => n3829);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           n_1321, QN => n3828);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => 
                           n_1322, QN => n3827);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => 
                           n_1323, QN => n3826);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => 
                           n_1324, QN => n3825);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => 
                           n_1325, QN => n3824);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => 
                           n_1326, QN => n3823);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => 
                           n_1327, QN => n3822);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => 
                           n_1328, QN => n3821);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => n_1329
                           , QN => n3820);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => n_1330
                           , QN => n3819);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => n_1331
                           , QN => n3818);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => n_1332
                           , QN => n3817);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => n_1333
                           , QN => n3816);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => n_1334
                           , QN => n3815);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => n_1335
                           , QN => n3814);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => n_1336
                           , QN => n3813);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => n_1337
                           , QN => n3812);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => n_1338
                           , QN => n3811);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           n_1339, QN => n3810);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           n_1340, QN => n3809);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           n_1341, QN => n3808);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           n_1342, QN => n3807);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           n_1343, QN => n3806);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           n_1344, QN => n3805);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           n_1345, QN => n3804);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           n_1346, QN => n3803);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           n_1347, QN => n3802);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           n_1348, QN => n3801);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           n_1349, QN => n3800);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           n_1350, QN => n3799);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           n_1351, QN => n3798);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => 
                           n_1352, QN => n3797);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => 
                           n_1353, QN => n3796);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => 
                           n_1354, QN => n3795);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => 
                           n_1355, QN => n3794);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => 
                           n_1356, QN => n3793);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => 
                           n_1357, QN => n3792);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => 
                           n_1358, QN => n3791);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => 
                           n_1359, QN => n3790);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => 
                           n_1360, QN => n3789);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => n_1361
                           , QN => n3788);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => n_1362
                           , QN => n3787);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => n_1363
                           , QN => n3786);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => n_1364
                           , QN => n3785);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => n_1365
                           , QN => n3784);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => n_1366
                           , QN => n3783);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => n_1367
                           , QN => n3782);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => n_1368
                           , QN => n3781);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => n_1369
                           , QN => n3780);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => n_1370
                           , QN => n3779);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           n_1371, QN => n3778);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           n_1372, QN => n3777);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           n_1373, QN => n3776);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           n_1374, QN => n3775);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           n_1375, QN => n3774);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           n_1376, QN => n3773);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           n_1377, QN => n3772);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           n_1378, QN => n3771);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           n_1379, QN => n3770);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           n_1380, QN => n3769);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           n_1381, QN => n3768);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           n_1382, QN => n3767);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           n_1383, QN => n3766);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           n_1384, QN => n3765);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           n_1385, QN => n3764);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           n_1386, QN => n3763);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           n_1387, QN => n3762);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           n_1388, QN => n3761);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           n_1389, QN => n3760);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           n_1390, QN => n3759);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           n_1391, QN => n3758);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           n_1392, QN => n3757);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           n_1393, QN => n3756);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           n_1394, QN => n3755);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           n_1395, QN => n3754);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           n_1396, QN => n3753);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           n_1397, QN => n3752);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           n_1398, QN => n3751);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           n_1399, QN => n3750);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           n_1400, QN => n3749);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           n_1401, QN => n3748);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           n_1402, QN => n3747);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           n_1403, QN => n3746);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           n_1404, QN => n3745);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           n_1405, QN => n3744);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           n_1406, QN => n3743);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           n_1407, QN => n3742);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           n_1408, QN => n3741);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           n_1409, QN => n3740);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           n_1410, QN => n3739);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           n_1411, QN => n3738);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           n_1412, QN => n3737);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           n_1413, QN => n3736);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           n_1414, QN => n3735);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           n_1415, QN => n3734);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           n_1416, QN => n3733);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           n_1417, QN => n3732);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           n_1418, QN => n3731);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           n_1419, QN => n3730);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           n_1420, QN => n3729);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           n_1421, QN => n3728);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           n_1422, QN => n3727);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           n_1423, QN => n3726);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => 
                           n_1424, QN => n3725);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => 
                           n_1425, QN => n3724);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           n_1426, QN => n3723);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           n_1427, QN => n3722);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           n_1428, QN => n3721);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           n_1429, QN => n3720);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           n_1430, QN => n3719);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           n_1431, QN => n3718);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           n_1432, QN => n3717);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           n_1433, QN => n3716);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           n_1434, QN => n3715);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           n_1435, QN => n3714);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           n_1436, QN => n3713);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           n_1437, QN => n3712);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           n_1438, QN => n3711);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           n_1439, QN => n3710);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           n_1440, QN => n3709);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           n_1441, QN => n3708);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           n_1442, QN => n3707);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           n_1443, QN => n3706);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           n_1444, QN => n3705);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           n_1445, QN => n3704);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           n_1446, QN => n3703);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           n_1447, QN => n3702);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           n_1448, QN => n3701);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           n_1449, QN => n3700);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           n_1450, QN => n3699);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           n_1451, QN => n3698);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           n_1452, QN => n3697);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           n_1453, QN => n3696);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           n_1454, QN => n3695);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           n_1455, QN => n3694);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => 
                           n_1456, QN => n3693);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => 
                           n_1457, QN => n3692);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           n_1458, QN => n3691);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           n_1459, QN => n3690);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           n_1460, QN => n3689);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           n_1461, QN => n3688);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           n_1462, QN => n3687);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           n_1463, QN => n3686);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           n_1464, QN => n3685);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           n_1465, QN => n3684);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           n_1466, QN => n3683);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           n_1467, QN => n3682);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           n_1468, QN => n3681);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           n_1469, QN => n3680);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           n_1470, QN => n3679);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           n_1471, QN => n3678);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           n_1472, QN => n3677);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           n_1473, QN => n3676);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           n_1474, QN => n3675);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           n_1475, QN => n3674);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           n_1476, QN => n3673);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           n_1477, QN => n3672);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           n_1478, QN => n3671);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           n_1479, QN => n3670);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           n_1480, QN => n3669);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           n_1481, QN => n3668);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           n_1482, QN => n3667);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           n_1483, QN => n3666);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           n_1484, QN => n3665);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           n_1485, QN => n3664);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           n_1486, QN => n3663);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           n_1487, QN => n3662);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           n_1488, QN => n3661);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           n_1489, QN => n3660);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           n_1490, QN => n3659);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           n_1491, QN => n3658);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           n_1492, QN => n3657);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           n_1493, QN => n3656);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           n_1494, QN => n3655);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           n_1495, QN => n3654);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           n_1496, QN => n3653);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           n_1497, QN => n3652);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           n_1498, QN => n3651);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           n_1499, QN => n3650);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           n_1500, QN => n3649);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           n_1501, QN => n3648);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           n_1502, QN => n3647);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           n_1503, QN => n3646);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           n_1504, QN => n3645);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           n_1505, QN => n3644);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           n_1506, QN => n3643);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           n_1507, QN => n3642);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           n_1508, QN => n3641);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           n_1509, QN => n3640);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           n_1510, QN => n3639);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           n_1511, QN => n3638);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           n_1512, QN => n3637);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           n_1513, QN => n3636);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           n_1514, QN => n3635);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           n_1515, QN => n3634);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           n_1516, QN => n3633);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           n_1517, QN => n3632);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           n_1518, QN => n3631);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           n_1519, QN => n3630);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           n_1520, QN => n3629);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           n_1521, QN => n3628);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           n_1522, QN => n3627);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           n_1523, QN => n3626);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           n_1524, QN => n3625);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           n_1525, QN => n3624);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           n_1526, QN => n3623);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           n_1527, QN => n3622);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           n_1528, QN => n3621);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           n_1529, QN => n3620);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           n_1530, QN => n3619);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           n_1531, QN => n3618);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           n_1532, QN => n3617);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           n_1533, QN => n3616);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           n_1534, QN => n3615);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           n_1535, QN => n3614);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           n_1536, QN => n3613);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           n_1537, QN => n3612);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           n_1538, QN => n3611);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           n_1539, QN => n3610);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           n_1540, QN => n3609);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           n_1541, QN => n3608);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           n_1542, QN => n3607);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           n_1543, QN => n3606);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           n_1544, QN => n3605);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           n_1545, QN => n3604);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           n_1546, QN => n3603);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           n_1547, QN => n3602);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           n_1548, QN => n3601);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           n_1549, QN => n3600);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           n_1550, QN => n3599);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           n_1551, QN => n3598);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => 
                           n_1552, QN => n3597);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => 
                           n_1553, QN => n3596);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           n_1554, QN => n3595);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           n_1555, QN => n3594);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           n_1556, QN => n3593);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           n_1557, QN => n3592);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           n_1558, QN => n3591);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           n_1559, QN => n3590);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           n_1560, QN => n3589);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           n_1561, QN => n3588);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           n_1562, QN => n3587);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           n4258, QN => n3586);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           n4257, QN => n3585);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           n4256, QN => n3584);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           n4255, QN => n3583);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           n4254, QN => n3582);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           n4253, QN => n3581);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           n4252, QN => n3580);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           n4251, QN => n3579);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           n4250, QN => n3578);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           n4249, QN => n3577);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           n4248, QN => n3576);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           n4247, QN => n3575);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           n4246, QN => n3574);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           n4245, QN => n3573);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           n4244, QN => n3572);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           n4243, QN => n3571);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           n4242, QN => n3570);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           n4241, QN => n3569);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           n4240, QN => n3568);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           n4239, QN => n3567);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           n4238, QN => n3566);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           n4237, QN => n3565);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => n4236
                           , QN => n3564);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => n4235
                           , QN => n3563);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => n4234
                           , QN => n3562);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => n4233
                           , QN => n3561);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => n4232
                           , QN => n3560);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => n4231
                           , QN => n3559);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => n4230
                           , QN => n3558);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => n4229
                           , QN => n3557);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => n4228
                           , QN => n3556);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => n4227
                           , QN => n3555);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           n_1563, QN => n3554);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           n_1564, QN => n3553);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           n_1565, QN => n3552);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           n_1566, QN => n3551);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           n_1567, QN => n3550);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           n_1568, QN => n3549);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           n_1569, QN => n3548);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           n_1570, QN => n3547);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           n_1571, QN => n3546);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           n_1572, QN => n3545);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           n_1573, QN => n3544);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           n_1574, QN => n3543);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           n_1575, QN => n3542);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           n_1576, QN => n3541);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           n_1577, QN => n3540);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           n_1578, QN => n3539);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           n_1579, QN => n3538);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           n_1580, QN => n3537);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           n_1581, QN => n3536);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           n_1582, QN => n3535);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           n_1583, QN => n3534);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           n_1584, QN => n3533);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           n_1585, QN => n3532);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           n_1586, QN => n3531);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           n_1587, QN => n3530);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           n_1588, QN => n3529);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           n_1589, QN => n3528);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           n_1590, QN => n3527);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           n_1591, QN => n3526);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           n_1592, QN => n3525);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           n_1593, QN => n3524);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           n_1594, QN => n3523);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           n4354, QN => n3522);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           n4353, QN => n3521);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           n4352, QN => n3520);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           n4351, QN => n3519);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           n4350, QN => n3518);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           n4349, QN => n3517);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           n4348, QN => n3516);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           n4347, QN => n3515);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           n4346, QN => n3514);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           n4345, QN => n3513);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           n4344, QN => n3512);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           n4343, QN => n3511);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           n4342, QN => n3510);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           n4341, QN => n3509);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           n4340, QN => n3508);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           n4339, QN => n3507);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           n4338, QN => n3506);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           n4337, QN => n3505);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           n4336, QN => n3504);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           n4335, QN => n3503);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           n4334, QN => n3502);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           n4333, QN => n3501);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => n4332
                           , QN => n3500);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => n4331
                           , QN => n3499);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => n4330
                           , QN => n3498);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => n4329
                           , QN => n3497);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => n4328
                           , QN => n3496);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => n4327
                           , QN => n3495);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => n4326
                           , QN => n3494);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => n4325
                           , QN => n3493);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => n4324
                           , QN => n3492);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => n4323
                           , QN => n3491);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           n_1595, QN => n3490);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           n_1596, QN => n3489);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           n_1597, QN => n3488);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           n_1598, QN => n3487);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           n_1599, QN => n3486);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           n_1600, QN => n3485);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           n_1601, QN => n3484);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           n_1602, QN => n3483);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           n_1603, QN => n3482);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           n_1604, QN => n3481);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           n_1605, QN => n3480);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           n_1606, QN => n3479);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           n_1607, QN => n3478);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           n_1608, QN => n3477);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           n_1609, QN => n3476);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           n_1610, QN => n3475);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           n_1611, QN => n3474);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           n_1612, QN => n3473);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           n_1613, QN => n3472);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           n_1614, QN => n3471);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           n_1615, QN => n3470);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           n_1616, QN => n3469);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           n_1617, QN => n3468);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           n_1618, QN => n3467);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           n_1619, QN => n3466);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           n_1620, QN => n3465);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           n_1621, QN => n3464);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           n_1622, QN => n3463);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           n_1623, QN => n3462);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           n_1624, QN => n3461);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           n_1625, QN => n3460);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           n_1626, QN => n3459);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           n4386, QN => n3458);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           n4385, QN => n3457);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           n4384, QN => n3456);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           n4383, QN => n3455);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           n4382, QN => n3454);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           n4381, QN => n3453);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           n4380, QN => n3452);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           n4379, QN => n3451);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           n4378, QN => n3450);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           n4377, QN => n3449);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           n4376, QN => n3448);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           n4375, QN => n3447);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           n4374, QN => n3446);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           n4373, QN => n3445);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           n4372, QN => n3444);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           n4371, QN => n3443);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           n4370, QN => n3442);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           n4369, QN => n3441);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           n4368, QN => n3440);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           n4367, QN => n3439);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           n4366, QN => n3438);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           n4365, QN => n3437);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => n4364
                           , QN => n3436);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => n4363
                           , QN => n3435);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => n4362
                           , QN => n3434);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => n4361
                           , QN => n3433);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => n4360
                           , QN => n3432);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => n4359
                           , QN => n3431);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => n4358
                           , QN => n3430);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => n4357
                           , QN => n3429);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => n4356
                           , QN => n3428);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => n4355
                           , QN => n3427);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           n4322, QN => n3426);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           n4321, QN => n3425);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           n4320, QN => n3424);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           n4319, QN => n3423);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           n4318, QN => n3422);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           n4317, QN => n3421);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           n4316, QN => n3420);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           n4315, QN => n3419);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           n4314, QN => n3418);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           n4313, QN => n3417);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           n4312, QN => n3416);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           n4311, QN => n3415);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           n4310, QN => n3414);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           n4309, QN => n3413);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           n4308, QN => n3412);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           n4307, QN => n3411);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           n4306, QN => n3410);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           n4305, QN => n3409);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           n4304, QN => n3408);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           n4303, QN => n3407);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           n4302, QN => n3406);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           n4301, QN => n3405);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => n4300
                           , QN => n3404);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => n4299
                           , QN => n3403);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => n4298
                           , QN => n3402);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => n4297
                           , QN => n3401);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n4296
                           , QN => n3400);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => n4295
                           , QN => n3399);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n4294
                           , QN => n3398);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => n4293
                           , QN => n3397);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n4292
                           , QN => n3396);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => n4291
                           , QN => n3395);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           n4194, QN => n3394);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           n4193, QN => n3393);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           n4192, QN => n3392);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           n4191, QN => n3391);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           n4190, QN => n3390);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           n4189, QN => n3389);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           n4188, QN => n3388);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           n4187, QN => n3387);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           n4186, QN => n3386);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           n4185, QN => n3385);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           n4184, QN => n3384);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           n4183, QN => n3383);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           n4182, QN => n3382);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           n4181, QN => n3381);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           n4180, QN => n3380);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           n4179, QN => n3379);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           n4178, QN => n3378);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           n4177, QN => n3377);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           n4176, QN => n3376);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           n4175, QN => n3375);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           n4174, QN => n3374);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           n4173, QN => n3373);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n4172
                           , QN => n3372);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => n4171
                           , QN => n3371);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n4170
                           , QN => n3370);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => n4169
                           , QN => n3369);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n4168
                           , QN => n3368);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => n4167
                           , QN => n3367);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n4166
                           , QN => n3366);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => n4165
                           , QN => n3365);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n4164
                           , QN => n3364);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => n4163
                           , QN => n3363);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           n4418, QN => n3362);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           n4417, QN => n3361);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           n4416, QN => n3360);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           n4415, QN => n3359);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           n4414, QN => n3358);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           n4413, QN => n3357);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           n4412, QN => n3356);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           n4411, QN => n3355);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           n4410, QN => n3354);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           n4409, QN => n3353);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           n4408, QN => n3352);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           n4407, QN => n3351);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           n4406, QN => n3350);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           n4405, QN => n3349);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           n4404, QN => n3348);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           n4403, QN => n3347);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           n4402, QN => n3346);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           n4401, QN => n3345);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           n4400, QN => n3344);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           n4399, QN => n3343);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           n4398, QN => n3342);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           n4397, QN => n3341);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n4396
                           , QN => n3340);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => n4395
                           , QN => n3339);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n4394
                           , QN => n3338);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => n4393
                           , QN => n3337);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n4392
                           , QN => n3336);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => n4391
                           , QN => n3335);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n4390
                           , QN => n3334);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => n4389
                           , QN => n3333);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n4388
                           , QN => n3332);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => n4387
                           , QN => n3331);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           n4226, QN => n3330);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           n4225, QN => n3329);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           n4224, QN => n3328);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           n4223, QN => n3327);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           n4222, QN => n3326);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           n4221, QN => n3325);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           n4220, QN => n3324);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           n4219, QN => n3323);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           n4218, QN => n3322);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           n4217, QN => n3321);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           n4216, QN => n3320);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           n4215, QN => n3319);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           n4214, QN => n3318);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           n4213, QN => n3317);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           n4212, QN => n3316);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           n4211, QN => n3315);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           n4210, QN => n3314);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           n4209, QN => n3313);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           n4208, QN => n3312);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           n4207, QN => n3311);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           n4206, QN => n3310);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           n4205, QN => n3309);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n4204
                           , QN => n3308);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => n4203
                           , QN => n3307);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n4202
                           , QN => n3306);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => n4201
                           , QN => n3305);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n4200
                           , QN => n3304);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => n4199
                           , QN => n3303);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n4198
                           , QN => n3302);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => n4197
                           , QN => n3301);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n4196
                           , QN => n3300);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => n4195
                           , QN => n3299);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           n_1627, QN => n3298);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           n_1628, QN => n3297);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           n_1629, QN => n3296);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           n_1630, QN => n3295);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           n_1631, QN => n3294);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           n_1632, QN => n3293);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           n_1633, QN => n3292);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           n_1634, QN => n3291);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           n_1635, QN => n3290);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           n_1636, QN => n3289);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           n_1637, QN => n3288);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           n_1638, QN => n3287);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           n_1639, QN => n3286);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           n_1640, QN => n3285);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           n_1641, QN => n3284);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           n_1642, QN => n3283);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           n_1643, QN => n3282);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           n_1644, QN => n3281);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           n_1645, QN => n3280);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           n_1646, QN => n3279);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           n_1647, QN => n3278);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           n_1648, QN => n3277);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           n_1649, QN => n3276);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           n_1650, QN => n3275);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           n_1651, QN => n3274);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           n_1652, QN => n3273);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           n_1653, QN => n3272);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           n_1654, QN => n3271);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           n_1655, QN => n3270);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           n_1656, QN => n3269);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           n_1657, QN => n3268);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           n_1658, QN => n3267);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           n4290, QN => n3266);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           n4289, QN => n3265);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           n4288, QN => n3264);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           n4287, QN => n3263);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           n4286, QN => n3262);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           n4285, QN => n3261);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           n4284, QN => n3260);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           n4283, QN => n3259);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           n4282, QN => n3258);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           n4281, QN => n3257);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           n4280, QN => n3256);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           n4279, QN => n3255);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           n4278, QN => n3254);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           n4277, QN => n3253);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           n4276, QN => n3252);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           n4275, QN => n3251);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           n4274, QN => n3250);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           n4273, QN => n3249);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           n4272, QN => n3248);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           n4271, QN => n3247);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           n4270, QN => n3246);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           n4269, QN => n3245);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n4268
                           , QN => n3244);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => n4267
                           , QN => n3243);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => n4266
                           , QN => n3242);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => n4265
                           , QN => n3241);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => n4264
                           , QN => n3240);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => n4263
                           , QN => n3239);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => n4262
                           , QN => n3238);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => n4261
                           , QN => n3237);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => n4260
                           , QN => n3236);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => n4259
                           , QN => n3235);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           n_1659, QN => n3234);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           n_1660, QN => n3233);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           n_1661, QN => n3232);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           n_1662, QN => n3231);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           n_1663, QN => n3230);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           n_1664, QN => n3229);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           n_1665, QN => n3228);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           n_1666, QN => n3227);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           n_1667, QN => n3226);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           n_1668, QN => n3225);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           n_1669, QN => n3224);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           n_1670, QN => n3223);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           n_1671, QN => n3222);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           n_1672, QN => n3221);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           n_1673, QN => n3220);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           n_1674, QN => n3219);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           n_1675, QN => n3218);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           n_1676, QN => n3217);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           n_1677, QN => n3216);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           n_1678, QN => n3215);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           n_1679, QN => n3214);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           n_1680, QN => n3213);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           n_1681, QN => n3212);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           n_1682, QN => n3211);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           n_1683, QN => n3210);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           n_1684, QN => n3209);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           n_1685, QN => n3208);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           n_1686, QN => n3207);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           n_1687, QN => n3206);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           n_1688, QN => n3205);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           n_1689, QN => n3204);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           n_1690, QN => n3203);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           n_1691, QN => n3202);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           n_1692, QN => n3201);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           n_1693, QN => n3200);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           n_1694, QN => n3199);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           n_1695, QN => n3198);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           n_1696, QN => n3197);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           n_1697, QN => n3196);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           n_1698, QN => n3195);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           n_1699, QN => n3194);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           n_1700, QN => n3193);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           n_1701, QN => n3192);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           n_1702, QN => n3191);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           n_1703, QN => n3190);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           n_1704, QN => n3189);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           n_1705, QN => n3188);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           n_1706, QN => n3187);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           n_1707, QN => n3186);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           n_1708, QN => n3185);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           n_1709, QN => n3184);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           n_1710, QN => n3183);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           n_1711, QN => n3182);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           n_1712, QN => n3181);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           n_1713, QN => n3180);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           n_1714, QN => n3179);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           n_1715, QN => n3178);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           n_1716, QN => n3177);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           n_1717, QN => n3176);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           n_1718, QN => n3175);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           n_1719, QN => n3174);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           n_1720, QN => n3173);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           n_1721, QN => n3172);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           n_1722, QN => n3171);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           n4482, QN => n3170);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           n4481, QN => n3169);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           n4480, QN => n3168);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           n4479, QN => n3167);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           n4478, QN => n3166);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           n4477, QN => n3165);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           n4476, QN => n3164);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           n4475, QN => n3163);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           n4474, QN => n3162);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           n4473, QN => n3161);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           n4472, QN => n3160);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           n4471, QN => n3159);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           n4470, QN => n3158);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           n4469, QN => n3157);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           n4468, QN => n3156);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           n4467, QN => n3155);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           n4466, QN => n3154);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           n4465, QN => n3153);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           n4464, QN => n3152);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           n4463, QN => n3151);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           n4462, QN => n3150);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => 
                           n4461, QN => n3149);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => n4460
                           , QN => n3148);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => n4459
                           , QN => n3147);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => n4458
                           , QN => n3146);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => n4457
                           , QN => n3145);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => n4456
                           , QN => n3144);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => n4455
                           , QN => n3143);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => n4454
                           , QN => n3142);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => n4453
                           , QN => n3141);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => n4452
                           , QN => n3140);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => n4451
                           , QN => n3139);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           n4450, QN => n3138);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           n4449, QN => n3137);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           n4448, QN => n3136);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           n4447, QN => n3135);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           n4446, QN => n3134);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           n4445, QN => n3133);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           n4444, QN => n3132);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           n4443, QN => n3131);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           n4442, QN => n3130);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           n4441, QN => n3129);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           n4440, QN => n3128);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           n4439, QN => n3127);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           n4438, QN => n3126);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           n4437, QN => n3125);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           n4436, QN => n3124);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           n4435, QN => n3123);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           n4434, QN => n3122);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           n4433, QN => n3121);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           n4432, QN => n3120);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           n4431, QN => n3119);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           n4430, QN => n3118);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => 
                           n4429, QN => n3117);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => n4428
                           , QN => n3116);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => n4427
                           , QN => n3115);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => n4426
                           , QN => n3114);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => n4425
                           , QN => n3113);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => n4424
                           , QN => n3112);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => n4423
                           , QN => n3111);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => n4422
                           , QN => n3110);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => n4421
                           , QN => n3109);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => n4420
                           , QN => n3108);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => n4419
                           , QN => n3107);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => 
                           n_1723, QN => n3106);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => 
                           n_1724, QN => n3105);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => 
                           n_1725, QN => n3104);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => 
                           n_1726, QN => n3103);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => 
                           n_1727, QN => n3102);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => 
                           n_1728, QN => n3101);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => 
                           n_1729, QN => n3100);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => 
                           n_1730, QN => n3099);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => 
                           n_1731, QN => n3098);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => 
                           n_1732, QN => n3097);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => 
                           n_1733, QN => n3096);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => 
                           n_1734, QN => n3095);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => 
                           n_1735, QN => n3094);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => 
                           n_1736, QN => n3093);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => 
                           n_1737, QN => n3092);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => 
                           n_1738, QN => n3091);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => 
                           n_1739, QN => n3090);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => 
                           n_1740, QN => n3089);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => 
                           n_1741, QN => n3088);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => 
                           n_1742, QN => n3087);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => 
                           n_1743, QN => n3086);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => 
                           n_1744, QN => n3085);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => 
                           n_1745, QN => n3084);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => 
                           n_1746, QN => n3083);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => 
                           n_1747, QN => n3082);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => 
                           n_1748, QN => n3081);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => 
                           n_1749, QN => n3080);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => 
                           n_1750, QN => n3079);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => 
                           n_1751, QN => n3078);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => 
                           n_1752, QN => n3077);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => 
                           n_1753, QN => n3076);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => 
                           n_1754, QN => n3075);
   OUT1_reg_31_inst : DFF_X1 port map( D => n4162, CK => CLK, Q => OUT1(31), QN
                           => n3042);
   OUT1_reg_30_inst : DFF_X1 port map( D => n4161, CK => CLK, Q => OUT1(30), QN
                           => n3041);
   OUT1_reg_29_inst : DFF_X1 port map( D => n4160, CK => CLK, Q => OUT1(29), QN
                           => n3040);
   OUT1_reg_28_inst : DFF_X1 port map( D => n4159, CK => CLK, Q => OUT1(28), QN
                           => n3039);
   OUT1_reg_27_inst : DFF_X1 port map( D => n4158, CK => CLK, Q => OUT1(27), QN
                           => n3038);
   OUT1_reg_26_inst : DFF_X1 port map( D => n4157, CK => CLK, Q => OUT1(26), QN
                           => n3037);
   OUT1_reg_25_inst : DFF_X1 port map( D => n4156, CK => CLK, Q => OUT1(25), QN
                           => n3036);
   OUT1_reg_24_inst : DFF_X1 port map( D => n4155, CK => CLK, Q => OUT1(24), QN
                           => n3035);
   OUT1_reg_23_inst : DFF_X1 port map( D => n4154, CK => CLK, Q => OUT1(23), QN
                           => n3034);
   OUT1_reg_22_inst : DFF_X1 port map( D => n4153, CK => CLK, Q => OUT1(22), QN
                           => n3033);
   OUT1_reg_21_inst : DFF_X1 port map( D => n4152, CK => CLK, Q => OUT1(21), QN
                           => n3032);
   OUT1_reg_20_inst : DFF_X1 port map( D => n4151, CK => CLK, Q => OUT1(20), QN
                           => n3031);
   OUT1_reg_19_inst : DFF_X1 port map( D => n4150, CK => CLK, Q => OUT1(19), QN
                           => n3030);
   OUT1_reg_18_inst : DFF_X1 port map( D => n4149, CK => CLK, Q => OUT1(18), QN
                           => n3029);
   OUT1_reg_17_inst : DFF_X1 port map( D => n4148, CK => CLK, Q => OUT1(17), QN
                           => n3028);
   OUT1_reg_16_inst : DFF_X1 port map( D => n4147, CK => CLK, Q => OUT1(16), QN
                           => n3027);
   OUT1_reg_15_inst : DFF_X1 port map( D => n4146, CK => CLK, Q => OUT1(15), QN
                           => n3026);
   OUT1_reg_14_inst : DFF_X1 port map( D => n4145, CK => CLK, Q => OUT1(14), QN
                           => n3025);
   OUT1_reg_13_inst : DFF_X1 port map( D => n4144, CK => CLK, Q => OUT1(13), QN
                           => n3024);
   OUT1_reg_12_inst : DFF_X1 port map( D => n4143, CK => CLK, Q => OUT1(12), QN
                           => n3023);
   OUT1_reg_11_inst : DFF_X1 port map( D => n4142, CK => CLK, Q => OUT1(11), QN
                           => n3022);
   OUT1_reg_10_inst : DFF_X1 port map( D => n4141, CK => CLK, Q => OUT1(10), QN
                           => n3021);
   OUT1_reg_9_inst : DFF_X1 port map( D => n4140, CK => CLK, Q => OUT1(9), QN 
                           => n3020);
   OUT1_reg_8_inst : DFF_X1 port map( D => n4139, CK => CLK, Q => OUT1(8), QN 
                           => n3019);
   OUT1_reg_7_inst : DFF_X1 port map( D => n4138, CK => CLK, Q => OUT1(7), QN 
                           => n3018);
   OUT1_reg_6_inst : DFF_X1 port map( D => n4137, CK => CLK, Q => OUT1(6), QN 
                           => n3017);
   OUT1_reg_5_inst : DFF_X1 port map( D => n4136, CK => CLK, Q => OUT1(5), QN 
                           => n3016);
   OUT1_reg_4_inst : DFF_X1 port map( D => n4135, CK => CLK, Q => OUT1(4), QN 
                           => n3015);
   OUT1_reg_3_inst : DFF_X1 port map( D => n4134, CK => CLK, Q => OUT1(3), QN 
                           => n3014);
   OUT1_reg_2_inst : DFF_X1 port map( D => n4133, CK => CLK, Q => OUT1(2), QN 
                           => n3013);
   OUT1_reg_1_inst : DFF_X1 port map( D => n4132, CK => CLK, Q => OUT1(1), QN 
                           => n3012);
   OUT1_reg_0_inst : DFF_X1 port map( D => n4131, CK => CLK, Q => OUT1(0), QN 
                           => n3011);
   U3 : BUF_X1 port map( A => n2685, Z => n4955);
   U4 : BUF_X1 port map( A => n2695, Z => n4931);
   U5 : BUF_X1 port map( A => n2692, Z => n4939);
   U6 : BUF_X1 port map( A => n2689, Z => n4947);
   U7 : BUF_X1 port map( A => n2748, Z => n4755);
   U8 : BUF_X1 port map( A => n2745, Z => n4763);
   U9 : BUF_X1 port map( A => n2735, Z => n4803);
   U10 : BUF_X1 port map( A => n2733, Z => n4811);
   U11 : BUF_X1 port map( A => n2731, Z => n4819);
   U12 : BUF_X1 port map( A => n2728, Z => n4827);
   U13 : BUF_X1 port map( A => n2718, Z => n4867);
   U14 : BUF_X1 port map( A => n2716, Z => n4875);
   U15 : BUF_X1 port map( A => n2714, Z => n4883);
   U16 : BUF_X1 port map( A => n2711, Z => n4891);
   U17 : BUF_X1 port map( A => n2752, Z => n4739);
   U18 : BUF_X1 port map( A => n2750, Z => n4747);
   U19 : BUF_X1 port map( A => n2707, Z => n4899);
   U20 : BUF_X1 port map( A => n2704, Z => n4907);
   U21 : BUF_X1 port map( A => n2701, Z => n4915);
   U22 : BUF_X1 port map( A => n2698, Z => n4923);
   U23 : BUF_X1 port map( A => n2726, Z => n4835);
   U24 : BUF_X1 port map( A => n2724, Z => n4843);
   U25 : BUF_X1 port map( A => n2722, Z => n4851);
   U26 : BUF_X1 port map( A => n2720, Z => n4859);
   U27 : BUF_X1 port map( A => n2743, Z => n4771);
   U28 : BUF_X1 port map( A => n2741, Z => n4779);
   U29 : BUF_X1 port map( A => n2739, Z => n4787);
   U30 : BUF_X1 port map( A => n2737, Z => n4795);
   U31 : BUF_X1 port map( A => n2758, Z => n4715);
   U32 : BUF_X1 port map( A => n2756, Z => n4723);
   U33 : BUF_X1 port map( A => n2754, Z => n4731);
   U34 : BUF_X1 port map( A => n2760, Z => n4707);
   U35 : BUF_X1 port map( A => n5128, Z => n4498);
   U36 : BUF_X1 port map( A => n5128, Z => n4497);
   U37 : BUF_X1 port map( A => n5141, Z => n4562);
   U38 : BUF_X1 port map( A => n5141, Z => n4561);
   U39 : BUF_X1 port map( A => n2684, Z => n4959);
   U40 : BUF_X1 port map( A => n2694, Z => n4935);
   U41 : BUF_X1 port map( A => n2691, Z => n4943);
   U42 : BUF_X1 port map( A => n2688, Z => n4951);
   U43 : BUF_X1 port map( A => n2747, Z => n4759);
   U44 : BUF_X1 port map( A => n2744, Z => n4767);
   U45 : BUF_X1 port map( A => n2734, Z => n4807);
   U46 : BUF_X1 port map( A => n2732, Z => n4815);
   U47 : BUF_X1 port map( A => n2730, Z => n4823);
   U48 : BUF_X1 port map( A => n2727, Z => n4831);
   U49 : BUF_X1 port map( A => n2717, Z => n4871);
   U50 : BUF_X1 port map( A => n2715, Z => n4879);
   U51 : BUF_X1 port map( A => n2713, Z => n4887);
   U52 : BUF_X1 port map( A => n2710, Z => n4895);
   U53 : BUF_X1 port map( A => n2751, Z => n4743);
   U54 : BUF_X1 port map( A => n2749, Z => n4751);
   U55 : BUF_X1 port map( A => n2706, Z => n4903);
   U56 : BUF_X1 port map( A => n2703, Z => n4911);
   U57 : BUF_X1 port map( A => n2700, Z => n4919);
   U58 : BUF_X1 port map( A => n2697, Z => n4927);
   U59 : BUF_X1 port map( A => n2725, Z => n4839);
   U60 : BUF_X1 port map( A => n2723, Z => n4847);
   U61 : BUF_X1 port map( A => n2721, Z => n4855);
   U62 : BUF_X1 port map( A => n2719, Z => n4863);
   U63 : BUF_X1 port map( A => n2742, Z => n4775);
   U64 : BUF_X1 port map( A => n2740, Z => n4783);
   U65 : BUF_X1 port map( A => n2738, Z => n4791);
   U66 : BUF_X1 port map( A => n2736, Z => n4799);
   U67 : BUF_X1 port map( A => n2757, Z => n4719);
   U68 : BUF_X1 port map( A => n2755, Z => n4727);
   U69 : BUF_X1 port map( A => n2753, Z => n4735);
   U70 : BUF_X1 port map( A => n2759, Z => n4711);
   U71 : BUF_X1 port map( A => n5140, Z => n4554);
   U72 : BUF_X1 port map( A => n5143, Z => n4578);
   U73 : BUF_X1 port map( A => n5140, Z => n4553);
   U74 : BUF_X1 port map( A => n5127, Z => n4490);
   U75 : BUF_X1 port map( A => n5127, Z => n4489);
   U76 : BUF_X1 port map( A => n5143, Z => n4577);
   U77 : BUF_X1 port map( A => n5130, Z => n4514);
   U78 : BUF_X1 port map( A => n5130, Z => n4513);
   U79 : BUF_X1 port map( A => n5142, Z => n4570);
   U80 : BUF_X1 port map( A => n5142, Z => n4569);
   U81 : BUF_X1 port map( A => n5129, Z => n4506);
   U82 : BUF_X1 port map( A => n5129, Z => n4505);
   U83 : BUF_X1 port map( A => n5133, Z => n4530);
   U84 : BUF_X1 port map( A => n5133, Z => n4529);
   U85 : BUF_X1 port map( A => n5146, Z => n4594);
   U86 : BUF_X1 port map( A => n5146, Z => n4593);
   U87 : BUF_X1 port map( A => n5132, Z => n4522);
   U88 : BUF_X1 port map( A => n5132, Z => n4521);
   U89 : BUF_X1 port map( A => n5145, Z => n4586);
   U90 : BUF_X1 port map( A => n5145, Z => n4585);
   U91 : BUF_X1 port map( A => n5147, Z => n4602);
   U92 : BUF_X1 port map( A => n5147, Z => n4601);
   U93 : BUF_X1 port map( A => n5134, Z => n4538);
   U94 : BUF_X1 port map( A => n5134, Z => n4537);
   U95 : BUF_X1 port map( A => n5148, Z => n4610);
   U96 : BUF_X1 port map( A => n5148, Z => n4609);
   U97 : BUF_X1 port map( A => n5135, Z => n4546);
   U98 : BUF_X1 port map( A => n5135, Z => n4545);
   U99 : BUF_X1 port map( A => n413, Z => n5071);
   U100 : BUF_X1 port map( A => n1051, Z => n4991);
   U101 : BUF_X1 port map( A => n384, Z => n5119);
   U102 : BUF_X1 port map( A => n1022, Z => n5039);
   U103 : BUF_X1 port map( A => n1049, Z => n5002);
   U104 : BUF_X1 port map( A => n411, Z => n5082);
   U105 : BUF_X1 port map( A => n410, Z => n5086);
   U106 : BUF_X1 port map( A => n1048, Z => n5006);
   U107 : BUF_X1 port map( A => n1060, Z => n4966);
   U108 : BUF_X1 port map( A => n422, Z => n5046);
   U109 : BUF_X1 port map( A => n1059, Z => n4970);
   U110 : BUF_X1 port map( A => n421, Z => n5050);
   U111 : BUF_X1 port map( A => n1047, Z => n5007);
   U112 : BUF_X1 port map( A => n397, Z => n5102);
   U113 : BUF_X1 port map( A => n396, Z => n5103);
   U114 : BUF_X1 port map( A => n409, Z => n5087);
   U115 : BUF_X1 port map( A => n1035, Z => n5022);
   U116 : BUF_X1 port map( A => n1034, Z => n5023);
   U117 : BUF_X1 port map( A => n1054, Z => n4986);
   U118 : BUF_X1 port map( A => n416, Z => n5066);
   U119 : BUF_X1 port map( A => n1058, Z => n4971);
   U120 : BUF_X1 port map( A => n420, Z => n5051);
   U121 : BUF_X1 port map( A => n1053, Z => n4987);
   U122 : BUF_X1 port map( A => n415, Z => n5067);
   U123 : BUF_X1 port map( A => n406, Z => n5095);
   U124 : BUF_X1 port map( A => n1044, Z => n5015);
   U125 : BUF_X1 port map( A => n412, Z => n5075);
   U126 : BUF_X1 port map( A => n1050, Z => n4995);
   U127 : BUF_X1 port map( A => n1055, Z => n4979);
   U128 : BUF_X1 port map( A => n417, Z => n5059);
   U129 : BUF_X1 port map( A => n407, Z => n5091);
   U130 : BUF_X1 port map( A => n1045, Z => n5011);
   U131 : BUF_X1 port map( A => n418, Z => n5055);
   U132 : BUF_X1 port map( A => n1056, Z => n4975);
   U133 : BUF_X1 port map( A => n1032, Z => n5027);
   U134 : BUF_X1 port map( A => n394, Z => n5107);
   U135 : BUF_X1 port map( A => n392, Z => n5111);
   U136 : BUF_X1 port map( A => n1030, Z => n5031);
   U137 : BUF_X1 port map( A => n386, Z => n5115);
   U138 : BUF_X1 port map( A => n1024, Z => n5035);
   U139 : BUF_X1 port map( A => n4955, Z => n4958);
   U140 : BUF_X1 port map( A => n4955, Z => n4956);
   U141 : BUF_X1 port map( A => n4955, Z => n4957);
   U142 : BUF_X1 port map( A => n4931, Z => n4934);
   U143 : BUF_X1 port map( A => n4939, Z => n4942);
   U144 : BUF_X1 port map( A => n4947, Z => n4950);
   U145 : BUF_X1 port map( A => n4931, Z => n4932);
   U146 : BUF_X1 port map( A => n4931, Z => n4933);
   U147 : BUF_X1 port map( A => n4939, Z => n4940);
   U148 : BUF_X1 port map( A => n4939, Z => n4941);
   U149 : BUF_X1 port map( A => n4947, Z => n4948);
   U150 : BUF_X1 port map( A => n4947, Z => n4949);
   U151 : BUF_X1 port map( A => n4755, Z => n4758);
   U152 : BUF_X1 port map( A => n4803, Z => n4806);
   U153 : BUF_X1 port map( A => n4867, Z => n4870);
   U154 : BUF_X1 port map( A => n4875, Z => n4878);
   U155 : BUF_X1 port map( A => n4883, Z => n4886);
   U156 : BUF_X1 port map( A => n4891, Z => n4894);
   U157 : BUF_X1 port map( A => n4739, Z => n4742);
   U158 : BUF_X1 port map( A => n4747, Z => n4750);
   U159 : BUF_X1 port map( A => n4763, Z => n4766);
   U160 : BUF_X1 port map( A => n4811, Z => n4814);
   U161 : BUF_X1 port map( A => n4819, Z => n4822);
   U162 : BUF_X1 port map( A => n4827, Z => n4830);
   U163 : BUF_X1 port map( A => n4755, Z => n4756);
   U164 : BUF_X1 port map( A => n4755, Z => n4757);
   U165 : BUF_X1 port map( A => n4803, Z => n4804);
   U166 : BUF_X1 port map( A => n4803, Z => n4805);
   U167 : BUF_X1 port map( A => n4739, Z => n4740);
   U168 : BUF_X1 port map( A => n4739, Z => n4741);
   U169 : BUF_X1 port map( A => n4747, Z => n4748);
   U170 : BUF_X1 port map( A => n4747, Z => n4749);
   U171 : BUF_X1 port map( A => n4763, Z => n4764);
   U172 : BUF_X1 port map( A => n4763, Z => n4765);
   U173 : BUF_X1 port map( A => n4811, Z => n4812);
   U174 : BUF_X1 port map( A => n4811, Z => n4813);
   U175 : BUF_X1 port map( A => n4819, Z => n4820);
   U176 : BUF_X1 port map( A => n4819, Z => n4821);
   U177 : BUF_X1 port map( A => n4827, Z => n4828);
   U178 : BUF_X1 port map( A => n4827, Z => n4829);
   U179 : BUF_X1 port map( A => n4867, Z => n4868);
   U180 : BUF_X1 port map( A => n4867, Z => n4869);
   U181 : BUF_X1 port map( A => n4875, Z => n4876);
   U182 : BUF_X1 port map( A => n4875, Z => n4877);
   U183 : BUF_X1 port map( A => n4883, Z => n4884);
   U184 : BUF_X1 port map( A => n4883, Z => n4885);
   U185 : BUF_X1 port map( A => n4891, Z => n4892);
   U186 : BUF_X1 port map( A => n4891, Z => n4893);
   U187 : BUF_X1 port map( A => n4899, Z => n4902);
   U188 : BUF_X1 port map( A => n4907, Z => n4910);
   U189 : BUF_X1 port map( A => n4915, Z => n4918);
   U190 : BUF_X1 port map( A => n4923, Z => n4926);
   U191 : BUF_X1 port map( A => n4899, Z => n4900);
   U192 : BUF_X1 port map( A => n4899, Z => n4901);
   U193 : BUF_X1 port map( A => n4907, Z => n4908);
   U194 : BUF_X1 port map( A => n4907, Z => n4909);
   U195 : BUF_X1 port map( A => n4915, Z => n4916);
   U196 : BUF_X1 port map( A => n4915, Z => n4917);
   U197 : BUF_X1 port map( A => n4923, Z => n4924);
   U198 : BUF_X1 port map( A => n4923, Z => n4925);
   U199 : BUF_X1 port map( A => n4835, Z => n4838);
   U200 : BUF_X1 port map( A => n4843, Z => n4846);
   U201 : BUF_X1 port map( A => n4851, Z => n4854);
   U202 : BUF_X1 port map( A => n4859, Z => n4862);
   U203 : BUF_X1 port map( A => n4771, Z => n4774);
   U204 : BUF_X1 port map( A => n4779, Z => n4782);
   U205 : BUF_X1 port map( A => n4787, Z => n4790);
   U206 : BUF_X1 port map( A => n4795, Z => n4798);
   U207 : BUF_X1 port map( A => n4835, Z => n4836);
   U208 : BUF_X1 port map( A => n4835, Z => n4837);
   U209 : BUF_X1 port map( A => n4843, Z => n4844);
   U210 : BUF_X1 port map( A => n4843, Z => n4845);
   U211 : BUF_X1 port map( A => n4851, Z => n4852);
   U212 : BUF_X1 port map( A => n4851, Z => n4853);
   U213 : BUF_X1 port map( A => n4859, Z => n4860);
   U214 : BUF_X1 port map( A => n4859, Z => n4861);
   U215 : BUF_X1 port map( A => n4771, Z => n4772);
   U216 : BUF_X1 port map( A => n4771, Z => n4773);
   U217 : BUF_X1 port map( A => n4779, Z => n4780);
   U218 : BUF_X1 port map( A => n4779, Z => n4781);
   U219 : BUF_X1 port map( A => n4787, Z => n4788);
   U220 : BUF_X1 port map( A => n4787, Z => n4789);
   U221 : BUF_X1 port map( A => n4795, Z => n4796);
   U222 : BUF_X1 port map( A => n4795, Z => n4797);
   U223 : BUF_X1 port map( A => n4715, Z => n4718);
   U224 : BUF_X1 port map( A => n4731, Z => n4734);
   U225 : BUF_X1 port map( A => n4723, Z => n4726);
   U226 : BUF_X1 port map( A => n4715, Z => n4716);
   U227 : BUF_X1 port map( A => n4715, Z => n4717);
   U228 : BUF_X1 port map( A => n4731, Z => n4732);
   U229 : BUF_X1 port map( A => n4731, Z => n4733);
   U230 : BUF_X1 port map( A => n4723, Z => n4724);
   U231 : BUF_X1 port map( A => n4723, Z => n4725);
   U232 : BUF_X1 port map( A => n4707, Z => n4710);
   U233 : BUF_X1 port map( A => n4707, Z => n4708);
   U234 : BUF_X1 port map( A => n4707, Z => n4709);
   U235 : NAND2_X1 port map( A1 => n5125, A2 => n4960, ZN => n2685);
   U236 : NAND2_X1 port map( A1 => n5125, A2 => n4936, ZN => n2695);
   U237 : NAND2_X1 port map( A1 => n5125, A2 => n4944, ZN => n2692);
   U238 : NAND2_X1 port map( A1 => n5125, A2 => n4952, ZN => n2689);
   U239 : NAND2_X1 port map( A1 => n5123, A2 => n4760, ZN => n2748);
   U240 : NAND2_X1 port map( A1 => n5124, A2 => n4808, ZN => n2735);
   U241 : NAND2_X1 port map( A1 => n5124, A2 => n4872, ZN => n2718);
   U242 : NAND2_X1 port map( A1 => n5124, A2 => n4880, ZN => n2716);
   U243 : NAND2_X1 port map( A1 => n5124, A2 => n4888, ZN => n2714);
   U244 : NAND2_X1 port map( A1 => n5124, A2 => n4896, ZN => n2711);
   U245 : NAND2_X1 port map( A1 => n5123, A2 => n4744, ZN => n2752);
   U246 : NAND2_X1 port map( A1 => n5123, A2 => n4752, ZN => n2750);
   U247 : NAND2_X1 port map( A1 => n5123, A2 => n4768, ZN => n2745);
   U248 : NAND2_X1 port map( A1 => n5124, A2 => n4816, ZN => n2733);
   U249 : NAND2_X1 port map( A1 => n5124, A2 => n4824, ZN => n2731);
   U250 : NAND2_X1 port map( A1 => n5124, A2 => n4832, ZN => n2728);
   U251 : NAND2_X1 port map( A1 => n5125, A2 => n4904, ZN => n2707);
   U252 : NAND2_X1 port map( A1 => n5125, A2 => n4912, ZN => n2704);
   U253 : NAND2_X1 port map( A1 => n5125, A2 => n4920, ZN => n2701);
   U254 : NAND2_X1 port map( A1 => n5125, A2 => n4928, ZN => n2698);
   U255 : NAND2_X1 port map( A1 => n5124, A2 => n4840, ZN => n2726);
   U256 : NAND2_X1 port map( A1 => n5124, A2 => n4848, ZN => n2724);
   U257 : NAND2_X1 port map( A1 => n5124, A2 => n4856, ZN => n2722);
   U258 : NAND2_X1 port map( A1 => n5124, A2 => n4864, ZN => n2720);
   U259 : NAND2_X1 port map( A1 => n5123, A2 => n4776, ZN => n2743);
   U260 : NAND2_X1 port map( A1 => n5123, A2 => n4784, ZN => n2741);
   U261 : NAND2_X1 port map( A1 => n5123, A2 => n4792, ZN => n2739);
   U262 : NAND2_X1 port map( A1 => n5123, A2 => n4800, ZN => n2737);
   U263 : NAND2_X1 port map( A1 => n5123, A2 => n4720, ZN => n2758);
   U264 : NAND2_X1 port map( A1 => n5123, A2 => n4736, ZN => n2754);
   U265 : NAND2_X1 port map( A1 => n5123, A2 => n4728, ZN => n2756);
   U266 : NAND2_X1 port map( A1 => n5123, A2 => n4712, ZN => n2760);
   U267 : BUF_X1 port map( A => n4562, Z => n4555);
   U268 : BUF_X1 port map( A => n4562, Z => n4556);
   U269 : BUF_X1 port map( A => n4562, Z => n4557);
   U270 : BUF_X1 port map( A => n4561, Z => n4558);
   U271 : BUF_X1 port map( A => n4561, Z => n4559);
   U272 : BUF_X1 port map( A => n4498, Z => n4491);
   U273 : BUF_X1 port map( A => n4498, Z => n4492);
   U274 : BUF_X1 port map( A => n4498, Z => n4493);
   U275 : BUF_X1 port map( A => n4497, Z => n4494);
   U276 : BUF_X1 port map( A => n4497, Z => n4495);
   U277 : BUF_X1 port map( A => n4561, Z => n4560);
   U278 : BUF_X1 port map( A => n4497, Z => n4496);
   U279 : BUF_X1 port map( A => n4959, Z => n4960);
   U280 : BUF_X1 port map( A => n4935, Z => n4936);
   U281 : BUF_X1 port map( A => n4943, Z => n4944);
   U282 : BUF_X1 port map( A => n4951, Z => n4952);
   U283 : BUF_X1 port map( A => n4759, Z => n4760);
   U284 : BUF_X1 port map( A => n4807, Z => n4808);
   U285 : BUF_X1 port map( A => n4871, Z => n4872);
   U286 : BUF_X1 port map( A => n4879, Z => n4880);
   U287 : BUF_X1 port map( A => n4887, Z => n4888);
   U288 : BUF_X1 port map( A => n4895, Z => n4896);
   U289 : BUF_X1 port map( A => n4743, Z => n4744);
   U290 : BUF_X1 port map( A => n4751, Z => n4752);
   U291 : BUF_X1 port map( A => n4767, Z => n4768);
   U292 : BUF_X1 port map( A => n4815, Z => n4816);
   U293 : BUF_X1 port map( A => n4823, Z => n4824);
   U294 : BUF_X1 port map( A => n4831, Z => n4832);
   U295 : BUF_X1 port map( A => n4903, Z => n4904);
   U296 : BUF_X1 port map( A => n4911, Z => n4912);
   U297 : BUF_X1 port map( A => n4919, Z => n4920);
   U298 : BUF_X1 port map( A => n4927, Z => n4928);
   U299 : BUF_X1 port map( A => n4839, Z => n4840);
   U300 : BUF_X1 port map( A => n4847, Z => n4848);
   U301 : BUF_X1 port map( A => n4855, Z => n4856);
   U302 : BUF_X1 port map( A => n4863, Z => n4864);
   U303 : BUF_X1 port map( A => n4775, Z => n4776);
   U304 : BUF_X1 port map( A => n4783, Z => n4784);
   U305 : BUF_X1 port map( A => n4791, Z => n4792);
   U306 : BUF_X1 port map( A => n4799, Z => n4800);
   U307 : BUF_X1 port map( A => n4719, Z => n4720);
   U308 : BUF_X1 port map( A => n4735, Z => n4736);
   U309 : BUF_X1 port map( A => n4727, Z => n4728);
   U310 : BUF_X1 port map( A => n4711, Z => n4712);
   U311 : BUF_X1 port map( A => n4490, Z => n4483);
   U312 : BUF_X1 port map( A => n4490, Z => n4484);
   U313 : BUF_X1 port map( A => n4490, Z => n4485);
   U314 : BUF_X1 port map( A => n4489, Z => n4486);
   U315 : BUF_X1 port map( A => n4489, Z => n4487);
   U316 : BUF_X1 port map( A => n4554, Z => n4547);
   U317 : BUF_X1 port map( A => n4554, Z => n4548);
   U318 : BUF_X1 port map( A => n4554, Z => n4549);
   U319 : BUF_X1 port map( A => n4553, Z => n4550);
   U320 : BUF_X1 port map( A => n4553, Z => n4551);
   U321 : BUF_X1 port map( A => n4514, Z => n4507);
   U322 : BUF_X1 port map( A => n4514, Z => n4508);
   U323 : BUF_X1 port map( A => n4514, Z => n4509);
   U324 : BUF_X1 port map( A => n4513, Z => n4510);
   U325 : BUF_X1 port map( A => n4513, Z => n4511);
   U326 : BUF_X1 port map( A => n4578, Z => n4571);
   U327 : BUF_X1 port map( A => n4578, Z => n4572);
   U328 : BUF_X1 port map( A => n4578, Z => n4573);
   U329 : BUF_X1 port map( A => n4577, Z => n4574);
   U330 : BUF_X1 port map( A => n4577, Z => n4575);
   U331 : BUF_X1 port map( A => n4506, Z => n4499);
   U332 : BUF_X1 port map( A => n4506, Z => n4500);
   U333 : BUF_X1 port map( A => n4506, Z => n4501);
   U334 : BUF_X1 port map( A => n4505, Z => n4502);
   U335 : BUF_X1 port map( A => n4505, Z => n4503);
   U336 : BUF_X1 port map( A => n4570, Z => n4563);
   U337 : BUF_X1 port map( A => n4570, Z => n4564);
   U338 : BUF_X1 port map( A => n4570, Z => n4565);
   U339 : BUF_X1 port map( A => n4569, Z => n4566);
   U340 : BUF_X1 port map( A => n4569, Z => n4567);
   U341 : BUF_X1 port map( A => n4489, Z => n4488);
   U342 : BUF_X1 port map( A => n4553, Z => n4552);
   U343 : BUF_X1 port map( A => n4513, Z => n4512);
   U344 : BUF_X1 port map( A => n4577, Z => n4576);
   U345 : BUF_X1 port map( A => n4505, Z => n4504);
   U346 : BUF_X1 port map( A => n4569, Z => n4568);
   U347 : BUF_X1 port map( A => n4530, Z => n4523);
   U348 : BUF_X1 port map( A => n4530, Z => n4524);
   U349 : BUF_X1 port map( A => n4530, Z => n4525);
   U350 : BUF_X1 port map( A => n4529, Z => n4526);
   U351 : BUF_X1 port map( A => n4529, Z => n4527);
   U352 : BUF_X1 port map( A => n4522, Z => n4515);
   U353 : BUF_X1 port map( A => n4522, Z => n4516);
   U354 : BUF_X1 port map( A => n4522, Z => n4517);
   U355 : BUF_X1 port map( A => n4521, Z => n4518);
   U356 : BUF_X1 port map( A => n4521, Z => n4519);
   U357 : BUF_X1 port map( A => n4594, Z => n4587);
   U358 : BUF_X1 port map( A => n4594, Z => n4588);
   U359 : BUF_X1 port map( A => n4594, Z => n4589);
   U360 : BUF_X1 port map( A => n4593, Z => n4590);
   U361 : BUF_X1 port map( A => n4593, Z => n4591);
   U362 : BUF_X1 port map( A => n4586, Z => n4579);
   U363 : BUF_X1 port map( A => n4586, Z => n4580);
   U364 : BUF_X1 port map( A => n4586, Z => n4581);
   U365 : BUF_X1 port map( A => n4585, Z => n4582);
   U366 : BUF_X1 port map( A => n4585, Z => n4583);
   U367 : BUF_X1 port map( A => n4529, Z => n4528);
   U368 : BUF_X1 port map( A => n4521, Z => n4520);
   U369 : BUF_X1 port map( A => n4593, Z => n4592);
   U370 : BUF_X1 port map( A => n4585, Z => n4584);
   U371 : BUF_X1 port map( A => n4538, Z => n4531);
   U372 : BUF_X1 port map( A => n4538, Z => n4532);
   U373 : BUF_X1 port map( A => n4538, Z => n4533);
   U374 : BUF_X1 port map( A => n4537, Z => n4534);
   U375 : BUF_X1 port map( A => n4537, Z => n4535);
   U376 : BUF_X1 port map( A => n4602, Z => n4595);
   U377 : BUF_X1 port map( A => n4602, Z => n4596);
   U378 : BUF_X1 port map( A => n4602, Z => n4597);
   U379 : BUF_X1 port map( A => n4601, Z => n4598);
   U380 : BUF_X1 port map( A => n4601, Z => n4599);
   U381 : BUF_X1 port map( A => n4537, Z => n4536);
   U382 : BUF_X1 port map( A => n4601, Z => n4600);
   U383 : BUF_X1 port map( A => n4610, Z => n4603);
   U384 : BUF_X1 port map( A => n4610, Z => n4604);
   U385 : BUF_X1 port map( A => n4610, Z => n4605);
   U386 : BUF_X1 port map( A => n4609, Z => n4606);
   U387 : BUF_X1 port map( A => n4609, Z => n4607);
   U388 : BUF_X1 port map( A => n4546, Z => n4539);
   U389 : BUF_X1 port map( A => n4546, Z => n4540);
   U390 : BUF_X1 port map( A => n4546, Z => n4541);
   U391 : BUF_X1 port map( A => n4545, Z => n4542);
   U392 : BUF_X1 port map( A => n4545, Z => n4543);
   U393 : BUF_X1 port map( A => n4609, Z => n4608);
   U394 : BUF_X1 port map( A => n4545, Z => n4544);
   U395 : BUF_X1 port map( A => n4935, Z => n4938);
   U396 : BUF_X1 port map( A => n4943, Z => n4946);
   U397 : BUF_X1 port map( A => n4951, Z => n4954);
   U398 : BUF_X1 port map( A => n4935, Z => n4937);
   U399 : BUF_X1 port map( A => n4943, Z => n4945);
   U400 : BUF_X1 port map( A => n4951, Z => n4953);
   U401 : BUF_X1 port map( A => n4743, Z => n4746);
   U402 : BUF_X1 port map( A => n4759, Z => n4762);
   U403 : BUF_X1 port map( A => n4807, Z => n4810);
   U404 : BUF_X1 port map( A => n4823, Z => n4826);
   U405 : BUF_X1 port map( A => n4871, Z => n4874);
   U406 : BUF_X1 port map( A => n4879, Z => n4882);
   U407 : BUF_X1 port map( A => n4887, Z => n4890);
   U408 : BUF_X1 port map( A => n4895, Z => n4898);
   U409 : BUF_X1 port map( A => n4751, Z => n4754);
   U410 : BUF_X1 port map( A => n4767, Z => n4770);
   U411 : BUF_X1 port map( A => n4815, Z => n4818);
   U412 : BUF_X1 port map( A => n4831, Z => n4834);
   U413 : BUF_X1 port map( A => n4743, Z => n4745);
   U414 : BUF_X1 port map( A => n4759, Z => n4761);
   U415 : BUF_X1 port map( A => n4807, Z => n4809);
   U416 : BUF_X1 port map( A => n4823, Z => n4825);
   U417 : BUF_X1 port map( A => n4871, Z => n4873);
   U418 : BUF_X1 port map( A => n4879, Z => n4881);
   U419 : BUF_X1 port map( A => n4887, Z => n4889);
   U420 : BUF_X1 port map( A => n4895, Z => n4897);
   U421 : BUF_X1 port map( A => n4751, Z => n4753);
   U422 : BUF_X1 port map( A => n4767, Z => n4769);
   U423 : BUF_X1 port map( A => n4815, Z => n4817);
   U424 : BUF_X1 port map( A => n4831, Z => n4833);
   U425 : BUF_X1 port map( A => n4959, Z => n4961);
   U426 : BUF_X1 port map( A => n4903, Z => n4906);
   U427 : BUF_X1 port map( A => n4911, Z => n4914);
   U428 : BUF_X1 port map( A => n4919, Z => n4922);
   U429 : BUF_X1 port map( A => n4927, Z => n4930);
   U430 : BUF_X1 port map( A => n4903, Z => n4905);
   U431 : BUF_X1 port map( A => n4911, Z => n4913);
   U432 : BUF_X1 port map( A => n4919, Z => n4921);
   U433 : BUF_X1 port map( A => n4927, Z => n4929);
   U434 : BUF_X1 port map( A => n4959, Z => n4962);
   U435 : BUF_X1 port map( A => n4839, Z => n4842);
   U436 : BUF_X1 port map( A => n4847, Z => n4850);
   U437 : BUF_X1 port map( A => n4855, Z => n4858);
   U438 : BUF_X1 port map( A => n4863, Z => n4866);
   U439 : BUF_X1 port map( A => n4775, Z => n4778);
   U440 : BUF_X1 port map( A => n4783, Z => n4786);
   U441 : BUF_X1 port map( A => n4791, Z => n4794);
   U442 : BUF_X1 port map( A => n4799, Z => n4802);
   U443 : BUF_X1 port map( A => n4719, Z => n4722);
   U444 : BUF_X1 port map( A => n4735, Z => n4738);
   U445 : BUF_X1 port map( A => n4839, Z => n4841);
   U446 : BUF_X1 port map( A => n4847, Z => n4849);
   U447 : BUF_X1 port map( A => n4855, Z => n4857);
   U448 : BUF_X1 port map( A => n4863, Z => n4865);
   U449 : BUF_X1 port map( A => n4727, Z => n4730);
   U450 : BUF_X1 port map( A => n4775, Z => n4777);
   U451 : BUF_X1 port map( A => n4783, Z => n4785);
   U452 : BUF_X1 port map( A => n4791, Z => n4793);
   U453 : BUF_X1 port map( A => n4799, Z => n4801);
   U454 : BUF_X1 port map( A => n4719, Z => n4721);
   U455 : BUF_X1 port map( A => n4735, Z => n4737);
   U456 : BUF_X1 port map( A => n4727, Z => n4729);
   U457 : BUF_X1 port map( A => n4711, Z => n4714);
   U458 : BUF_X1 port map( A => n4711, Z => n4713);
   U459 : BUF_X1 port map( A => n5071, Z => n5074);
   U460 : BUF_X1 port map( A => n4991, Z => n4994);
   U461 : BUF_X1 port map( A => n5071, Z => n5072);
   U462 : BUF_X1 port map( A => n5071, Z => n5073);
   U463 : BUF_X1 port map( A => n4991, Z => n4992);
   U464 : BUF_X1 port map( A => n4991, Z => n4993);
   U465 : BUF_X1 port map( A => n5119, Z => n5120);
   U466 : BUF_X1 port map( A => n5119, Z => n5121);
   U467 : BUF_X1 port map( A => n5039, Z => n5040);
   U468 : BUF_X1 port map( A => n5039, Z => n5041);
   U469 : BUF_X1 port map( A => n5126, Z => n5123);
   U470 : BUF_X1 port map( A => n5126, Z => n5124);
   U471 : BUF_X1 port map( A => n5126, Z => n5125);
   U472 : BUF_X1 port map( A => n5119, Z => n5122);
   U473 : BUF_X1 port map( A => n5039, Z => n5042);
   U474 : NAND2_X1 port map( A1 => n2686, A2 => n2687, ZN => n2684);
   U475 : NAND2_X1 port map( A1 => n2696, A2 => n2687, ZN => n2694);
   U476 : NAND2_X1 port map( A1 => n2693, A2 => n2687, ZN => n2691);
   U477 : NAND2_X1 port map( A1 => n2690, A2 => n2687, ZN => n2688);
   U478 : NAND2_X1 port map( A1 => n2746, A2 => n2690, ZN => n2747);
   U479 : NAND2_X1 port map( A1 => n2729, A2 => n2696, ZN => n2734);
   U480 : NAND2_X1 port map( A1 => n2712, A2 => n2696, ZN => n2717);
   U481 : NAND2_X1 port map( A1 => n2712, A2 => n2693, ZN => n2715);
   U482 : NAND2_X1 port map( A1 => n2712, A2 => n2690, ZN => n2713);
   U483 : NAND2_X1 port map( A1 => n2712, A2 => n2686, ZN => n2710);
   U484 : NAND2_X1 port map( A1 => n2746, A2 => n2696, ZN => n2751);
   U485 : NAND2_X1 port map( A1 => n2746, A2 => n2693, ZN => n2749);
   U486 : NAND2_X1 port map( A1 => n2746, A2 => n2686, ZN => n2744);
   U487 : NAND2_X1 port map( A1 => n2729, A2 => n2693, ZN => n2732);
   U488 : NAND2_X1 port map( A1 => n2729, A2 => n2690, ZN => n2730);
   U489 : NAND2_X1 port map( A1 => n2729, A2 => n2686, ZN => n2727);
   U490 : NAND2_X1 port map( A1 => n2708, A2 => n2687, ZN => n2706);
   U491 : NAND2_X1 port map( A1 => n2705, A2 => n2687, ZN => n2703);
   U492 : NAND2_X1 port map( A1 => n2702, A2 => n2687, ZN => n2700);
   U493 : NAND2_X1 port map( A1 => n2699, A2 => n2687, ZN => n2697);
   U494 : NAND2_X1 port map( A1 => n2712, A2 => n2708, ZN => n2725);
   U495 : NAND2_X1 port map( A1 => n2712, A2 => n2705, ZN => n2723);
   U496 : NAND2_X1 port map( A1 => n2712, A2 => n2702, ZN => n2721);
   U497 : NAND2_X1 port map( A1 => n2712, A2 => n2699, ZN => n2719);
   U498 : NAND2_X1 port map( A1 => n2729, A2 => n2708, ZN => n2742);
   U499 : NAND2_X1 port map( A1 => n2729, A2 => n2705, ZN => n2740);
   U500 : NAND2_X1 port map( A1 => n2729, A2 => n2702, ZN => n2738);
   U501 : NAND2_X1 port map( A1 => n2729, A2 => n2699, ZN => n2736);
   U502 : NAND2_X1 port map( A1 => n2746, A2 => n2705, ZN => n2757);
   U503 : NAND2_X1 port map( A1 => n2746, A2 => n2699, ZN => n2753);
   U504 : NAND2_X1 port map( A1 => n2746, A2 => n2702, ZN => n2755);
   U505 : NAND2_X1 port map( A1 => n2746, A2 => n2708, ZN => n2759);
   U506 : INV_X1 port map( A => n1003, ZN => n5141);
   U507 : INV_X1 port map( A => n2665, ZN => n5128);
   U508 : BUF_X1 port map( A => n5007, Z => n5010);
   U509 : BUF_X1 port map( A => n5002, Z => n5001);
   U510 : BUF_X1 port map( A => n5007, Z => n5008);
   U511 : BUF_X1 port map( A => n5007, Z => n5009);
   U512 : BUF_X1 port map( A => n5002, Z => n5000);
   U513 : BUF_X1 port map( A => n5002, Z => n4999);
   U514 : BUF_X1 port map( A => n5103, Z => n5106);
   U515 : BUF_X1 port map( A => n5023, Z => n5026);
   U516 : BUF_X1 port map( A => n5103, Z => n5104);
   U517 : BUF_X1 port map( A => n5103, Z => n5105);
   U518 : BUF_X1 port map( A => n5023, Z => n5024);
   U519 : BUF_X1 port map( A => n5023, Z => n5025);
   U520 : BUF_X1 port map( A => n5102, Z => n5101);
   U521 : BUF_X1 port map( A => n5022, Z => n5021);
   U522 : BUF_X1 port map( A => n5087, Z => n5090);
   U523 : BUF_X1 port map( A => n5082, Z => n5081);
   U524 : BUF_X1 port map( A => n5102, Z => n5100);
   U525 : BUF_X1 port map( A => n5102, Z => n5099);
   U526 : BUF_X1 port map( A => n5022, Z => n5020);
   U527 : BUF_X1 port map( A => n5022, Z => n5019);
   U528 : BUF_X1 port map( A => n5087, Z => n5088);
   U529 : BUF_X1 port map( A => n5087, Z => n5089);
   U530 : BUF_X1 port map( A => n5082, Z => n5080);
   U531 : BUF_X1 port map( A => n5082, Z => n5079);
   U532 : BUF_X1 port map( A => n4970, Z => n4969);
   U533 : BUF_X1 port map( A => n4970, Z => n4968);
   U534 : BUF_X1 port map( A => n4970, Z => n4967);
   U535 : BUF_X1 port map( A => n4986, Z => n4985);
   U536 : BUF_X1 port map( A => n5067, Z => n5070);
   U537 : BUF_X1 port map( A => n4987, Z => n4990);
   U538 : BUF_X1 port map( A => n4986, Z => n4984);
   U539 : BUF_X1 port map( A => n4986, Z => n4983);
   U540 : BUF_X1 port map( A => n5067, Z => n5068);
   U541 : BUF_X1 port map( A => n5067, Z => n5069);
   U542 : BUF_X1 port map( A => n4971, Z => n4974);
   U543 : BUF_X1 port map( A => n4987, Z => n4988);
   U544 : BUF_X1 port map( A => n4987, Z => n4989);
   U545 : BUF_X1 port map( A => n4971, Z => n4972);
   U546 : BUF_X1 port map( A => n4971, Z => n4973);
   U547 : BUF_X1 port map( A => n5050, Z => n5049);
   U548 : BUF_X1 port map( A => n5050, Z => n5048);
   U549 : BUF_X1 port map( A => n5050, Z => n5047);
   U550 : BUF_X1 port map( A => n5066, Z => n5065);
   U551 : BUF_X1 port map( A => n5066, Z => n5064);
   U552 : BUF_X1 port map( A => n5066, Z => n5063);
   U553 : BUF_X1 port map( A => n5051, Z => n5054);
   U554 : BUF_X1 port map( A => n5051, Z => n5052);
   U555 : BUF_X1 port map( A => n5051, Z => n5053);
   U556 : BUF_X1 port map( A => n5046, Z => n5045);
   U557 : BUF_X1 port map( A => n4966, Z => n4965);
   U558 : BUF_X1 port map( A => n5046, Z => n5044);
   U559 : BUF_X1 port map( A => n5046, Z => n5043);
   U560 : BUF_X1 port map( A => n4966, Z => n4964);
   U561 : BUF_X1 port map( A => n4966, Z => n4963);
   U562 : BUF_X1 port map( A => n5086, Z => n5085);
   U563 : BUF_X1 port map( A => n5006, Z => n5005);
   U564 : BUF_X1 port map( A => n5086, Z => n5084);
   U565 : BUF_X1 port map( A => n5086, Z => n5083);
   U566 : BUF_X1 port map( A => n5006, Z => n5004);
   U567 : BUF_X1 port map( A => n5006, Z => n5003);
   U568 : BUF_X1 port map( A => n5095, Z => n5098);
   U569 : BUF_X1 port map( A => n5015, Z => n5018);
   U570 : BUF_X1 port map( A => n5095, Z => n5096);
   U571 : BUF_X1 port map( A => n5095, Z => n5097);
   U572 : BUF_X1 port map( A => n5015, Z => n5016);
   U573 : BUF_X1 port map( A => n5015, Z => n5017);
   U574 : BUF_X1 port map( A => n5075, Z => n5078);
   U575 : BUF_X1 port map( A => n4995, Z => n4998);
   U576 : BUF_X1 port map( A => n5075, Z => n5076);
   U577 : BUF_X1 port map( A => n5075, Z => n5077);
   U578 : BUF_X1 port map( A => n4995, Z => n4996);
   U579 : BUF_X1 port map( A => n4995, Z => n4997);
   U580 : BUF_X1 port map( A => n5091, Z => n5094);
   U581 : BUF_X1 port map( A => n5011, Z => n5014);
   U582 : BUF_X1 port map( A => n5091, Z => n5092);
   U583 : BUF_X1 port map( A => n5091, Z => n5093);
   U584 : BUF_X1 port map( A => n5011, Z => n5012);
   U585 : BUF_X1 port map( A => n5011, Z => n5013);
   U586 : BUF_X1 port map( A => n4979, Z => n4982);
   U587 : BUF_X1 port map( A => n4979, Z => n4980);
   U588 : BUF_X1 port map( A => n4979, Z => n4981);
   U589 : BUF_X1 port map( A => n5055, Z => n5058);
   U590 : BUF_X1 port map( A => n4975, Z => n4978);
   U591 : BUF_X1 port map( A => n5055, Z => n5056);
   U592 : BUF_X1 port map( A => n5055, Z => n5057);
   U593 : BUF_X1 port map( A => n4975, Z => n4976);
   U594 : BUF_X1 port map( A => n4975, Z => n4977);
   U595 : BUF_X1 port map( A => n5059, Z => n5062);
   U596 : BUF_X1 port map( A => n5059, Z => n5060);
   U597 : BUF_X1 port map( A => n5059, Z => n5061);
   U598 : NAND2_X1 port map( A1 => n1003, A2 => n1020, ZN => n413);
   U599 : NAND2_X1 port map( A1 => n2665, A2 => n2682, ZN => n1051);
   U600 : BUF_X1 port map( A => n5107, Z => n5110);
   U601 : BUF_X1 port map( A => n5027, Z => n5030);
   U602 : BUF_X1 port map( A => n5107, Z => n5108);
   U603 : BUF_X1 port map( A => n5107, Z => n5109);
   U604 : BUF_X1 port map( A => n5027, Z => n5028);
   U605 : BUF_X1 port map( A => n5027, Z => n5029);
   U606 : NAND2_X1 port map( A1 => n5125, A2 => n5116, ZN => n384);
   U607 : NAND2_X1 port map( A1 => n5125, A2 => n5036, ZN => n1022);
   U608 : INV_X1 port map( A => RESET, ZN => n5126);
   U609 : BUF_X1 port map( A => n5156, Z => n4620);
   U610 : BUF_X1 port map( A => n5157, Z => n4623);
   U611 : BUF_X1 port map( A => n5158, Z => n4626);
   U612 : BUF_X1 port map( A => n5159, Z => n4629);
   U613 : BUF_X1 port map( A => n5160, Z => n4632);
   U614 : BUF_X1 port map( A => n5161, Z => n4635);
   U615 : BUF_X1 port map( A => n5184, Z => n4704);
   U616 : BUF_X1 port map( A => n5153, Z => n4611);
   U617 : BUF_X1 port map( A => n5154, Z => n4614);
   U618 : BUF_X1 port map( A => n5155, Z => n4617);
   U619 : BUF_X1 port map( A => n5163, Z => n4641);
   U620 : BUF_X1 port map( A => n5164, Z => n4644);
   U621 : BUF_X1 port map( A => n5165, Z => n4647);
   U622 : BUF_X1 port map( A => n5166, Z => n4650);
   U623 : BUF_X1 port map( A => n5167, Z => n4653);
   U624 : BUF_X1 port map( A => n5168, Z => n4656);
   U625 : BUF_X1 port map( A => n5169, Z => n4659);
   U626 : BUF_X1 port map( A => n5170, Z => n4662);
   U627 : BUF_X1 port map( A => n5171, Z => n4665);
   U628 : BUF_X1 port map( A => n5172, Z => n4668);
   U629 : BUF_X1 port map( A => n5173, Z => n4671);
   U630 : BUF_X1 port map( A => n5174, Z => n4674);
   U631 : BUF_X1 port map( A => n5175, Z => n4677);
   U632 : BUF_X1 port map( A => n5176, Z => n4680);
   U633 : BUF_X1 port map( A => n5177, Z => n4683);
   U634 : BUF_X1 port map( A => n5178, Z => n4686);
   U635 : BUF_X1 port map( A => n5179, Z => n4689);
   U636 : BUF_X1 port map( A => n5180, Z => n4692);
   U637 : BUF_X1 port map( A => n5181, Z => n4695);
   U638 : BUF_X1 port map( A => n5182, Z => n4698);
   U639 : BUF_X1 port map( A => n5183, Z => n4701);
   U640 : BUF_X1 port map( A => n5156, Z => n4621);
   U641 : BUF_X1 port map( A => n5157, Z => n4624);
   U642 : BUF_X1 port map( A => n5158, Z => n4627);
   U643 : BUF_X1 port map( A => n5159, Z => n4630);
   U644 : BUF_X1 port map( A => n5160, Z => n4633);
   U645 : BUF_X1 port map( A => n5161, Z => n4636);
   U646 : BUF_X1 port map( A => n5184, Z => n4705);
   U647 : BUF_X1 port map( A => n5153, Z => n4612);
   U648 : BUF_X1 port map( A => n5154, Z => n4615);
   U649 : BUF_X1 port map( A => n5155, Z => n4618);
   U650 : BUF_X1 port map( A => n5163, Z => n4642);
   U651 : BUF_X1 port map( A => n5164, Z => n4645);
   U652 : BUF_X1 port map( A => n5165, Z => n4648);
   U653 : BUF_X1 port map( A => n5166, Z => n4651);
   U654 : BUF_X1 port map( A => n5167, Z => n4654);
   U655 : BUF_X1 port map( A => n5168, Z => n4657);
   U656 : BUF_X1 port map( A => n5169, Z => n4660);
   U657 : BUF_X1 port map( A => n5170, Z => n4663);
   U658 : BUF_X1 port map( A => n5171, Z => n4666);
   U659 : BUF_X1 port map( A => n5172, Z => n4669);
   U660 : BUF_X1 port map( A => n5173, Z => n4672);
   U661 : BUF_X1 port map( A => n5174, Z => n4675);
   U662 : BUF_X1 port map( A => n5175, Z => n4678);
   U663 : BUF_X1 port map( A => n5176, Z => n4681);
   U664 : BUF_X1 port map( A => n5177, Z => n4684);
   U665 : BUF_X1 port map( A => n5178, Z => n4687);
   U666 : BUF_X1 port map( A => n5179, Z => n4690);
   U667 : BUF_X1 port map( A => n5180, Z => n4693);
   U668 : BUF_X1 port map( A => n5181, Z => n4696);
   U669 : BUF_X1 port map( A => n5182, Z => n4699);
   U670 : BUF_X1 port map( A => n5183, Z => n4702);
   U671 : BUF_X1 port map( A => n5162, Z => n4638);
   U672 : BUF_X1 port map( A => n5162, Z => n4639);
   U673 : BUF_X1 port map( A => n5156, Z => n4622);
   U674 : BUF_X1 port map( A => n5157, Z => n4625);
   U675 : BUF_X1 port map( A => n5158, Z => n4628);
   U676 : BUF_X1 port map( A => n5159, Z => n4631);
   U677 : BUF_X1 port map( A => n5160, Z => n4634);
   U678 : BUF_X1 port map( A => n5161, Z => n4637);
   U679 : BUF_X1 port map( A => n5184, Z => n4706);
   U680 : BUF_X1 port map( A => n5153, Z => n4613);
   U681 : BUF_X1 port map( A => n5154, Z => n4616);
   U682 : BUF_X1 port map( A => n5155, Z => n4619);
   U683 : BUF_X1 port map( A => n5163, Z => n4643);
   U684 : BUF_X1 port map( A => n5164, Z => n4646);
   U685 : BUF_X1 port map( A => n5165, Z => n4649);
   U686 : BUF_X1 port map( A => n5166, Z => n4652);
   U687 : BUF_X1 port map( A => n5167, Z => n4655);
   U688 : BUF_X1 port map( A => n5168, Z => n4658);
   U689 : BUF_X1 port map( A => n5169, Z => n4661);
   U690 : BUF_X1 port map( A => n5170, Z => n4664);
   U691 : BUF_X1 port map( A => n5171, Z => n4667);
   U692 : BUF_X1 port map( A => n5172, Z => n4670);
   U693 : BUF_X1 port map( A => n5173, Z => n4673);
   U694 : BUF_X1 port map( A => n5174, Z => n4676);
   U695 : BUF_X1 port map( A => n5175, Z => n4679);
   U696 : BUF_X1 port map( A => n5176, Z => n4682);
   U697 : BUF_X1 port map( A => n5177, Z => n4685);
   U698 : BUF_X1 port map( A => n5178, Z => n4688);
   U699 : BUF_X1 port map( A => n5179, Z => n4691);
   U700 : BUF_X1 port map( A => n5180, Z => n4694);
   U701 : BUF_X1 port map( A => n5181, Z => n4697);
   U702 : BUF_X1 port map( A => n5182, Z => n4700);
   U703 : BUF_X1 port map( A => n5183, Z => n4703);
   U704 : BUF_X1 port map( A => n5162, Z => n4640);
   U705 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => ADD_WR(0), 
                           ZN => n2686);
   U706 : NOR3_X1 port map( A1 => n5185, A2 => ADD_WR(2), A3 => n5186, ZN => 
                           n2696);
   U707 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n5186, ZN 
                           => n2693);
   U708 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n5185, ZN 
                           => n2690);
   U709 : AND3_X1 port map( A1 => n5187, A2 => n5188, A3 => n2709, ZN => n2687)
                           ;
   U710 : INV_X1 port map( A => ADD_WR(4), ZN => n5188);
   U711 : INV_X1 port map( A => ADD_WR(3), ZN => n5187);
   U712 : INV_X1 port map( A => ADD_WR(1), ZN => n5186);
   U713 : INV_X1 port map( A => ADD_WR(0), ZN => n5185);
   U714 : AND3_X1 port map( A1 => n2709, A2 => n5187, A3 => ADD_WR(4), ZN => 
                           n2729);
   U715 : AND3_X1 port map( A1 => n2709, A2 => n5188, A3 => ADD_WR(3), ZN => 
                           n2712);
   U716 : AND3_X1 port map( A1 => ADD_WR(1), A2 => n5185, A3 => ADD_WR(2), ZN 
                           => n2705);
   U717 : AND3_X1 port map( A1 => n5185, A2 => n5186, A3 => ADD_WR(2), ZN => 
                           n2699);
   U718 : AND3_X1 port map( A1 => ADD_WR(0), A2 => n5186, A3 => ADD_WR(2), ZN 
                           => n2702);
   U719 : AND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2), 
                           ZN => n2708);
   U720 : AND3_X1 port map( A1 => ADD_WR(3), A2 => n2709, A3 => ADD_WR(4), ZN 
                           => n2746);
   U721 : OAI221_X1 port map( B1 => n2660, B2 => n5032, C1 => n2661, C2 => 
                           n5028, A => n2662, ZN => n2659);
   U722 : AOI22_X1 port map( A1 => n5024, A2 => n4387, B1 => n5021, B2 => n4291
                           , ZN => n2662);
   U723 : NOR4_X1 port map( A1 => n2666, A2 => n2667, A3 => n2668, A4 => n2669,
                           ZN => n2661);
   U724 : NOR4_X1 port map( A1 => n2670, A2 => n2671, A3 => n2672, A4 => n2673,
                           ZN => n2660);
   U725 : OAI221_X1 port map( B1 => n2641, B2 => n5032, C1 => n2642, C2 => 
                           n5028, A => n2643, ZN => n2640);
   U726 : AOI22_X1 port map( A1 => n5024, A2 => n4388, B1 => n5021, B2 => n4292
                           , ZN => n2643);
   U727 : NOR4_X1 port map( A1 => n2644, A2 => n2645, A3 => n2646, A4 => n2647,
                           ZN => n2642);
   U728 : NOR4_X1 port map( A1 => n2648, A2 => n2649, A3 => n2650, A4 => n2651,
                           ZN => n2641);
   U729 : OAI221_X1 port map( B1 => n2622, B2 => n5032, C1 => n2623, C2 => 
                           n5028, A => n2624, ZN => n2621);
   U730 : AOI22_X1 port map( A1 => n5024, A2 => n4389, B1 => n5021, B2 => n4293
                           , ZN => n2624);
   U731 : NOR4_X1 port map( A1 => n2625, A2 => n2626, A3 => n2627, A4 => n2628,
                           ZN => n2623);
   U732 : NOR4_X1 port map( A1 => n2629, A2 => n2630, A3 => n2631, A4 => n2632,
                           ZN => n2622);
   U733 : OAI221_X1 port map( B1 => n2603, B2 => n5032, C1 => n2604, C2 => 
                           n5028, A => n2605, ZN => n2602);
   U734 : AOI22_X1 port map( A1 => n5024, A2 => n4390, B1 => n5021, B2 => n4294
                           , ZN => n2605);
   U735 : NOR4_X1 port map( A1 => n2606, A2 => n2607, A3 => n2608, A4 => n2609,
                           ZN => n2604);
   U736 : NOR4_X1 port map( A1 => n2610, A2 => n2611, A3 => n2612, A4 => n2613,
                           ZN => n2603);
   U737 : OAI221_X1 port map( B1 => n2584, B2 => n5032, C1 => n2585, C2 => 
                           n5028, A => n2586, ZN => n2583);
   U738 : AOI22_X1 port map( A1 => n5024, A2 => n4391, B1 => n5021, B2 => n4295
                           , ZN => n2586);
   U739 : NOR4_X1 port map( A1 => n2587, A2 => n2588, A3 => n2589, A4 => n2590,
                           ZN => n2585);
   U740 : NOR4_X1 port map( A1 => n2591, A2 => n2592, A3 => n2593, A4 => n2594,
                           ZN => n2584);
   U741 : OAI221_X1 port map( B1 => n2565, B2 => n5032, C1 => n2566, C2 => 
                           n5028, A => n2567, ZN => n2564);
   U742 : AOI22_X1 port map( A1 => n5024, A2 => n4392, B1 => n5021, B2 => n4296
                           , ZN => n2567);
   U743 : NOR4_X1 port map( A1 => n2568, A2 => n2569, A3 => n2570, A4 => n2571,
                           ZN => n2566);
   U744 : NOR4_X1 port map( A1 => n2572, A2 => n2573, A3 => n2574, A4 => n2575,
                           ZN => n2565);
   U745 : OAI221_X1 port map( B1 => n2546, B2 => n5032, C1 => n2547, C2 => 
                           n5028, A => n2548, ZN => n2545);
   U746 : AOI22_X1 port map( A1 => n5024, A2 => n4393, B1 => n5021, B2 => n4297
                           , ZN => n2548);
   U747 : NOR4_X1 port map( A1 => n2549, A2 => n2550, A3 => n2551, A4 => n2552,
                           ZN => n2547);
   U748 : NOR4_X1 port map( A1 => n2553, A2 => n2554, A3 => n2555, A4 => n2556,
                           ZN => n2546);
   U749 : OAI221_X1 port map( B1 => n2527, B2 => n5032, C1 => n2528, C2 => 
                           n5028, A => n2529, ZN => n2526);
   U750 : AOI22_X1 port map( A1 => n5024, A2 => n4394, B1 => n5021, B2 => n4298
                           , ZN => n2529);
   U751 : NOR4_X1 port map( A1 => n2530, A2 => n2531, A3 => n2532, A4 => n2533,
                           ZN => n2528);
   U752 : NOR4_X1 port map( A1 => n2534, A2 => n2535, A3 => n2536, A4 => n2537,
                           ZN => n2527);
   U753 : OAI221_X1 port map( B1 => n2508, B2 => n5032, C1 => n2509, C2 => 
                           n5028, A => n2510, ZN => n2507);
   U754 : AOI22_X1 port map( A1 => n5024, A2 => n4395, B1 => n5020, B2 => n4299
                           , ZN => n2510);
   U755 : NOR4_X1 port map( A1 => n2511, A2 => n2512, A3 => n2513, A4 => n2514,
                           ZN => n2509);
   U756 : NOR4_X1 port map( A1 => n2515, A2 => n2516, A3 => n2517, A4 => n2518,
                           ZN => n2508);
   U757 : OAI221_X1 port map( B1 => n2489, B2 => n5032, C1 => n2490, C2 => 
                           n5028, A => n2491, ZN => n2488);
   U758 : AOI22_X1 port map( A1 => n5024, A2 => n4396, B1 => n5020, B2 => n4300
                           , ZN => n2491);
   U759 : NOR4_X1 port map( A1 => n2492, A2 => n2493, A3 => n2494, A4 => n2495,
                           ZN => n2490);
   U760 : NOR4_X1 port map( A1 => n2496, A2 => n2497, A3 => n2498, A4 => n2499,
                           ZN => n2489);
   U761 : OAI221_X1 port map( B1 => n2470, B2 => n5032, C1 => n2471, C2 => 
                           n5028, A => n2472, ZN => n2469);
   U762 : AOI22_X1 port map( A1 => n5024, A2 => n4397, B1 => n5020, B2 => n4301
                           , ZN => n2472);
   U763 : NOR4_X1 port map( A1 => n2473, A2 => n2474, A3 => n2475, A4 => n2476,
                           ZN => n2471);
   U764 : NOR4_X1 port map( A1 => n2477, A2 => n2478, A3 => n2479, A4 => n2480,
                           ZN => n2470);
   U765 : OAI221_X1 port map( B1 => n2451, B2 => n5032, C1 => n2452, C2 => 
                           n5028, A => n2453, ZN => n2450);
   U766 : AOI22_X1 port map( A1 => n5024, A2 => n4398, B1 => n5020, B2 => n4302
                           , ZN => n2453);
   U767 : NOR4_X1 port map( A1 => n2454, A2 => n2455, A3 => n2456, A4 => n2457,
                           ZN => n2452);
   U768 : NOR4_X1 port map( A1 => n2458, A2 => n2459, A3 => n2460, A4 => n2461,
                           ZN => n2451);
   U769 : OAI221_X1 port map( B1 => n2432, B2 => n5033, C1 => n2433, C2 => 
                           n5029, A => n2434, ZN => n2431);
   U770 : AOI22_X1 port map( A1 => n5025, A2 => n4399, B1 => n5020, B2 => n4303
                           , ZN => n2434);
   U771 : NOR4_X1 port map( A1 => n2435, A2 => n2436, A3 => n2437, A4 => n2438,
                           ZN => n2433);
   U772 : NOR4_X1 port map( A1 => n2439, A2 => n2440, A3 => n2441, A4 => n2442,
                           ZN => n2432);
   U773 : OAI221_X1 port map( B1 => n2413, B2 => n5033, C1 => n2414, C2 => 
                           n5029, A => n2415, ZN => n2412);
   U774 : AOI22_X1 port map( A1 => n5025, A2 => n4400, B1 => n5020, B2 => n4304
                           , ZN => n2415);
   U775 : NOR4_X1 port map( A1 => n2416, A2 => n2417, A3 => n2418, A4 => n2419,
                           ZN => n2414);
   U776 : NOR4_X1 port map( A1 => n2420, A2 => n2421, A3 => n2422, A4 => n2423,
                           ZN => n2413);
   U777 : OAI221_X1 port map( B1 => n2394, B2 => n5033, C1 => n2395, C2 => 
                           n5029, A => n2396, ZN => n2393);
   U778 : AOI22_X1 port map( A1 => n5025, A2 => n4401, B1 => n5020, B2 => n4305
                           , ZN => n2396);
   U779 : NOR4_X1 port map( A1 => n2397, A2 => n2398, A3 => n2399, A4 => n2400,
                           ZN => n2395);
   U780 : NOR4_X1 port map( A1 => n2401, A2 => n2402, A3 => n2403, A4 => n2404,
                           ZN => n2394);
   U781 : OAI221_X1 port map( B1 => n2375, B2 => n5033, C1 => n2376, C2 => 
                           n5029, A => n2377, ZN => n2374);
   U782 : AOI22_X1 port map( A1 => n5025, A2 => n4402, B1 => n5020, B2 => n4306
                           , ZN => n2377);
   U783 : NOR4_X1 port map( A1 => n2378, A2 => n2379, A3 => n2380, A4 => n2381,
                           ZN => n2376);
   U784 : NOR4_X1 port map( A1 => n2382, A2 => n2383, A3 => n2384, A4 => n2385,
                           ZN => n2375);
   U785 : OAI221_X1 port map( B1 => n2356, B2 => n5033, C1 => n2357, C2 => 
                           n5029, A => n2358, ZN => n2355);
   U786 : AOI22_X1 port map( A1 => n5025, A2 => n4403, B1 => n5020, B2 => n4307
                           , ZN => n2358);
   U787 : NOR4_X1 port map( A1 => n2359, A2 => n2360, A3 => n2361, A4 => n2362,
                           ZN => n2357);
   U788 : NOR4_X1 port map( A1 => n2363, A2 => n2364, A3 => n2365, A4 => n2366,
                           ZN => n2356);
   U789 : OAI221_X1 port map( B1 => n2337, B2 => n5033, C1 => n2338, C2 => 
                           n5029, A => n2339, ZN => n2336);
   U790 : AOI22_X1 port map( A1 => n5025, A2 => n4404, B1 => n5020, B2 => n4308
                           , ZN => n2339);
   U791 : NOR4_X1 port map( A1 => n2340, A2 => n2341, A3 => n2342, A4 => n2343,
                           ZN => n2338);
   U792 : NOR4_X1 port map( A1 => n2344, A2 => n2345, A3 => n2346, A4 => n2347,
                           ZN => n2337);
   U793 : OAI221_X1 port map( B1 => n1294, B2 => n5033, C1 => n1295, C2 => 
                           n5029, A => n1296, ZN => n1293);
   U794 : AOI22_X1 port map( A1 => n5025, A2 => n4405, B1 => n5020, B2 => n4309
                           , ZN => n1296);
   U795 : NOR4_X1 port map( A1 => n1297, A2 => n1298, A3 => n1299, A4 => n1300,
                           ZN => n1295);
   U796 : NOR4_X1 port map( A1 => n1301, A2 => n1302, A3 => n2327, A4 => n2328,
                           ZN => n1294);
   U797 : OAI221_X1 port map( B1 => n1275, B2 => n5033, C1 => n1276, C2 => 
                           n5029, A => n1277, ZN => n1274);
   U798 : AOI22_X1 port map( A1 => n5025, A2 => n4406, B1 => n5020, B2 => n4310
                           , ZN => n1277);
   U799 : NOR4_X1 port map( A1 => n1278, A2 => n1279, A3 => n1280, A4 => n1281,
                           ZN => n1276);
   U800 : NOR4_X1 port map( A1 => n1282, A2 => n1283, A3 => n1284, A4 => n1285,
                           ZN => n1275);
   U801 : OAI221_X1 port map( B1 => n1256, B2 => n5033, C1 => n1257, C2 => 
                           n5029, A => n1258, ZN => n1255);
   U802 : AOI22_X1 port map( A1 => n5025, A2 => n4407, B1 => n5019, B2 => n4311
                           , ZN => n1258);
   U803 : NOR4_X1 port map( A1 => n1259, A2 => n1260, A3 => n1261, A4 => n1262,
                           ZN => n1257);
   U804 : NOR4_X1 port map( A1 => n1263, A2 => n1264, A3 => n1265, A4 => n1266,
                           ZN => n1256);
   U805 : OAI221_X1 port map( B1 => n1237, B2 => n5033, C1 => n1238, C2 => 
                           n5029, A => n1239, ZN => n1236);
   U806 : AOI22_X1 port map( A1 => n5025, A2 => n4408, B1 => n5019, B2 => n4312
                           , ZN => n1239);
   U807 : NOR4_X1 port map( A1 => n1240, A2 => n1241, A3 => n1242, A4 => n1243,
                           ZN => n1238);
   U808 : NOR4_X1 port map( A1 => n1244, A2 => n1245, A3 => n1246, A4 => n1247,
                           ZN => n1237);
   U809 : OAI221_X1 port map( B1 => n1218, B2 => n5033, C1 => n1219, C2 => 
                           n5029, A => n1220, ZN => n1217);
   U810 : AOI22_X1 port map( A1 => n5025, A2 => n4409, B1 => n5019, B2 => n4313
                           , ZN => n1220);
   U811 : NOR4_X1 port map( A1 => n1221, A2 => n1222, A3 => n1223, A4 => n1224,
                           ZN => n1219);
   U812 : NOR4_X1 port map( A1 => n1225, A2 => n1226, A3 => n1227, A4 => n1228,
                           ZN => n1218);
   U813 : OAI221_X1 port map( B1 => n1199, B2 => n5033, C1 => n1200, C2 => 
                           n5029, A => n1201, ZN => n1198);
   U814 : AOI22_X1 port map( A1 => n5025, A2 => n4410, B1 => n5019, B2 => n4314
                           , ZN => n1201);
   U815 : NOR4_X1 port map( A1 => n1202, A2 => n1203, A3 => n1204, A4 => n1205,
                           ZN => n1200);
   U816 : NOR4_X1 port map( A1 => n1206, A2 => n1207, A3 => n1208, A4 => n1209,
                           ZN => n1199);
   U817 : OAI221_X1 port map( B1 => n1180, B2 => n5034, C1 => n1181, C2 => 
                           n5030, A => n1182, ZN => n1179);
   U818 : AOI22_X1 port map( A1 => n5026, A2 => n4411, B1 => n5019, B2 => n4315
                           , ZN => n1182);
   U819 : NOR4_X1 port map( A1 => n1183, A2 => n1184, A3 => n1185, A4 => n1186,
                           ZN => n1181);
   U820 : NOR4_X1 port map( A1 => n1187, A2 => n1188, A3 => n1189, A4 => n1190,
                           ZN => n1180);
   U821 : OAI221_X1 port map( B1 => n1161, B2 => n5034, C1 => n1162, C2 => 
                           n5030, A => n1163, ZN => n1160);
   U822 : AOI22_X1 port map( A1 => n5026, A2 => n4412, B1 => n5019, B2 => n4316
                           , ZN => n1163);
   U823 : NOR4_X1 port map( A1 => n1164, A2 => n1165, A3 => n1166, A4 => n1167,
                           ZN => n1162);
   U824 : NOR4_X1 port map( A1 => n1168, A2 => n1169, A3 => n1170, A4 => n1171,
                           ZN => n1161);
   U825 : OAI221_X1 port map( B1 => n1142, B2 => n5034, C1 => n1143, C2 => 
                           n5030, A => n1144, ZN => n1141);
   U826 : AOI22_X1 port map( A1 => n5026, A2 => n4413, B1 => n5019, B2 => n4317
                           , ZN => n1144);
   U827 : NOR4_X1 port map( A1 => n1145, A2 => n1146, A3 => n1147, A4 => n1148,
                           ZN => n1143);
   U828 : NOR4_X1 port map( A1 => n1149, A2 => n1150, A3 => n1151, A4 => n1152,
                           ZN => n1142);
   U829 : OAI221_X1 port map( B1 => n1123, B2 => n5034, C1 => n1124, C2 => 
                           n5030, A => n1125, ZN => n1122);
   U830 : AOI22_X1 port map( A1 => n5026, A2 => n4414, B1 => n5019, B2 => n4318
                           , ZN => n1125);
   U831 : NOR4_X1 port map( A1 => n1126, A2 => n1127, A3 => n1128, A4 => n1129,
                           ZN => n1124);
   U832 : NOR4_X1 port map( A1 => n1130, A2 => n1131, A3 => n1132, A4 => n1133,
                           ZN => n1123);
   U833 : OAI221_X1 port map( B1 => n1104, B2 => n5034, C1 => n1105, C2 => 
                           n5030, A => n1106, ZN => n1103);
   U834 : AOI22_X1 port map( A1 => n5026, A2 => n4415, B1 => n5019, B2 => n4319
                           , ZN => n1106);
   U835 : NOR4_X1 port map( A1 => n1107, A2 => n1108, A3 => n1109, A4 => n1110,
                           ZN => n1105);
   U836 : NOR4_X1 port map( A1 => n1111, A2 => n1112, A3 => n1113, A4 => n1114,
                           ZN => n1104);
   U837 : OAI221_X1 port map( B1 => n1085, B2 => n5034, C1 => n1086, C2 => 
                           n5030, A => n1087, ZN => n1084);
   U838 : AOI22_X1 port map( A1 => n5026, A2 => n4416, B1 => n5019, B2 => n4320
                           , ZN => n1087);
   U839 : NOR4_X1 port map( A1 => n1088, A2 => n1089, A3 => n1090, A4 => n1091,
                           ZN => n1086);
   U840 : NOR4_X1 port map( A1 => n1092, A2 => n1093, A3 => n1094, A4 => n1095,
                           ZN => n1085);
   U841 : INV_X1 port map( A => n2664, ZN => n5127);
   U842 : OAI221_X1 port map( B1 => n998, B2 => n5112, C1 => n999, C2 => n5108,
                           A => n1000, ZN => n997);
   U843 : AOI22_X1 port map( A1 => n5104, A2 => n4387, B1 => n5101, B2 => n4291
                           , ZN => n1000);
   U844 : NOR4_X1 port map( A1 => n1004, A2 => n1005, A3 => n1006, A4 => n1007,
                           ZN => n999);
   U845 : NOR4_X1 port map( A1 => n1008, A2 => n1009, A3 => n1010, A4 => n1011,
                           ZN => n998);
   U846 : OAI221_X1 port map( B1 => n979, B2 => n5112, C1 => n980, C2 => n5108,
                           A => n981, ZN => n978);
   U847 : AOI22_X1 port map( A1 => n5104, A2 => n4388, B1 => n5101, B2 => n4292
                           , ZN => n981);
   U848 : NOR4_X1 port map( A1 => n982, A2 => n983, A3 => n984, A4 => n985, ZN 
                           => n980);
   U849 : NOR4_X1 port map( A1 => n986, A2 => n987, A3 => n988, A4 => n989, ZN 
                           => n979);
   U850 : OAI221_X1 port map( B1 => n960, B2 => n5112, C1 => n961, C2 => n5108,
                           A => n962, ZN => n959);
   U851 : AOI22_X1 port map( A1 => n5104, A2 => n4389, B1 => n5101, B2 => n4293
                           , ZN => n962);
   U852 : NOR4_X1 port map( A1 => n963, A2 => n964, A3 => n965, A4 => n966, ZN 
                           => n961);
   U853 : NOR4_X1 port map( A1 => n967, A2 => n968, A3 => n969, A4 => n970, ZN 
                           => n960);
   U854 : OAI221_X1 port map( B1 => n941, B2 => n5112, C1 => n942, C2 => n5108,
                           A => n943, ZN => n940);
   U855 : AOI22_X1 port map( A1 => n5104, A2 => n4390, B1 => n5101, B2 => n4294
                           , ZN => n943);
   U856 : NOR4_X1 port map( A1 => n944, A2 => n945, A3 => n946, A4 => n947, ZN 
                           => n942);
   U857 : NOR4_X1 port map( A1 => n948, A2 => n949, A3 => n950, A4 => n951, ZN 
                           => n941);
   U858 : OAI221_X1 port map( B1 => n922, B2 => n5112, C1 => n923, C2 => n5108,
                           A => n924, ZN => n921);
   U859 : AOI22_X1 port map( A1 => n5104, A2 => n4391, B1 => n5101, B2 => n4295
                           , ZN => n924);
   U860 : NOR4_X1 port map( A1 => n925, A2 => n926, A3 => n927, A4 => n928, ZN 
                           => n923);
   U861 : NOR4_X1 port map( A1 => n929, A2 => n930, A3 => n931, A4 => n932, ZN 
                           => n922);
   U862 : OAI221_X1 port map( B1 => n903, B2 => n5112, C1 => n904, C2 => n5108,
                           A => n905, ZN => n902);
   U863 : AOI22_X1 port map( A1 => n5104, A2 => n4392, B1 => n5101, B2 => n4296
                           , ZN => n905);
   U864 : NOR4_X1 port map( A1 => n906, A2 => n907, A3 => n908, A4 => n909, ZN 
                           => n904);
   U865 : NOR4_X1 port map( A1 => n910, A2 => n911, A3 => n912, A4 => n913, ZN 
                           => n903);
   U866 : OAI221_X1 port map( B1 => n884, B2 => n5112, C1 => n885, C2 => n5108,
                           A => n886, ZN => n883);
   U867 : AOI22_X1 port map( A1 => n5104, A2 => n4393, B1 => n5101, B2 => n4297
                           , ZN => n886);
   U868 : NOR4_X1 port map( A1 => n887, A2 => n888, A3 => n889, A4 => n890, ZN 
                           => n885);
   U869 : NOR4_X1 port map( A1 => n891, A2 => n892, A3 => n893, A4 => n894, ZN 
                           => n884);
   U870 : OAI221_X1 port map( B1 => n865, B2 => n5112, C1 => n866, C2 => n5108,
                           A => n867, ZN => n864);
   U871 : AOI22_X1 port map( A1 => n5104, A2 => n4394, B1 => n5101, B2 => n4298
                           , ZN => n867);
   U872 : NOR4_X1 port map( A1 => n868, A2 => n869, A3 => n870, A4 => n871, ZN 
                           => n866);
   U873 : NOR4_X1 port map( A1 => n872, A2 => n873, A3 => n874, A4 => n875, ZN 
                           => n865);
   U874 : OAI221_X1 port map( B1 => n846, B2 => n5112, C1 => n847, C2 => n5108,
                           A => n848, ZN => n845);
   U875 : AOI22_X1 port map( A1 => n5104, A2 => n4395, B1 => n5100, B2 => n4299
                           , ZN => n848);
   U876 : NOR4_X1 port map( A1 => n849, A2 => n850, A3 => n851, A4 => n852, ZN 
                           => n847);
   U877 : NOR4_X1 port map( A1 => n853, A2 => n854, A3 => n855, A4 => n856, ZN 
                           => n846);
   U878 : OAI221_X1 port map( B1 => n827, B2 => n5112, C1 => n828, C2 => n5108,
                           A => n829, ZN => n826);
   U879 : AOI22_X1 port map( A1 => n5104, A2 => n4396, B1 => n5100, B2 => n4300
                           , ZN => n829);
   U880 : NOR4_X1 port map( A1 => n830, A2 => n831, A3 => n832, A4 => n833, ZN 
                           => n828);
   U881 : NOR4_X1 port map( A1 => n834, A2 => n835, A3 => n836, A4 => n837, ZN 
                           => n827);
   U882 : OAI221_X1 port map( B1 => n808, B2 => n5112, C1 => n809, C2 => n5108,
                           A => n810, ZN => n807);
   U883 : AOI22_X1 port map( A1 => n5104, A2 => n4397, B1 => n5100, B2 => n4301
                           , ZN => n810);
   U884 : NOR4_X1 port map( A1 => n811, A2 => n812, A3 => n813, A4 => n814, ZN 
                           => n809);
   U885 : NOR4_X1 port map( A1 => n815, A2 => n816, A3 => n817, A4 => n818, ZN 
                           => n808);
   U886 : OAI221_X1 port map( B1 => n789, B2 => n5112, C1 => n790, C2 => n5108,
                           A => n791, ZN => n788);
   U887 : AOI22_X1 port map( A1 => n5104, A2 => n4398, B1 => n5100, B2 => n4302
                           , ZN => n791);
   U888 : NOR4_X1 port map( A1 => n792, A2 => n793, A3 => n794, A4 => n795, ZN 
                           => n790);
   U889 : NOR4_X1 port map( A1 => n796, A2 => n797, A3 => n798, A4 => n799, ZN 
                           => n789);
   U890 : OAI221_X1 port map( B1 => n770, B2 => n5113, C1 => n771, C2 => n5109,
                           A => n772, ZN => n769);
   U891 : AOI22_X1 port map( A1 => n5105, A2 => n4399, B1 => n5100, B2 => n4303
                           , ZN => n772);
   U892 : NOR4_X1 port map( A1 => n773, A2 => n774, A3 => n775, A4 => n776, ZN 
                           => n771);
   U893 : NOR4_X1 port map( A1 => n777, A2 => n778, A3 => n779, A4 => n780, ZN 
                           => n770);
   U894 : OAI221_X1 port map( B1 => n751, B2 => n5113, C1 => n752, C2 => n5109,
                           A => n753, ZN => n750);
   U895 : AOI22_X1 port map( A1 => n5105, A2 => n4400, B1 => n5100, B2 => n4304
                           , ZN => n753);
   U896 : NOR4_X1 port map( A1 => n754, A2 => n755, A3 => n756, A4 => n757, ZN 
                           => n752);
   U897 : NOR4_X1 port map( A1 => n758, A2 => n759, A3 => n760, A4 => n761, ZN 
                           => n751);
   U898 : OAI221_X1 port map( B1 => n732, B2 => n5113, C1 => n733, C2 => n5109,
                           A => n734, ZN => n731);
   U899 : AOI22_X1 port map( A1 => n5105, A2 => n4401, B1 => n5100, B2 => n4305
                           , ZN => n734);
   U900 : NOR4_X1 port map( A1 => n735, A2 => n736, A3 => n737, A4 => n738, ZN 
                           => n733);
   U901 : NOR4_X1 port map( A1 => n739, A2 => n740, A3 => n741, A4 => n742, ZN 
                           => n732);
   U902 : OAI221_X1 port map( B1 => n713, B2 => n5113, C1 => n714, C2 => n5109,
                           A => n715, ZN => n712);
   U903 : AOI22_X1 port map( A1 => n5105, A2 => n4402, B1 => n5100, B2 => n4306
                           , ZN => n715);
   U904 : NOR4_X1 port map( A1 => n716, A2 => n717, A3 => n718, A4 => n719, ZN 
                           => n714);
   U905 : NOR4_X1 port map( A1 => n720, A2 => n721, A3 => n722, A4 => n723, ZN 
                           => n713);
   U906 : OAI221_X1 port map( B1 => n694, B2 => n5113, C1 => n695, C2 => n5109,
                           A => n696, ZN => n693);
   U907 : AOI22_X1 port map( A1 => n5105, A2 => n4403, B1 => n5100, B2 => n4307
                           , ZN => n696);
   U908 : NOR4_X1 port map( A1 => n697, A2 => n698, A3 => n699, A4 => n700, ZN 
                           => n695);
   U909 : NOR4_X1 port map( A1 => n701, A2 => n702, A3 => n703, A4 => n704, ZN 
                           => n694);
   U910 : OAI221_X1 port map( B1 => n675, B2 => n5113, C1 => n676, C2 => n5109,
                           A => n677, ZN => n674);
   U911 : AOI22_X1 port map( A1 => n5105, A2 => n4404, B1 => n5100, B2 => n4308
                           , ZN => n677);
   U912 : NOR4_X1 port map( A1 => n678, A2 => n679, A3 => n680, A4 => n681, ZN 
                           => n676);
   U913 : NOR4_X1 port map( A1 => n682, A2 => n683, A3 => n684, A4 => n685, ZN 
                           => n675);
   U914 : OAI221_X1 port map( B1 => n656, B2 => n5113, C1 => n657, C2 => n5109,
                           A => n658, ZN => n655);
   U915 : AOI22_X1 port map( A1 => n5105, A2 => n4405, B1 => n5100, B2 => n4309
                           , ZN => n658);
   U916 : NOR4_X1 port map( A1 => n659, A2 => n660, A3 => n661, A4 => n662, ZN 
                           => n657);
   U917 : NOR4_X1 port map( A1 => n663, A2 => n664, A3 => n665, A4 => n666, ZN 
                           => n656);
   U918 : OAI221_X1 port map( B1 => n637, B2 => n5113, C1 => n638, C2 => n5109,
                           A => n639, ZN => n636);
   U919 : AOI22_X1 port map( A1 => n5105, A2 => n4406, B1 => n5100, B2 => n4310
                           , ZN => n639);
   U920 : NOR4_X1 port map( A1 => n640, A2 => n641, A3 => n642, A4 => n643, ZN 
                           => n638);
   U921 : NOR4_X1 port map( A1 => n644, A2 => n645, A3 => n646, A4 => n647, ZN 
                           => n637);
   U922 : OAI221_X1 port map( B1 => n618, B2 => n5113, C1 => n619, C2 => n5109,
                           A => n620, ZN => n617);
   U923 : AOI22_X1 port map( A1 => n5105, A2 => n4407, B1 => n5099, B2 => n4311
                           , ZN => n620);
   U924 : NOR4_X1 port map( A1 => n621, A2 => n622, A3 => n623, A4 => n624, ZN 
                           => n619);
   U925 : NOR4_X1 port map( A1 => n625, A2 => n626, A3 => n627, A4 => n628, ZN 
                           => n618);
   U926 : OAI221_X1 port map( B1 => n599, B2 => n5113, C1 => n600, C2 => n5109,
                           A => n601, ZN => n598);
   U927 : AOI22_X1 port map( A1 => n5105, A2 => n4408, B1 => n5099, B2 => n4312
                           , ZN => n601);
   U928 : NOR4_X1 port map( A1 => n602, A2 => n603, A3 => n604, A4 => n605, ZN 
                           => n600);
   U929 : NOR4_X1 port map( A1 => n606, A2 => n607, A3 => n608, A4 => n609, ZN 
                           => n599);
   U930 : OAI221_X1 port map( B1 => n580, B2 => n5113, C1 => n581, C2 => n5109,
                           A => n582, ZN => n579);
   U931 : AOI22_X1 port map( A1 => n5105, A2 => n4409, B1 => n5099, B2 => n4313
                           , ZN => n582);
   U932 : NOR4_X1 port map( A1 => n583, A2 => n584, A3 => n585, A4 => n586, ZN 
                           => n581);
   U933 : NOR4_X1 port map( A1 => n587, A2 => n588, A3 => n589, A4 => n590, ZN 
                           => n580);
   U934 : OAI221_X1 port map( B1 => n561, B2 => n5113, C1 => n562, C2 => n5109,
                           A => n563, ZN => n560);
   U935 : AOI22_X1 port map( A1 => n5105, A2 => n4410, B1 => n5099, B2 => n4314
                           , ZN => n563);
   U936 : NOR4_X1 port map( A1 => n564, A2 => n565, A3 => n566, A4 => n567, ZN 
                           => n562);
   U937 : NOR4_X1 port map( A1 => n568, A2 => n569, A3 => n570, A4 => n571, ZN 
                           => n561);
   U938 : OAI221_X1 port map( B1 => n542, B2 => n5114, C1 => n543, C2 => n5110,
                           A => n544, ZN => n541);
   U939 : AOI22_X1 port map( A1 => n5106, A2 => n4411, B1 => n5099, B2 => n4315
                           , ZN => n544);
   U940 : NOR4_X1 port map( A1 => n545, A2 => n546, A3 => n547, A4 => n548, ZN 
                           => n543);
   U941 : NOR4_X1 port map( A1 => n549, A2 => n550, A3 => n551, A4 => n552, ZN 
                           => n542);
   U942 : OAI221_X1 port map( B1 => n523, B2 => n5114, C1 => n524, C2 => n5110,
                           A => n525, ZN => n522);
   U943 : AOI22_X1 port map( A1 => n5106, A2 => n4412, B1 => n5099, B2 => n4316
                           , ZN => n525);
   U944 : NOR4_X1 port map( A1 => n526, A2 => n527, A3 => n528, A4 => n529, ZN 
                           => n524);
   U945 : NOR4_X1 port map( A1 => n530, A2 => n531, A3 => n532, A4 => n533, ZN 
                           => n523);
   U946 : OAI221_X1 port map( B1 => n504, B2 => n5114, C1 => n505, C2 => n5110,
                           A => n506, ZN => n503);
   U947 : AOI22_X1 port map( A1 => n5106, A2 => n4413, B1 => n5099, B2 => n4317
                           , ZN => n506);
   U948 : NOR4_X1 port map( A1 => n507, A2 => n508, A3 => n509, A4 => n510, ZN 
                           => n505);
   U949 : NOR4_X1 port map( A1 => n511, A2 => n512, A3 => n513, A4 => n514, ZN 
                           => n504);
   U950 : OAI221_X1 port map( B1 => n485, B2 => n5114, C1 => n486, C2 => n5110,
                           A => n487, ZN => n484);
   U951 : AOI22_X1 port map( A1 => n5106, A2 => n4414, B1 => n5099, B2 => n4318
                           , ZN => n487);
   U952 : NOR4_X1 port map( A1 => n488, A2 => n489, A3 => n490, A4 => n491, ZN 
                           => n486);
   U953 : NOR4_X1 port map( A1 => n492, A2 => n493, A3 => n494, A4 => n495, ZN 
                           => n485);
   U954 : OAI221_X1 port map( B1 => n466, B2 => n5114, C1 => n467, C2 => n5110,
                           A => n468, ZN => n465);
   U955 : AOI22_X1 port map( A1 => n5106, A2 => n4415, B1 => n5099, B2 => n4319
                           , ZN => n468);
   U956 : NOR4_X1 port map( A1 => n469, A2 => n470, A3 => n471, A4 => n472, ZN 
                           => n467);
   U957 : NOR4_X1 port map( A1 => n473, A2 => n474, A3 => n475, A4 => n476, ZN 
                           => n466);
   U958 : OAI221_X1 port map( B1 => n447, B2 => n5114, C1 => n448, C2 => n5110,
                           A => n449, ZN => n446);
   U959 : AOI22_X1 port map( A1 => n5106, A2 => n4416, B1 => n5099, B2 => n4320
                           , ZN => n449);
   U960 : NOR4_X1 port map( A1 => n450, A2 => n451, A3 => n452, A4 => n453, ZN 
                           => n448);
   U961 : NOR4_X1 port map( A1 => n454, A2 => n455, A3 => n456, A4 => n457, ZN 
                           => n447);
   U962 : INV_X1 port map( A => n1002, ZN => n5140);
   U963 : NOR3_X1 port map( A1 => n5150, A2 => n5149, A3 => n5144, ZN => n1003)
                           ;
   U964 : NOR3_X1 port map( A1 => n5137, A2 => n5136, A3 => n5131, ZN => n2665)
                           ;
   U965 : INV_X1 port map( A => n2674, ZN => n5130);
   U966 : INV_X1 port map( A => n1012, ZN => n5143);
   U967 : INV_X1 port map( A => n2675, ZN => n5129);
   U968 : INV_X1 port map( A => n1013, ZN => n5142);
   U969 : OAI221_X1 port map( B1 => n1066, B2 => n5034, C1 => n1067, C2 => 
                           n5030, A => n1068, ZN => n1065);
   U970 : AOI22_X1 port map( A1 => n5026, A2 => n4417, B1 => n5019, B2 => n4321
                           , ZN => n1068);
   U971 : NOR4_X1 port map( A1 => n1069, A2 => n1070, A3 => n1071, A4 => n1072,
                           ZN => n1067);
   U972 : NOR4_X1 port map( A1 => n1073, A2 => n1074, A3 => n1075, A4 => n1076,
                           ZN => n1066);
   U973 : OAI221_X1 port map( B1 => n1029, B2 => n5034, C1 => n1031, C2 => 
                           n5030, A => n1033, ZN => n1028);
   U974 : AOI22_X1 port map( A1 => n5026, A2 => n4418, B1 => n5019, B2 => n4322
                           , ZN => n1033);
   U975 : NOR4_X1 port map( A1 => n1036, A2 => n1037, A3 => n1038, A4 => n1039,
                           ZN => n1031);
   U976 : NOR4_X1 port map( A1 => n1040, A2 => n1041, A3 => n1042, A4 => n1043,
                           ZN => n1029);
   U977 : OAI221_X1 port map( B1 => n428, B2 => n5114, C1 => n429, C2 => n5110,
                           A => n430, ZN => n427);
   U978 : AOI22_X1 port map( A1 => n5106, A2 => n4417, B1 => n5099, B2 => n4321
                           , ZN => n430);
   U979 : NOR4_X1 port map( A1 => n431, A2 => n432, A3 => n433, A4 => n434, ZN 
                           => n429);
   U980 : NOR4_X1 port map( A1 => n435, A2 => n436, A3 => n437, A4 => n438, ZN 
                           => n428);
   U981 : OAI221_X1 port map( B1 => n391, B2 => n5114, C1 => n393, C2 => n5110,
                           A => n395, ZN => n390);
   U982 : AOI22_X1 port map( A1 => n5106, A2 => n4418, B1 => n5099, B2 => n4322
                           , ZN => n395);
   U983 : NOR4_X1 port map( A1 => n398, A2 => n399, A3 => n400, A4 => n401, ZN 
                           => n393);
   U984 : NOR4_X1 port map( A1 => n402, A2 => n403, A3 => n404, A4 => n405, ZN 
                           => n391);
   U985 : INV_X1 port map( A => n2676, ZN => n5133);
   U986 : INV_X1 port map( A => n2677, ZN => n5132);
   U987 : INV_X1 port map( A => n1014, ZN => n5146);
   U988 : INV_X1 port map( A => n1015, ZN => n5145);
   U989 : INV_X1 port map( A => n2678, ZN => n5134);
   U990 : INV_X1 port map( A => n1016, ZN => n5147);
   U991 : INV_X1 port map( A => n1017, ZN => n5148);
   U992 : INV_X1 port map( A => n2679, ZN => n5135);
   U993 : AND2_X1 port map( A1 => n2663, A2 => n2677, ZN => n1047);
   U994 : AND2_X1 port map( A1 => n2663, A2 => n2676, ZN => n1049);
   U995 : AND2_X1 port map( A1 => n1001, A2 => n1003, ZN => n396);
   U996 : AND2_X1 port map( A1 => n2663, A2 => n2665, ZN => n1034);
   U997 : AND2_X1 port map( A1 => n1001, A2 => n1002, ZN => n397);
   U998 : AND2_X1 port map( A1 => n2663, A2 => n2664, ZN => n1035);
   U999 : AND2_X1 port map( A1 => n1001, A2 => n1015, ZN => n409);
   U1000 : AND2_X1 port map( A1 => n1001, A2 => n1014, ZN => n411);
   U1001 : AOI222_X1 port map( A1 => n4972, A2 => n4419, B1 => n4969, B2 => 
                           n4259, C1 => n4965, C2 => n4195, ZN => n2683);
   U1002 : AOI222_X1 port map( A1 => n4972, A2 => n4420, B1 => n4969, B2 => 
                           n4260, C1 => n4965, C2 => n4196, ZN => n2654);
   U1003 : AOI222_X1 port map( A1 => n4972, A2 => n4421, B1 => n4969, B2 => 
                           n4261, C1 => n4965, C2 => n4197, ZN => n2635);
   U1004 : AOI222_X1 port map( A1 => n4972, A2 => n4422, B1 => n4969, B2 => 
                           n4262, C1 => n4965, C2 => n4198, ZN => n2616);
   U1005 : AOI222_X1 port map( A1 => n4972, A2 => n4423, B1 => n4969, B2 => 
                           n4263, C1 => n4965, C2 => n4199, ZN => n2597);
   U1006 : AOI222_X1 port map( A1 => n4972, A2 => n4424, B1 => n4969, B2 => 
                           n4264, C1 => n4965, C2 => n4200, ZN => n2578);
   U1007 : AOI222_X1 port map( A1 => n4972, A2 => n4425, B1 => n4969, B2 => 
                           n4265, C1 => n4965, C2 => n4201, ZN => n2559);
   U1008 : AOI222_X1 port map( A1 => n4972, A2 => n4426, B1 => n4969, B2 => 
                           n4266, C1 => n4965, C2 => n4202, ZN => n2540);
   U1009 : AND2_X1 port map( A1 => n2678, A2 => n2682, ZN => n1059);
   U1010 : AOI222_X1 port map( A1 => n4972, A2 => n4427, B1 => n4968, B2 => 
                           n4267, C1 => n4964, C2 => n4203, ZN => n2521);
   U1011 : AOI222_X1 port map( A1 => n4972, A2 => n4428, B1 => n4968, B2 => 
                           n4268, C1 => n4964, C2 => n4204, ZN => n2502);
   U1012 : AOI222_X1 port map( A1 => n4972, A2 => n4429, B1 => n4968, B2 => 
                           n4269, C1 => n4964, C2 => n4205, ZN => n2483);
   U1013 : AOI222_X1 port map( A1 => n4972, A2 => n4430, B1 => n4968, B2 => 
                           n4270, C1 => n4964, C2 => n4206, ZN => n2464);
   U1014 : AOI222_X1 port map( A1 => n4973, A2 => n4431, B1 => n4968, B2 => 
                           n4271, C1 => n4964, C2 => n4207, ZN => n2445);
   U1015 : AOI222_X1 port map( A1 => n4973, A2 => n4432, B1 => n4968, B2 => 
                           n4272, C1 => n4964, C2 => n4208, ZN => n2426);
   U1016 : AOI222_X1 port map( A1 => n4973, A2 => n4433, B1 => n4968, B2 => 
                           n4273, C1 => n4964, C2 => n4209, ZN => n2407);
   U1017 : AOI222_X1 port map( A1 => n4973, A2 => n4434, B1 => n4968, B2 => 
                           n4274, C1 => n4964, C2 => n4210, ZN => n2388);
   U1018 : AOI222_X1 port map( A1 => n4973, A2 => n4435, B1 => n4968, B2 => 
                           n4275, C1 => n4964, C2 => n4211, ZN => n2369);
   U1019 : AOI222_X1 port map( A1 => n4973, A2 => n4436, B1 => n4968, B2 => 
                           n4276, C1 => n4964, C2 => n4212, ZN => n2350);
   U1020 : AOI222_X1 port map( A1 => n4973, A2 => n4437, B1 => n4968, B2 => 
                           n4277, C1 => n4964, C2 => n4213, ZN => n2331);
   U1021 : AOI222_X1 port map( A1 => n4973, A2 => n4438, B1 => n4968, B2 => 
                           n4278, C1 => n4964, C2 => n4214, ZN => n1288);
   U1022 : AOI222_X1 port map( A1 => n4973, A2 => n4439, B1 => n4967, B2 => 
                           n4279, C1 => n4963, C2 => n4215, ZN => n1269);
   U1023 : AOI222_X1 port map( A1 => n4973, A2 => n4440, B1 => n4967, B2 => 
                           n4280, C1 => n4963, C2 => n4216, ZN => n1250);
   U1024 : AOI222_X1 port map( A1 => n4973, A2 => n4441, B1 => n4967, B2 => 
                           n4281, C1 => n4963, C2 => n4217, ZN => n1231);
   U1025 : AOI222_X1 port map( A1 => n4973, A2 => n4442, B1 => n4967, B2 => 
                           n4282, C1 => n4963, C2 => n4218, ZN => n1212);
   U1026 : AOI222_X1 port map( A1 => n4974, A2 => n4443, B1 => n4967, B2 => 
                           n4283, C1 => n4963, C2 => n4219, ZN => n1193);
   U1027 : AOI222_X1 port map( A1 => n4974, A2 => n4444, B1 => n4967, B2 => 
                           n4284, C1 => n4963, C2 => n4220, ZN => n1174);
   U1028 : AOI222_X1 port map( A1 => n4974, A2 => n4445, B1 => n4967, B2 => 
                           n4285, C1 => n4963, C2 => n4221, ZN => n1155);
   U1029 : AOI222_X1 port map( A1 => n4974, A2 => n4446, B1 => n4967, B2 => 
                           n4286, C1 => n4963, C2 => n4222, ZN => n1136);
   U1030 : AOI222_X1 port map( A1 => n4974, A2 => n4447, B1 => n4967, B2 => 
                           n4287, C1 => n4963, C2 => n4223, ZN => n1117);
   U1031 : AOI222_X1 port map( A1 => n4974, A2 => n4448, B1 => n4967, B2 => 
                           n4288, C1 => n4963, C2 => n4224, ZN => n1098);
   U1032 : AOI222_X1 port map( A1 => n4974, A2 => n4449, B1 => n4967, B2 => 
                           n4289, C1 => n4963, C2 => n4225, ZN => n1079);
   U1033 : AOI222_X1 port map( A1 => n4974, A2 => n4450, B1 => n4967, B2 => 
                           n4290, C1 => n4963, C2 => n4226, ZN => n1057);
   U1034 : AND2_X1 port map( A1 => n2663, A2 => n2678, ZN => n1054);
   U1035 : AOI22_X1 port map( A1 => n4988, A2 => n4451, B1 => n4985, B2 => 
                           n4323, ZN => n2681);
   U1036 : AOI22_X1 port map( A1 => n4988, A2 => n4452, B1 => n4985, B2 => 
                           n4324, ZN => n2653);
   U1037 : AOI22_X1 port map( A1 => n4988, A2 => n4453, B1 => n4985, B2 => 
                           n4325, ZN => n2634);
   U1038 : AOI22_X1 port map( A1 => n4988, A2 => n4454, B1 => n4985, B2 => 
                           n4326, ZN => n2615);
   U1039 : AOI22_X1 port map( A1 => n4988, A2 => n4455, B1 => n4985, B2 => 
                           n4327, ZN => n2596);
   U1040 : AOI22_X1 port map( A1 => n4988, A2 => n4456, B1 => n4985, B2 => 
                           n4328, ZN => n2577);
   U1041 : AOI22_X1 port map( A1 => n4988, A2 => n4457, B1 => n4985, B2 => 
                           n4329, ZN => n2558);
   U1042 : AOI22_X1 port map( A1 => n4988, A2 => n4458, B1 => n4985, B2 => 
                           n4330, ZN => n2539);
   U1043 : AND2_X1 port map( A1 => n1002, A2 => n1020, ZN => n415);
   U1044 : AOI22_X1 port map( A1 => n5070, A2 => n4475, B1 => n5063, B2 => 
                           n4347, ZN => n554);
   U1045 : AOI22_X1 port map( A1 => n5070, A2 => n4476, B1 => n5063, B2 => 
                           n4348, ZN => n535);
   U1046 : AOI22_X1 port map( A1 => n5070, A2 => n4477, B1 => n5063, B2 => 
                           n4349, ZN => n516);
   U1047 : AOI22_X1 port map( A1 => n5070, A2 => n4478, B1 => n5063, B2 => 
                           n4350, ZN => n497);
   U1048 : AOI22_X1 port map( A1 => n5070, A2 => n4479, B1 => n5063, B2 => 
                           n4351, ZN => n478);
   U1049 : AOI22_X1 port map( A1 => n5070, A2 => n4480, B1 => n5063, B2 => 
                           n4352, ZN => n459);
   U1050 : AOI22_X1 port map( A1 => n5070, A2 => n4481, B1 => n5063, B2 => 
                           n4353, ZN => n440);
   U1051 : AOI22_X1 port map( A1 => n5070, A2 => n4482, B1 => n5063, B2 => 
                           n4354, ZN => n414);
   U1052 : AND2_X1 port map( A1 => n2664, A2 => n2682, ZN => n1053);
   U1053 : AOI22_X1 port map( A1 => n4990, A2 => n4475, B1 => n4983, B2 => 
                           n4347, ZN => n1192);
   U1054 : AOI22_X1 port map( A1 => n4990, A2 => n4476, B1 => n4983, B2 => 
                           n4348, ZN => n1173);
   U1055 : AOI22_X1 port map( A1 => n4990, A2 => n4477, B1 => n4983, B2 => 
                           n4349, ZN => n1154);
   U1056 : AOI22_X1 port map( A1 => n4990, A2 => n4478, B1 => n4983, B2 => 
                           n4350, ZN => n1135);
   U1057 : AOI22_X1 port map( A1 => n4990, A2 => n4479, B1 => n4983, B2 => 
                           n4351, ZN => n1116);
   U1058 : AOI22_X1 port map( A1 => n4990, A2 => n4480, B1 => n4983, B2 => 
                           n4352, ZN => n1097);
   U1059 : AOI22_X1 port map( A1 => n4990, A2 => n4481, B1 => n4983, B2 => 
                           n4353, ZN => n1078);
   U1060 : AOI22_X1 port map( A1 => n4990, A2 => n4482, B1 => n4983, B2 => 
                           n4354, ZN => n1052);
   U1061 : AOI22_X1 port map( A1 => n4988, A2 => n4459, B1 => n4984, B2 => 
                           n4331, ZN => n2520);
   U1062 : AOI22_X1 port map( A1 => n4988, A2 => n4460, B1 => n4984, B2 => 
                           n4332, ZN => n2501);
   U1063 : AOI22_X1 port map( A1 => n4988, A2 => n4461, B1 => n4984, B2 => 
                           n4333, ZN => n2482);
   U1064 : AOI22_X1 port map( A1 => n4988, A2 => n4462, B1 => n4984, B2 => 
                           n4334, ZN => n2463);
   U1065 : AOI22_X1 port map( A1 => n4989, A2 => n4463, B1 => n4984, B2 => 
                           n4335, ZN => n2444);
   U1066 : AOI22_X1 port map( A1 => n4989, A2 => n4464, B1 => n4984, B2 => 
                           n4336, ZN => n2425);
   U1067 : AOI22_X1 port map( A1 => n4989, A2 => n4465, B1 => n4984, B2 => 
                           n4337, ZN => n2406);
   U1068 : AOI22_X1 port map( A1 => n4989, A2 => n4466, B1 => n4984, B2 => 
                           n4338, ZN => n2387);
   U1069 : AOI22_X1 port map( A1 => n4989, A2 => n4467, B1 => n4984, B2 => 
                           n4339, ZN => n2368);
   U1070 : AOI22_X1 port map( A1 => n4989, A2 => n4468, B1 => n4984, B2 => 
                           n4340, ZN => n2349);
   U1071 : AOI22_X1 port map( A1 => n4989, A2 => n4469, B1 => n4984, B2 => 
                           n4341, ZN => n2330);
   U1072 : AOI22_X1 port map( A1 => n4989, A2 => n4470, B1 => n4984, B2 => 
                           n4342, ZN => n1287);
   U1073 : AOI22_X1 port map( A1 => n4989, A2 => n4471, B1 => n4983, B2 => 
                           n4343, ZN => n1268);
   U1074 : AOI22_X1 port map( A1 => n4989, A2 => n4472, B1 => n4983, B2 => 
                           n4344, ZN => n1249);
   U1075 : AOI22_X1 port map( A1 => n4989, A2 => n4473, B1 => n4983, B2 => 
                           n4345, ZN => n1230);
   U1076 : AOI22_X1 port map( A1 => n4989, A2 => n4474, B1 => n4983, B2 => 
                           n4346, ZN => n1211);
   U1077 : AOI22_X1 port map( A1 => n5068, A2 => n4451, B1 => n5065, B2 => 
                           n4323, ZN => n1019);
   U1078 : AOI22_X1 port map( A1 => n5068, A2 => n4452, B1 => n5065, B2 => 
                           n4324, ZN => n991);
   U1079 : AOI22_X1 port map( A1 => n5068, A2 => n4453, B1 => n5065, B2 => 
                           n4325, ZN => n972);
   U1080 : AOI22_X1 port map( A1 => n5068, A2 => n4454, B1 => n5065, B2 => 
                           n4326, ZN => n953);
   U1081 : AOI22_X1 port map( A1 => n5068, A2 => n4455, B1 => n5065, B2 => 
                           n4327, ZN => n934);
   U1082 : AOI22_X1 port map( A1 => n5068, A2 => n4456, B1 => n5065, B2 => 
                           n4328, ZN => n915);
   U1083 : AOI22_X1 port map( A1 => n5068, A2 => n4457, B1 => n5065, B2 => 
                           n4329, ZN => n896);
   U1084 : AOI22_X1 port map( A1 => n5068, A2 => n4458, B1 => n5065, B2 => 
                           n4330, ZN => n877);
   U1085 : AOI22_X1 port map( A1 => n5068, A2 => n4459, B1 => n5064, B2 => 
                           n4331, ZN => n858);
   U1086 : AOI22_X1 port map( A1 => n5068, A2 => n4460, B1 => n5064, B2 => 
                           n4332, ZN => n839);
   U1087 : AOI22_X1 port map( A1 => n5068, A2 => n4461, B1 => n5064, B2 => 
                           n4333, ZN => n820);
   U1088 : AOI22_X1 port map( A1 => n5068, A2 => n4462, B1 => n5064, B2 => 
                           n4334, ZN => n801);
   U1089 : AOI22_X1 port map( A1 => n5069, A2 => n4463, B1 => n5064, B2 => 
                           n4335, ZN => n782);
   U1090 : AOI22_X1 port map( A1 => n5069, A2 => n4464, B1 => n5064, B2 => 
                           n4336, ZN => n763);
   U1091 : AOI22_X1 port map( A1 => n5069, A2 => n4465, B1 => n5064, B2 => 
                           n4337, ZN => n744);
   U1092 : AOI22_X1 port map( A1 => n5069, A2 => n4466, B1 => n5064, B2 => 
                           n4338, ZN => n725);
   U1093 : AOI22_X1 port map( A1 => n5069, A2 => n4467, B1 => n5064, B2 => 
                           n4339, ZN => n706);
   U1094 : AOI22_X1 port map( A1 => n5069, A2 => n4468, B1 => n5064, B2 => 
                           n4340, ZN => n687);
   U1095 : AOI22_X1 port map( A1 => n5069, A2 => n4469, B1 => n5064, B2 => 
                           n4341, ZN => n668);
   U1096 : AOI22_X1 port map( A1 => n5069, A2 => n4470, B1 => n5064, B2 => 
                           n4342, ZN => n649);
   U1097 : AOI22_X1 port map( A1 => n5069, A2 => n4471, B1 => n5063, B2 => 
                           n4343, ZN => n630);
   U1098 : AOI22_X1 port map( A1 => n5069, A2 => n4472, B1 => n5063, B2 => 
                           n4344, ZN => n611);
   U1099 : AOI22_X1 port map( A1 => n5069, A2 => n4473, B1 => n5063, B2 => 
                           n4345, ZN => n592);
   U1100 : AOI22_X1 port map( A1 => n5069, A2 => n4474, B1 => n5063, B2 => 
                           n4346, ZN => n573);
   U1101 : AND2_X1 port map( A1 => n2676, A2 => n2682, ZN => n1058);
   U1102 : AOI222_X1 port map( A1 => n5052, A2 => n4419, B1 => n5049, B2 => 
                           n4259, C1 => n5045, C2 => n4195, ZN => n1021);
   U1103 : AOI222_X1 port map( A1 => n5052, A2 => n4420, B1 => n5049, B2 => 
                           n4260, C1 => n5045, C2 => n4196, ZN => n992);
   U1104 : AOI222_X1 port map( A1 => n5052, A2 => n4421, B1 => n5049, B2 => 
                           n4261, C1 => n5045, C2 => n4197, ZN => n973);
   U1105 : AOI222_X1 port map( A1 => n5052, A2 => n4422, B1 => n5049, B2 => 
                           n4262, C1 => n5045, C2 => n4198, ZN => n954);
   U1106 : AOI222_X1 port map( A1 => n5052, A2 => n4423, B1 => n5049, B2 => 
                           n4263, C1 => n5045, C2 => n4199, ZN => n935);
   U1107 : AOI222_X1 port map( A1 => n5052, A2 => n4424, B1 => n5049, B2 => 
                           n4264, C1 => n5045, C2 => n4200, ZN => n916);
   U1108 : AOI222_X1 port map( A1 => n5052, A2 => n4425, B1 => n5049, B2 => 
                           n4265, C1 => n5045, C2 => n4201, ZN => n897);
   U1109 : AOI222_X1 port map( A1 => n5052, A2 => n4426, B1 => n5049, B2 => 
                           n4266, C1 => n5045, C2 => n4202, ZN => n878);
   U1110 : AND2_X1 port map( A1 => n1016, A2 => n1020, ZN => n421);
   U1111 : AOI222_X1 port map( A1 => n5052, A2 => n4427, B1 => n5048, B2 => 
                           n4267, C1 => n5044, C2 => n4203, ZN => n859);
   U1112 : AOI222_X1 port map( A1 => n5052, A2 => n4428, B1 => n5048, B2 => 
                           n4268, C1 => n5044, C2 => n4204, ZN => n840);
   U1113 : AOI222_X1 port map( A1 => n5052, A2 => n4429, B1 => n5048, B2 => 
                           n4269, C1 => n5044, C2 => n4205, ZN => n821);
   U1114 : AOI222_X1 port map( A1 => n5052, A2 => n4430, B1 => n5048, B2 => 
                           n4270, C1 => n5044, C2 => n4206, ZN => n802);
   U1115 : AOI222_X1 port map( A1 => n5053, A2 => n4431, B1 => n5048, B2 => 
                           n4271, C1 => n5044, C2 => n4207, ZN => n783);
   U1116 : AOI222_X1 port map( A1 => n5053, A2 => n4432, B1 => n5048, B2 => 
                           n4272, C1 => n5044, C2 => n4208, ZN => n764);
   U1117 : AOI222_X1 port map( A1 => n5053, A2 => n4433, B1 => n5048, B2 => 
                           n4273, C1 => n5044, C2 => n4209, ZN => n745);
   U1118 : AOI222_X1 port map( A1 => n5053, A2 => n4434, B1 => n5048, B2 => 
                           n4274, C1 => n5044, C2 => n4210, ZN => n726);
   U1119 : AOI222_X1 port map( A1 => n5053, A2 => n4435, B1 => n5048, B2 => 
                           n4275, C1 => n5044, C2 => n4211, ZN => n707);
   U1120 : AOI222_X1 port map( A1 => n5053, A2 => n4436, B1 => n5048, B2 => 
                           n4276, C1 => n5044, C2 => n4212, ZN => n688);
   U1121 : AOI222_X1 port map( A1 => n5053, A2 => n4437, B1 => n5048, B2 => 
                           n4277, C1 => n5044, C2 => n4213, ZN => n669);
   U1122 : AOI222_X1 port map( A1 => n5053, A2 => n4438, B1 => n5048, B2 => 
                           n4278, C1 => n5044, C2 => n4214, ZN => n650);
   U1123 : AOI222_X1 port map( A1 => n5053, A2 => n4439, B1 => n5047, B2 => 
                           n4279, C1 => n5043, C2 => n4215, ZN => n631);
   U1124 : AOI222_X1 port map( A1 => n5053, A2 => n4440, B1 => n5047, B2 => 
                           n4280, C1 => n5043, C2 => n4216, ZN => n612);
   U1125 : AOI222_X1 port map( A1 => n5053, A2 => n4441, B1 => n5047, B2 => 
                           n4281, C1 => n5043, C2 => n4217, ZN => n593);
   U1126 : AOI222_X1 port map( A1 => n5053, A2 => n4442, B1 => n5047, B2 => 
                           n4282, C1 => n5043, C2 => n4218, ZN => n574);
   U1127 : AOI222_X1 port map( A1 => n5054, A2 => n4443, B1 => n5047, B2 => 
                           n4283, C1 => n5043, C2 => n4219, ZN => n555);
   U1128 : AOI222_X1 port map( A1 => n5054, A2 => n4444, B1 => n5047, B2 => 
                           n4284, C1 => n5043, C2 => n4220, ZN => n536);
   U1129 : AOI222_X1 port map( A1 => n5054, A2 => n4445, B1 => n5047, B2 => 
                           n4285, C1 => n5043, C2 => n4221, ZN => n517);
   U1130 : AOI222_X1 port map( A1 => n5054, A2 => n4446, B1 => n5047, B2 => 
                           n4286, C1 => n5043, C2 => n4222, ZN => n498);
   U1131 : AOI222_X1 port map( A1 => n5054, A2 => n4447, B1 => n5047, B2 => 
                           n4287, C1 => n5043, C2 => n4223, ZN => n479);
   U1132 : AOI222_X1 port map( A1 => n5054, A2 => n4448, B1 => n5047, B2 => 
                           n4288, C1 => n5043, C2 => n4224, ZN => n460);
   U1133 : AOI222_X1 port map( A1 => n5054, A2 => n4449, B1 => n5047, B2 => 
                           n4289, C1 => n5043, C2 => n4225, ZN => n441);
   U1134 : AOI222_X1 port map( A1 => n5054, A2 => n4450, B1 => n5047, B2 => 
                           n4290, C1 => n5043, C2 => n4226, ZN => n419);
   U1135 : AND2_X1 port map( A1 => n1001, A2 => n1016, ZN => n416);
   U1136 : AND2_X1 port map( A1 => n1014, A2 => n1020, ZN => n420);
   U1137 : NOR2_X1 port map( A1 => n5152, A2 => n5151, ZN => n1020);
   U1138 : AND2_X1 port map( A1 => n1017, A2 => n1020, ZN => n422);
   U1139 : NOR2_X1 port map( A1 => n5139, A2 => n5138, ZN => n2682);
   U1140 : AND2_X1 port map( A1 => n2679, A2 => n2682, ZN => n1060);
   U1141 : AND2_X1 port map( A1 => n1001, A2 => n1017, ZN => n410);
   U1142 : AND2_X1 port map( A1 => n2663, A2 => n2679, ZN => n1048);
   U1143 : NAND2_X1 port map( A1 => n1001, A2 => n1012, ZN => n406);
   U1144 : NAND2_X1 port map( A1 => n2663, A2 => n2674, ZN => n1044);
   U1145 : NAND2_X1 port map( A1 => n1013, A2 => n1020, ZN => n412);
   U1146 : NAND2_X1 port map( A1 => n2675, A2 => n2682, ZN => n1050);
   U1147 : NAND2_X1 port map( A1 => n1001, A2 => n1013, ZN => n407);
   U1148 : NAND2_X1 port map( A1 => n2663, A2 => n2675, ZN => n1045);
   U1149 : NAND2_X1 port map( A1 => n2677, A2 => n2682, ZN => n1055);
   U1150 : NAND2_X1 port map( A1 => n1012, A2 => n1020, ZN => n418);
   U1151 : NAND2_X1 port map( A1 => n2674, A2 => n2682, ZN => n1056);
   U1152 : NAND2_X1 port map( A1 => n1015, A2 => n1020, ZN => n417);
   U1153 : NAND2_X1 port map( A1 => n5151, A2 => n5152, ZN => n394);
   U1154 : NAND2_X1 port map( A1 => n5138, A2 => n5139, ZN => n1032);
   U1155 : BUF_X1 port map( A => n5111, Z => n5114);
   U1156 : BUF_X1 port map( A => n5031, Z => n5034);
   U1157 : BUF_X1 port map( A => n5111, Z => n5112);
   U1158 : BUF_X1 port map( A => n5111, Z => n5113);
   U1159 : BUF_X1 port map( A => n5031, Z => n5032);
   U1160 : BUF_X1 port map( A => n5031, Z => n5033);
   U1161 : BUF_X1 port map( A => n5115, Z => n5116);
   U1162 : BUF_X1 port map( A => n5035, Z => n5036);
   U1163 : BUF_X1 port map( A => n5115, Z => n5117);
   U1164 : BUF_X1 port map( A => n5035, Z => n5037);
   U1165 : BUF_X1 port map( A => n5115, Z => n5118);
   U1166 : BUF_X1 port map( A => n5035, Z => n5038);
   U1167 : OAI22_X1 port map( A1 => n4960, A2 => n4620, B1 => n4070, B2 => 
                           n4956, ZN => n2298);
   U1168 : OAI22_X1 port map( A1 => n4960, A2 => n4623, B1 => n4071, B2 => 
                           n4956, ZN => n2299);
   U1169 : OAI22_X1 port map( A1 => n4960, A2 => n4626, B1 => n4072, B2 => 
                           n4956, ZN => n2300);
   U1170 : OAI22_X1 port map( A1 => n4960, A2 => n4629, B1 => n4073, B2 => 
                           n4956, ZN => n2301);
   U1171 : OAI22_X1 port map( A1 => n4960, A2 => n4632, B1 => n4074, B2 => 
                           n4956, ZN => n2302);
   U1172 : OAI22_X1 port map( A1 => n4960, A2 => n4635, B1 => n4075, B2 => 
                           n4956, ZN => n2303);
   U1173 : OAI22_X1 port map( A1 => n4962, A2 => n4704, B1 => n4098, B2 => 
                           n4958, ZN => n2326);
   U1174 : INV_X1 port map( A => DATAIN(3), ZN => n5156);
   U1175 : INV_X1 port map( A => DATAIN(4), ZN => n5157);
   U1176 : INV_X1 port map( A => DATAIN(5), ZN => n5158);
   U1177 : INV_X1 port map( A => DATAIN(6), ZN => n5159);
   U1178 : INV_X1 port map( A => DATAIN(7), ZN => n5160);
   U1179 : INV_X1 port map( A => DATAIN(8), ZN => n5161);
   U1180 : INV_X1 port map( A => DATAIN(31), ZN => n5184);
   U1181 : OAI22_X1 port map( A1 => n4960, A2 => n4611, B1 => n4067, B2 => 
                           n4956, ZN => n2295);
   U1182 : OAI22_X1 port map( A1 => n4960, A2 => n4614, B1 => n4068, B2 => 
                           n4956, ZN => n2296);
   U1183 : OAI22_X1 port map( A1 => n4960, A2 => n4617, B1 => n4069, B2 => 
                           n4956, ZN => n2297);
   U1184 : OAI22_X1 port map( A1 => n4960, A2 => n4641, B1 => n4077, B2 => 
                           n4956, ZN => n2305);
   U1185 : OAI22_X1 port map( A1 => n4960, A2 => n4644, B1 => n4078, B2 => 
                           n4956, ZN => n2306);
   U1186 : OAI22_X1 port map( A1 => n4961, A2 => n4647, B1 => n4079, B2 => 
                           n4957, ZN => n2307);
   U1187 : OAI22_X1 port map( A1 => n4961, A2 => n4650, B1 => n4080, B2 => 
                           n4957, ZN => n2308);
   U1188 : OAI22_X1 port map( A1 => n4961, A2 => n4653, B1 => n4081, B2 => 
                           n4957, ZN => n2309);
   U1189 : OAI22_X1 port map( A1 => n4961, A2 => n4656, B1 => n4082, B2 => 
                           n4957, ZN => n2310);
   U1190 : OAI22_X1 port map( A1 => n4961, A2 => n4659, B1 => n4083, B2 => 
                           n4957, ZN => n2311);
   U1191 : OAI22_X1 port map( A1 => n4961, A2 => n4662, B1 => n4084, B2 => 
                           n4957, ZN => n2312);
   U1192 : OAI22_X1 port map( A1 => n4961, A2 => n4665, B1 => n4085, B2 => 
                           n4957, ZN => n2313);
   U1193 : OAI22_X1 port map( A1 => n4961, A2 => n4668, B1 => n4086, B2 => 
                           n4957, ZN => n2314);
   U1194 : OAI22_X1 port map( A1 => n4961, A2 => n4671, B1 => n4087, B2 => 
                           n4957, ZN => n2315);
   U1195 : OAI22_X1 port map( A1 => n4961, A2 => n4674, B1 => n4088, B2 => 
                           n4957, ZN => n2316);
   U1196 : OAI22_X1 port map( A1 => n4961, A2 => n4677, B1 => n4089, B2 => 
                           n4957, ZN => n2317);
   U1197 : OAI22_X1 port map( A1 => n4961, A2 => n4680, B1 => n4090, B2 => 
                           n4957, ZN => n2318);
   U1198 : OAI22_X1 port map( A1 => n4961, A2 => n4683, B1 => n4091, B2 => 
                           n4958, ZN => n2319);
   U1199 : OAI22_X1 port map( A1 => n4962, A2 => n4686, B1 => n4092, B2 => 
                           n4958, ZN => n2320);
   U1200 : OAI22_X1 port map( A1 => n4962, A2 => n4689, B1 => n4093, B2 => 
                           n4958, ZN => n2321);
   U1201 : OAI22_X1 port map( A1 => n4962, A2 => n4692, B1 => n4094, B2 => 
                           n4958, ZN => n2322);
   U1202 : OAI22_X1 port map( A1 => n4962, A2 => n4695, B1 => n4095, B2 => 
                           n4958, ZN => n2323);
   U1203 : OAI22_X1 port map( A1 => n4962, A2 => n4698, B1 => n4096, B2 => 
                           n4958, ZN => n2324);
   U1204 : OAI22_X1 port map( A1 => n4962, A2 => n4701, B1 => n4097, B2 => 
                           n4958, ZN => n2325);
   U1205 : INV_X1 port map( A => DATAIN(0), ZN => n5153);
   U1206 : INV_X1 port map( A => DATAIN(1), ZN => n5154);
   U1207 : INV_X1 port map( A => DATAIN(2), ZN => n5155);
   U1208 : INV_X1 port map( A => DATAIN(10), ZN => n5163);
   U1209 : INV_X1 port map( A => DATAIN(11), ZN => n5164);
   U1210 : INV_X1 port map( A => DATAIN(12), ZN => n5165);
   U1211 : INV_X1 port map( A => DATAIN(13), ZN => n5166);
   U1212 : INV_X1 port map( A => DATAIN(14), ZN => n5167);
   U1213 : INV_X1 port map( A => DATAIN(15), ZN => n5168);
   U1214 : INV_X1 port map( A => DATAIN(16), ZN => n5169);
   U1215 : INV_X1 port map( A => DATAIN(17), ZN => n5170);
   U1216 : INV_X1 port map( A => DATAIN(18), ZN => n5171);
   U1217 : INV_X1 port map( A => DATAIN(19), ZN => n5172);
   U1218 : INV_X1 port map( A => DATAIN(20), ZN => n5173);
   U1219 : INV_X1 port map( A => DATAIN(21), ZN => n5174);
   U1220 : INV_X1 port map( A => DATAIN(22), ZN => n5175);
   U1221 : INV_X1 port map( A => DATAIN(23), ZN => n5176);
   U1222 : INV_X1 port map( A => DATAIN(24), ZN => n5177);
   U1223 : INV_X1 port map( A => DATAIN(25), ZN => n5178);
   U1224 : INV_X1 port map( A => DATAIN(26), ZN => n5179);
   U1225 : INV_X1 port map( A => DATAIN(27), ZN => n5180);
   U1226 : INV_X1 port map( A => DATAIN(28), ZN => n5181);
   U1227 : INV_X1 port map( A => DATAIN(29), ZN => n5182);
   U1228 : INV_X1 port map( A => DATAIN(30), ZN => n5183);
   U1229 : OAI22_X1 port map( A1 => n4621, A2 => n4760, B1 => n3270, B2 => 
                           n4756, ZN => n1498);
   U1230 : OAI22_X1 port map( A1 => n4624, A2 => n4760, B1 => n3271, B2 => 
                           n4756, ZN => n1499);
   U1231 : OAI22_X1 port map( A1 => n4627, A2 => n4760, B1 => n3272, B2 => 
                           n4756, ZN => n1500);
   U1232 : OAI22_X1 port map( A1 => n4630, A2 => n4760, B1 => n3273, B2 => 
                           n4756, ZN => n1501);
   U1233 : OAI22_X1 port map( A1 => n4633, A2 => n4760, B1 => n3274, B2 => 
                           n4756, ZN => n1502);
   U1234 : OAI22_X1 port map( A1 => n4636, A2 => n4760, B1 => n3275, B2 => 
                           n4756, ZN => n1503);
   U1235 : OAI22_X1 port map( A1 => n4705, A2 => n4762, B1 => n3298, B2 => 
                           n4758, ZN => n1526);
   U1236 : OAI22_X1 port map( A1 => n4621, A2 => n4808, B1 => n3462, B2 => 
                           n4804, ZN => n1690);
   U1237 : OAI22_X1 port map( A1 => n4624, A2 => n4808, B1 => n3463, B2 => 
                           n4804, ZN => n1691);
   U1238 : OAI22_X1 port map( A1 => n4627, A2 => n4808, B1 => n3464, B2 => 
                           n4804, ZN => n1692);
   U1239 : OAI22_X1 port map( A1 => n4630, A2 => n4808, B1 => n3465, B2 => 
                           n4804, ZN => n1693);
   U1240 : OAI22_X1 port map( A1 => n4633, A2 => n4808, B1 => n3466, B2 => 
                           n4804, ZN => n1694);
   U1241 : OAI22_X1 port map( A1 => n4636, A2 => n4808, B1 => n3467, B2 => 
                           n4804, ZN => n1695);
   U1242 : OAI22_X1 port map( A1 => n4705, A2 => n4810, B1 => n3490, B2 => 
                           n4806, ZN => n1718);
   U1243 : OAI22_X1 port map( A1 => n4620, A2 => n4864, B1 => n3686, B2 => 
                           n4860, ZN => n1914);
   U1244 : OAI22_X1 port map( A1 => n4623, A2 => n4864, B1 => n3687, B2 => 
                           n4860, ZN => n1915);
   U1245 : OAI22_X1 port map( A1 => n4626, A2 => n4864, B1 => n3688, B2 => 
                           n4860, ZN => n1916);
   U1246 : OAI22_X1 port map( A1 => n4629, A2 => n4864, B1 => n3689, B2 => 
                           n4860, ZN => n1917);
   U1247 : OAI22_X1 port map( A1 => n4632, A2 => n4864, B1 => n3690, B2 => 
                           n4860, ZN => n1918);
   U1248 : OAI22_X1 port map( A1 => n4635, A2 => n4864, B1 => n3691, B2 => 
                           n4860, ZN => n1919);
   U1249 : OAI22_X1 port map( A1 => n4704, A2 => n4866, B1 => n3714, B2 => 
                           n4862, ZN => n1942);
   U1250 : OAI22_X1 port map( A1 => n4620, A2 => n4888, B1 => n3782, B2 => 
                           n4884, ZN => n2010);
   U1251 : OAI22_X1 port map( A1 => n4623, A2 => n4888, B1 => n3783, B2 => 
                           n4884, ZN => n2011);
   U1252 : OAI22_X1 port map( A1 => n4626, A2 => n4888, B1 => n3784, B2 => 
                           n4884, ZN => n2012);
   U1253 : OAI22_X1 port map( A1 => n4629, A2 => n4888, B1 => n3785, B2 => 
                           n4884, ZN => n2013);
   U1254 : OAI22_X1 port map( A1 => n4632, A2 => n4888, B1 => n3786, B2 => 
                           n4884, ZN => n2014);
   U1255 : OAI22_X1 port map( A1 => n4635, A2 => n4888, B1 => n3787, B2 => 
                           n4884, ZN => n2015);
   U1256 : OAI22_X1 port map( A1 => n4704, A2 => n4890, B1 => n3810, B2 => 
                           n4886, ZN => n2038);
   U1257 : OAI22_X1 port map( A1 => n4620, A2 => n4896, B1 => n3814, B2 => 
                           n4892, ZN => n2042);
   U1258 : OAI22_X1 port map( A1 => n4623, A2 => n4896, B1 => n3815, B2 => 
                           n4892, ZN => n2043);
   U1259 : OAI22_X1 port map( A1 => n4626, A2 => n4896, B1 => n3816, B2 => 
                           n4892, ZN => n2044);
   U1260 : OAI22_X1 port map( A1 => n4629, A2 => n4896, B1 => n3817, B2 => 
                           n4892, ZN => n2045);
   U1261 : OAI22_X1 port map( A1 => n4632, A2 => n4896, B1 => n3818, B2 => 
                           n4892, ZN => n2046);
   U1262 : OAI22_X1 port map( A1 => n4635, A2 => n4896, B1 => n3819, B2 => 
                           n4892, ZN => n2047);
   U1263 : OAI22_X1 port map( A1 => n4704, A2 => n4898, B1 => n3842, B2 => 
                           n4894, ZN => n2070);
   U1264 : OAI22_X1 port map( A1 => n4620, A2 => n4920, B1 => n3910, B2 => 
                           n4916, ZN => n2138);
   U1265 : OAI22_X1 port map( A1 => n4623, A2 => n4920, B1 => n3911, B2 => 
                           n4916, ZN => n2139);
   U1266 : OAI22_X1 port map( A1 => n4626, A2 => n4920, B1 => n3912, B2 => 
                           n4916, ZN => n2140);
   U1267 : OAI22_X1 port map( A1 => n4629, A2 => n4920, B1 => n3913, B2 => 
                           n4916, ZN => n2141);
   U1268 : OAI22_X1 port map( A1 => n4632, A2 => n4920, B1 => n3914, B2 => 
                           n4916, ZN => n2142);
   U1269 : OAI22_X1 port map( A1 => n4635, A2 => n4920, B1 => n3915, B2 => 
                           n4916, ZN => n2143);
   U1270 : OAI22_X1 port map( A1 => n4704, A2 => n4922, B1 => n3938, B2 => 
                           n4918, ZN => n2166);
   U1271 : OAI22_X1 port map( A1 => n4620, A2 => n4928, B1 => n3942, B2 => 
                           n4924, ZN => n2170);
   U1272 : OAI22_X1 port map( A1 => n4623, A2 => n4928, B1 => n3943, B2 => 
                           n4924, ZN => n2171);
   U1273 : OAI22_X1 port map( A1 => n4626, A2 => n4928, B1 => n3944, B2 => 
                           n4924, ZN => n2172);
   U1274 : OAI22_X1 port map( A1 => n4629, A2 => n4928, B1 => n3945, B2 => 
                           n4924, ZN => n2173);
   U1275 : OAI22_X1 port map( A1 => n4632, A2 => n4928, B1 => n3946, B2 => 
                           n4924, ZN => n2174);
   U1276 : OAI22_X1 port map( A1 => n4635, A2 => n4928, B1 => n3947, B2 => 
                           n4924, ZN => n2175);
   U1277 : OAI22_X1 port map( A1 => n4704, A2 => n4930, B1 => n3970, B2 => 
                           n4926, ZN => n2198);
   U1278 : OAI22_X1 port map( A1 => n4620, A2 => n4952, B1 => n4038, B2 => 
                           n4948, ZN => n2266);
   U1279 : OAI22_X1 port map( A1 => n4623, A2 => n4952, B1 => n4039, B2 => 
                           n4948, ZN => n2267);
   U1280 : OAI22_X1 port map( A1 => n4626, A2 => n4952, B1 => n4040, B2 => 
                           n4948, ZN => n2268);
   U1281 : OAI22_X1 port map( A1 => n4629, A2 => n4952, B1 => n4041, B2 => 
                           n4948, ZN => n2269);
   U1282 : OAI22_X1 port map( A1 => n4632, A2 => n4952, B1 => n4042, B2 => 
                           n4948, ZN => n2270);
   U1283 : OAI22_X1 port map( A1 => n4635, A2 => n4952, B1 => n4043, B2 => 
                           n4948, ZN => n2271);
   U1284 : OAI22_X1 port map( A1 => n4704, A2 => n4954, B1 => n4066, B2 => 
                           n4950, ZN => n2294);
   U1285 : OAI22_X1 port map( A1 => n4620, A2 => n4872, B1 => n3718, B2 => 
                           n4868, ZN => n1946);
   U1286 : OAI22_X1 port map( A1 => n4623, A2 => n4872, B1 => n3719, B2 => 
                           n4868, ZN => n1947);
   U1287 : OAI22_X1 port map( A1 => n4626, A2 => n4872, B1 => n3720, B2 => 
                           n4868, ZN => n1948);
   U1288 : OAI22_X1 port map( A1 => n4629, A2 => n4872, B1 => n3721, B2 => 
                           n4868, ZN => n1949);
   U1289 : OAI22_X1 port map( A1 => n4632, A2 => n4872, B1 => n3722, B2 => 
                           n4868, ZN => n1950);
   U1290 : OAI22_X1 port map( A1 => n4635, A2 => n4872, B1 => n3723, B2 => 
                           n4868, ZN => n1951);
   U1291 : OAI22_X1 port map( A1 => n4704, A2 => n4874, B1 => n3746, B2 => 
                           n4870, ZN => n1974);
   U1292 : OAI22_X1 port map( A1 => n4620, A2 => n4880, B1 => n3750, B2 => 
                           n4876, ZN => n1978);
   U1293 : OAI22_X1 port map( A1 => n4623, A2 => n4880, B1 => n3751, B2 => 
                           n4876, ZN => n1979);
   U1294 : OAI22_X1 port map( A1 => n4626, A2 => n4880, B1 => n3752, B2 => 
                           n4876, ZN => n1980);
   U1295 : OAI22_X1 port map( A1 => n4629, A2 => n4880, B1 => n3753, B2 => 
                           n4876, ZN => n1981);
   U1296 : OAI22_X1 port map( A1 => n4632, A2 => n4880, B1 => n3754, B2 => 
                           n4876, ZN => n1982);
   U1297 : OAI22_X1 port map( A1 => n4635, A2 => n4880, B1 => n3755, B2 => 
                           n4876, ZN => n1983);
   U1298 : OAI22_X1 port map( A1 => n4704, A2 => n4882, B1 => n3778, B2 => 
                           n4878, ZN => n2006);
   U1299 : OAI22_X1 port map( A1 => n4620, A2 => n4904, B1 => n3846, B2 => 
                           n4900, ZN => n2074);
   U1300 : OAI22_X1 port map( A1 => n4623, A2 => n4904, B1 => n3847, B2 => 
                           n4900, ZN => n2075);
   U1301 : OAI22_X1 port map( A1 => n4626, A2 => n4904, B1 => n3848, B2 => 
                           n4900, ZN => n2076);
   U1302 : OAI22_X1 port map( A1 => n4629, A2 => n4904, B1 => n3849, B2 => 
                           n4900, ZN => n2077);
   U1303 : OAI22_X1 port map( A1 => n4632, A2 => n4904, B1 => n3850, B2 => 
                           n4900, ZN => n2078);
   U1304 : OAI22_X1 port map( A1 => n4635, A2 => n4904, B1 => n3851, B2 => 
                           n4900, ZN => n2079);
   U1305 : OAI22_X1 port map( A1 => n4704, A2 => n4906, B1 => n3874, B2 => 
                           n4902, ZN => n2102);
   U1306 : OAI22_X1 port map( A1 => n4620, A2 => n4912, B1 => n3878, B2 => 
                           n4908, ZN => n2106);
   U1307 : OAI22_X1 port map( A1 => n4623, A2 => n4912, B1 => n3879, B2 => 
                           n4908, ZN => n2107);
   U1308 : OAI22_X1 port map( A1 => n4626, A2 => n4912, B1 => n3880, B2 => 
                           n4908, ZN => n2108);
   U1309 : OAI22_X1 port map( A1 => n4629, A2 => n4912, B1 => n3881, B2 => 
                           n4908, ZN => n2109);
   U1310 : OAI22_X1 port map( A1 => n4632, A2 => n4912, B1 => n3882, B2 => 
                           n4908, ZN => n2110);
   U1311 : OAI22_X1 port map( A1 => n4635, A2 => n4912, B1 => n3883, B2 => 
                           n4908, ZN => n2111);
   U1312 : OAI22_X1 port map( A1 => n4704, A2 => n4914, B1 => n3906, B2 => 
                           n4910, ZN => n2134);
   U1313 : OAI22_X1 port map( A1 => n4620, A2 => n4936, B1 => n3974, B2 => 
                           n4932, ZN => n2202);
   U1314 : OAI22_X1 port map( A1 => n4623, A2 => n4936, B1 => n3975, B2 => 
                           n4932, ZN => n2203);
   U1315 : OAI22_X1 port map( A1 => n4626, A2 => n4936, B1 => n3976, B2 => 
                           n4932, ZN => n2204);
   U1316 : OAI22_X1 port map( A1 => n4629, A2 => n4936, B1 => n3977, B2 => 
                           n4932, ZN => n2205);
   U1317 : OAI22_X1 port map( A1 => n4632, A2 => n4936, B1 => n3978, B2 => 
                           n4932, ZN => n2206);
   U1318 : OAI22_X1 port map( A1 => n4635, A2 => n4936, B1 => n3979, B2 => 
                           n4932, ZN => n2207);
   U1319 : OAI22_X1 port map( A1 => n4704, A2 => n4938, B1 => n4002, B2 => 
                           n4934, ZN => n2230);
   U1320 : OAI22_X1 port map( A1 => n4620, A2 => n4944, B1 => n4006, B2 => 
                           n4940, ZN => n2234);
   U1321 : OAI22_X1 port map( A1 => n4623, A2 => n4944, B1 => n4007, B2 => 
                           n4940, ZN => n2235);
   U1322 : OAI22_X1 port map( A1 => n4626, A2 => n4944, B1 => n4008, B2 => 
                           n4940, ZN => n2236);
   U1323 : OAI22_X1 port map( A1 => n4629, A2 => n4944, B1 => n4009, B2 => 
                           n4940, ZN => n2237);
   U1324 : OAI22_X1 port map( A1 => n4632, A2 => n4944, B1 => n4010, B2 => 
                           n4940, ZN => n2238);
   U1325 : OAI22_X1 port map( A1 => n4635, A2 => n4944, B1 => n4011, B2 => 
                           n4940, ZN => n2239);
   U1326 : OAI22_X1 port map( A1 => n4704, A2 => n4946, B1 => n4034, B2 => 
                           n4942, ZN => n2262);
   U1327 : OAI22_X1 port map( A1 => n4621, A2 => n4824, B1 => n3526, B2 => 
                           n4820, ZN => n1754);
   U1328 : OAI22_X1 port map( A1 => n4624, A2 => n4824, B1 => n3527, B2 => 
                           n4820, ZN => n1755);
   U1329 : OAI22_X1 port map( A1 => n4627, A2 => n4824, B1 => n3528, B2 => 
                           n4820, ZN => n1756);
   U1330 : OAI22_X1 port map( A1 => n4630, A2 => n4824, B1 => n3529, B2 => 
                           n4820, ZN => n1757);
   U1331 : OAI22_X1 port map( A1 => n4633, A2 => n4824, B1 => n3530, B2 => 
                           n4820, ZN => n1758);
   U1332 : OAI22_X1 port map( A1 => n4636, A2 => n4824, B1 => n3531, B2 => 
                           n4820, ZN => n1759);
   U1333 : OAI22_X1 port map( A1 => n4705, A2 => n4826, B1 => n3554, B2 => 
                           n4822, ZN => n1782);
   U1334 : OAI22_X1 port map( A1 => n4621, A2 => n4856, B1 => n3654, B2 => 
                           n4852, ZN => n1882);
   U1335 : OAI22_X1 port map( A1 => n4624, A2 => n4856, B1 => n3655, B2 => 
                           n4852, ZN => n1883);
   U1336 : OAI22_X1 port map( A1 => n4627, A2 => n4856, B1 => n3656, B2 => 
                           n4852, ZN => n1884);
   U1337 : OAI22_X1 port map( A1 => n4630, A2 => n4856, B1 => n3657, B2 => 
                           n4852, ZN => n1885);
   U1338 : OAI22_X1 port map( A1 => n4633, A2 => n4856, B1 => n3658, B2 => 
                           n4852, ZN => n1886);
   U1339 : OAI22_X1 port map( A1 => n4636, A2 => n4856, B1 => n3659, B2 => 
                           n4852, ZN => n1887);
   U1340 : OAI22_X1 port map( A1 => n4705, A2 => n4858, B1 => n3682, B2 => 
                           n4854, ZN => n1910);
   U1341 : OAI22_X1 port map( A1 => n4621, A2 => n4840, B1 => n3590, B2 => 
                           n4836, ZN => n1818);
   U1342 : OAI22_X1 port map( A1 => n4624, A2 => n4840, B1 => n3591, B2 => 
                           n4836, ZN => n1819);
   U1343 : OAI22_X1 port map( A1 => n4627, A2 => n4840, B1 => n3592, B2 => 
                           n4836, ZN => n1820);
   U1344 : OAI22_X1 port map( A1 => n4630, A2 => n4840, B1 => n3593, B2 => 
                           n4836, ZN => n1821);
   U1345 : OAI22_X1 port map( A1 => n4633, A2 => n4840, B1 => n3594, B2 => 
                           n4836, ZN => n1822);
   U1346 : OAI22_X1 port map( A1 => n4636, A2 => n4840, B1 => n3595, B2 => 
                           n4836, ZN => n1823);
   U1347 : OAI22_X1 port map( A1 => n4705, A2 => n4842, B1 => n3618, B2 => 
                           n4838, ZN => n1846);
   U1348 : OAI22_X1 port map( A1 => n4621, A2 => n4848, B1 => n3622, B2 => 
                           n4844, ZN => n1850);
   U1349 : OAI22_X1 port map( A1 => n4624, A2 => n4848, B1 => n3623, B2 => 
                           n4844, ZN => n1851);
   U1350 : OAI22_X1 port map( A1 => n4627, A2 => n4848, B1 => n3624, B2 => 
                           n4844, ZN => n1852);
   U1351 : OAI22_X1 port map( A1 => n4630, A2 => n4848, B1 => n3625, B2 => 
                           n4844, ZN => n1853);
   U1352 : OAI22_X1 port map( A1 => n4633, A2 => n4848, B1 => n3626, B2 => 
                           n4844, ZN => n1854);
   U1353 : OAI22_X1 port map( A1 => n4636, A2 => n4848, B1 => n3627, B2 => 
                           n4844, ZN => n1855);
   U1354 : OAI22_X1 port map( A1 => n4705, A2 => n4850, B1 => n3650, B2 => 
                           n4846, ZN => n1878);
   U1355 : OAI22_X1 port map( A1 => n4621, A2 => n4768, B1 => n3302, B2 => 
                           n4764, ZN => n1530);
   U1356 : OAI22_X1 port map( A1 => n4624, A2 => n4768, B1 => n3303, B2 => 
                           n4764, ZN => n1531);
   U1357 : OAI22_X1 port map( A1 => n4627, A2 => n4768, B1 => n3304, B2 => 
                           n4764, ZN => n1532);
   U1358 : OAI22_X1 port map( A1 => n4630, A2 => n4768, B1 => n3305, B2 => 
                           n4764, ZN => n1533);
   U1359 : OAI22_X1 port map( A1 => n4633, A2 => n4768, B1 => n3306, B2 => 
                           n4764, ZN => n1534);
   U1360 : OAI22_X1 port map( A1 => n4636, A2 => n4768, B1 => n3307, B2 => 
                           n4764, ZN => n1535);
   U1361 : OAI22_X1 port map( A1 => n4705, A2 => n4770, B1 => n3330, B2 => 
                           n4766, ZN => n1558);
   U1362 : OAI22_X1 port map( A1 => n4621, A2 => n4776, B1 => n3334, B2 => 
                           n4772, ZN => n1562);
   U1363 : OAI22_X1 port map( A1 => n4624, A2 => n4776, B1 => n3335, B2 => 
                           n4772, ZN => n1563);
   U1364 : OAI22_X1 port map( A1 => n4627, A2 => n4776, B1 => n3336, B2 => 
                           n4772, ZN => n1564);
   U1365 : OAI22_X1 port map( A1 => n4630, A2 => n4776, B1 => n3337, B2 => 
                           n4772, ZN => n1565);
   U1366 : OAI22_X1 port map( A1 => n4633, A2 => n4776, B1 => n3338, B2 => 
                           n4772, ZN => n1566);
   U1367 : OAI22_X1 port map( A1 => n4636, A2 => n4776, B1 => n3339, B2 => 
                           n4772, ZN => n1567);
   U1368 : OAI22_X1 port map( A1 => n4705, A2 => n4778, B1 => n3362, B2 => 
                           n4774, ZN => n1590);
   U1369 : OAI22_X1 port map( A1 => n4621, A2 => n4784, B1 => n3366, B2 => 
                           n4780, ZN => n1594);
   U1370 : OAI22_X1 port map( A1 => n4624, A2 => n4784, B1 => n3367, B2 => 
                           n4780, ZN => n1595);
   U1371 : OAI22_X1 port map( A1 => n4627, A2 => n4784, B1 => n3368, B2 => 
                           n4780, ZN => n1596);
   U1372 : OAI22_X1 port map( A1 => n4630, A2 => n4784, B1 => n3369, B2 => 
                           n4780, ZN => n1597);
   U1373 : OAI22_X1 port map( A1 => n4633, A2 => n4784, B1 => n3370, B2 => 
                           n4780, ZN => n1598);
   U1374 : OAI22_X1 port map( A1 => n4636, A2 => n4784, B1 => n3371, B2 => 
                           n4780, ZN => n1599);
   U1375 : OAI22_X1 port map( A1 => n4705, A2 => n4786, B1 => n3394, B2 => 
                           n4782, ZN => n1622);
   U1376 : OAI22_X1 port map( A1 => n4621, A2 => n4792, B1 => n3398, B2 => 
                           n4788, ZN => n1626);
   U1377 : OAI22_X1 port map( A1 => n4624, A2 => n4792, B1 => n3399, B2 => 
                           n4788, ZN => n1627);
   U1378 : OAI22_X1 port map( A1 => n4627, A2 => n4792, B1 => n3400, B2 => 
                           n4788, ZN => n1628);
   U1379 : OAI22_X1 port map( A1 => n4630, A2 => n4792, B1 => n3401, B2 => 
                           n4788, ZN => n1629);
   U1380 : OAI22_X1 port map( A1 => n4633, A2 => n4792, B1 => n3402, B2 => 
                           n4788, ZN => n1630);
   U1381 : OAI22_X1 port map( A1 => n4636, A2 => n4792, B1 => n3403, B2 => 
                           n4788, ZN => n1631);
   U1382 : OAI22_X1 port map( A1 => n4705, A2 => n4794, B1 => n3426, B2 => 
                           n4790, ZN => n1654);
   U1383 : OAI22_X1 port map( A1 => n4621, A2 => n4800, B1 => n3430, B2 => 
                           n4796, ZN => n1658);
   U1384 : OAI22_X1 port map( A1 => n4624, A2 => n4800, B1 => n3431, B2 => 
                           n4796, ZN => n1659);
   U1385 : OAI22_X1 port map( A1 => n4627, A2 => n4800, B1 => n3432, B2 => 
                           n4796, ZN => n1660);
   U1386 : OAI22_X1 port map( A1 => n4630, A2 => n4800, B1 => n3433, B2 => 
                           n4796, ZN => n1661);
   U1387 : OAI22_X1 port map( A1 => n4633, A2 => n4800, B1 => n3434, B2 => 
                           n4796, ZN => n1662);
   U1388 : OAI22_X1 port map( A1 => n4636, A2 => n4800, B1 => n3435, B2 => 
                           n4796, ZN => n1663);
   U1389 : OAI22_X1 port map( A1 => n4705, A2 => n4802, B1 => n3458, B2 => 
                           n4798, ZN => n1686);
   U1390 : OAI22_X1 port map( A1 => n4621, A2 => n4816, B1 => n3494, B2 => 
                           n4812, ZN => n1722);
   U1391 : OAI22_X1 port map( A1 => n4624, A2 => n4816, B1 => n3495, B2 => 
                           n4812, ZN => n1723);
   U1392 : OAI22_X1 port map( A1 => n4627, A2 => n4816, B1 => n3496, B2 => 
                           n4812, ZN => n1724);
   U1393 : OAI22_X1 port map( A1 => n4630, A2 => n4816, B1 => n3497, B2 => 
                           n4812, ZN => n1725);
   U1394 : OAI22_X1 port map( A1 => n4633, A2 => n4816, B1 => n3498, B2 => 
                           n4812, ZN => n1726);
   U1395 : OAI22_X1 port map( A1 => n4636, A2 => n4816, B1 => n3499, B2 => 
                           n4812, ZN => n1727);
   U1396 : OAI22_X1 port map( A1 => n4705, A2 => n4818, B1 => n3522, B2 => 
                           n4814, ZN => n1750);
   U1397 : OAI22_X1 port map( A1 => n4621, A2 => n4832, B1 => n3558, B2 => 
                           n4828, ZN => n1786);
   U1398 : OAI22_X1 port map( A1 => n4624, A2 => n4832, B1 => n3559, B2 => 
                           n4828, ZN => n1787);
   U1399 : OAI22_X1 port map( A1 => n4627, A2 => n4832, B1 => n3560, B2 => 
                           n4828, ZN => n1788);
   U1400 : OAI22_X1 port map( A1 => n4630, A2 => n4832, B1 => n3561, B2 => 
                           n4828, ZN => n1789);
   U1401 : OAI22_X1 port map( A1 => n4633, A2 => n4832, B1 => n3562, B2 => 
                           n4828, ZN => n1790);
   U1402 : OAI22_X1 port map( A1 => n4636, A2 => n4832, B1 => n3563, B2 => 
                           n4828, ZN => n1791);
   U1403 : OAI22_X1 port map( A1 => n4705, A2 => n4834, B1 => n3586, B2 => 
                           n4830, ZN => n1814);
   U1404 : OAI22_X1 port map( A1 => n4612, A2 => n4760, B1 => n3267, B2 => 
                           n4756, ZN => n1495);
   U1405 : OAI22_X1 port map( A1 => n4615, A2 => n4760, B1 => n3268, B2 => 
                           n4756, ZN => n1496);
   U1406 : OAI22_X1 port map( A1 => n4618, A2 => n4760, B1 => n3269, B2 => 
                           n4756, ZN => n1497);
   U1407 : OAI22_X1 port map( A1 => n4642, A2 => n4760, B1 => n3277, B2 => 
                           n4756, ZN => n1505);
   U1408 : OAI22_X1 port map( A1 => n4645, A2 => n4761, B1 => n3278, B2 => 
                           n4756, ZN => n1506);
   U1409 : OAI22_X1 port map( A1 => n4648, A2 => n4761, B1 => n3279, B2 => 
                           n4757, ZN => n1507);
   U1410 : OAI22_X1 port map( A1 => n4651, A2 => n4761, B1 => n3280, B2 => 
                           n4757, ZN => n1508);
   U1411 : OAI22_X1 port map( A1 => n4654, A2 => n4761, B1 => n3281, B2 => 
                           n4757, ZN => n1509);
   U1412 : OAI22_X1 port map( A1 => n4657, A2 => n4761, B1 => n3282, B2 => 
                           n4757, ZN => n1510);
   U1413 : OAI22_X1 port map( A1 => n4660, A2 => n4761, B1 => n3283, B2 => 
                           n4757, ZN => n1511);
   U1414 : OAI22_X1 port map( A1 => n4663, A2 => n4761, B1 => n3284, B2 => 
                           n4757, ZN => n1512);
   U1415 : OAI22_X1 port map( A1 => n4666, A2 => n4761, B1 => n3285, B2 => 
                           n4757, ZN => n1513);
   U1416 : OAI22_X1 port map( A1 => n4669, A2 => n4761, B1 => n3286, B2 => 
                           n4757, ZN => n1514);
   U1417 : OAI22_X1 port map( A1 => n4672, A2 => n4761, B1 => n3287, B2 => 
                           n4757, ZN => n1515);
   U1418 : OAI22_X1 port map( A1 => n4675, A2 => n4761, B1 => n3288, B2 => 
                           n4757, ZN => n1516);
   U1419 : OAI22_X1 port map( A1 => n4678, A2 => n4761, B1 => n3289, B2 => 
                           n4757, ZN => n1517);
   U1420 : OAI22_X1 port map( A1 => n4681, A2 => n4762, B1 => n3290, B2 => 
                           n4757, ZN => n1518);
   U1421 : OAI22_X1 port map( A1 => n4684, A2 => n4762, B1 => n3291, B2 => 
                           n4758, ZN => n1519);
   U1422 : OAI22_X1 port map( A1 => n4687, A2 => n4762, B1 => n3292, B2 => 
                           n4758, ZN => n1520);
   U1423 : OAI22_X1 port map( A1 => n4690, A2 => n4762, B1 => n3293, B2 => 
                           n4758, ZN => n1521);
   U1424 : OAI22_X1 port map( A1 => n4693, A2 => n4762, B1 => n3294, B2 => 
                           n4758, ZN => n1522);
   U1425 : OAI22_X1 port map( A1 => n4696, A2 => n4762, B1 => n3295, B2 => 
                           n4758, ZN => n1523);
   U1426 : OAI22_X1 port map( A1 => n4699, A2 => n4762, B1 => n3296, B2 => 
                           n4758, ZN => n1524);
   U1427 : OAI22_X1 port map( A1 => n4702, A2 => n4762, B1 => n3297, B2 => 
                           n4758, ZN => n1525);
   U1428 : OAI22_X1 port map( A1 => n4612, A2 => n4808, B1 => n3459, B2 => 
                           n4804, ZN => n1687);
   U1429 : OAI22_X1 port map( A1 => n4615, A2 => n4808, B1 => n3460, B2 => 
                           n4804, ZN => n1688);
   U1430 : OAI22_X1 port map( A1 => n4618, A2 => n4808, B1 => n3461, B2 => 
                           n4804, ZN => n1689);
   U1431 : OAI22_X1 port map( A1 => n4642, A2 => n4808, B1 => n3469, B2 => 
                           n4804, ZN => n1697);
   U1432 : OAI22_X1 port map( A1 => n4645, A2 => n4809, B1 => n3470, B2 => 
                           n4804, ZN => n1698);
   U1433 : OAI22_X1 port map( A1 => n4648, A2 => n4809, B1 => n3471, B2 => 
                           n4805, ZN => n1699);
   U1434 : OAI22_X1 port map( A1 => n4651, A2 => n4809, B1 => n3472, B2 => 
                           n4805, ZN => n1700);
   U1435 : OAI22_X1 port map( A1 => n4654, A2 => n4809, B1 => n3473, B2 => 
                           n4805, ZN => n1701);
   U1436 : OAI22_X1 port map( A1 => n4657, A2 => n4809, B1 => n3474, B2 => 
                           n4805, ZN => n1702);
   U1437 : OAI22_X1 port map( A1 => n4660, A2 => n4809, B1 => n3475, B2 => 
                           n4805, ZN => n1703);
   U1438 : OAI22_X1 port map( A1 => n4663, A2 => n4809, B1 => n3476, B2 => 
                           n4805, ZN => n1704);
   U1439 : OAI22_X1 port map( A1 => n4666, A2 => n4809, B1 => n3477, B2 => 
                           n4805, ZN => n1705);
   U1440 : OAI22_X1 port map( A1 => n4669, A2 => n4809, B1 => n3478, B2 => 
                           n4805, ZN => n1706);
   U1441 : OAI22_X1 port map( A1 => n4672, A2 => n4809, B1 => n3479, B2 => 
                           n4805, ZN => n1707);
   U1442 : OAI22_X1 port map( A1 => n4675, A2 => n4809, B1 => n3480, B2 => 
                           n4805, ZN => n1708);
   U1443 : OAI22_X1 port map( A1 => n4678, A2 => n4809, B1 => n3481, B2 => 
                           n4805, ZN => n1709);
   U1444 : OAI22_X1 port map( A1 => n4681, A2 => n4810, B1 => n3482, B2 => 
                           n4805, ZN => n1710);
   U1445 : OAI22_X1 port map( A1 => n4684, A2 => n4810, B1 => n3483, B2 => 
                           n4806, ZN => n1711);
   U1446 : OAI22_X1 port map( A1 => n4687, A2 => n4810, B1 => n3484, B2 => 
                           n4806, ZN => n1712);
   U1447 : OAI22_X1 port map( A1 => n4690, A2 => n4810, B1 => n3485, B2 => 
                           n4806, ZN => n1713);
   U1448 : OAI22_X1 port map( A1 => n4693, A2 => n4810, B1 => n3486, B2 => 
                           n4806, ZN => n1714);
   U1449 : OAI22_X1 port map( A1 => n4696, A2 => n4810, B1 => n3487, B2 => 
                           n4806, ZN => n1715);
   U1450 : OAI22_X1 port map( A1 => n4699, A2 => n4810, B1 => n3488, B2 => 
                           n4806, ZN => n1716);
   U1451 : OAI22_X1 port map( A1 => n4702, A2 => n4810, B1 => n3489, B2 => 
                           n4806, ZN => n1717);
   U1452 : OAI22_X1 port map( A1 => n4611, A2 => n4864, B1 => n3683, B2 => 
                           n4860, ZN => n1911);
   U1453 : OAI22_X1 port map( A1 => n4614, A2 => n4864, B1 => n3684, B2 => 
                           n4860, ZN => n1912);
   U1454 : OAI22_X1 port map( A1 => n4617, A2 => n4864, B1 => n3685, B2 => 
                           n4860, ZN => n1913);
   U1455 : OAI22_X1 port map( A1 => n4641, A2 => n4864, B1 => n3693, B2 => 
                           n4860, ZN => n1921);
   U1456 : OAI22_X1 port map( A1 => n4644, A2 => n4865, B1 => n3694, B2 => 
                           n4860, ZN => n1922);
   U1457 : OAI22_X1 port map( A1 => n4647, A2 => n4865, B1 => n3695, B2 => 
                           n4861, ZN => n1923);
   U1458 : OAI22_X1 port map( A1 => n4650, A2 => n4865, B1 => n3696, B2 => 
                           n4861, ZN => n1924);
   U1459 : OAI22_X1 port map( A1 => n4653, A2 => n4865, B1 => n3697, B2 => 
                           n4861, ZN => n1925);
   U1460 : OAI22_X1 port map( A1 => n4656, A2 => n4865, B1 => n3698, B2 => 
                           n4861, ZN => n1926);
   U1461 : OAI22_X1 port map( A1 => n4659, A2 => n4865, B1 => n3699, B2 => 
                           n4861, ZN => n1927);
   U1462 : OAI22_X1 port map( A1 => n4662, A2 => n4865, B1 => n3700, B2 => 
                           n4861, ZN => n1928);
   U1463 : OAI22_X1 port map( A1 => n4665, A2 => n4865, B1 => n3701, B2 => 
                           n4861, ZN => n1929);
   U1464 : OAI22_X1 port map( A1 => n4668, A2 => n4865, B1 => n3702, B2 => 
                           n4861, ZN => n1930);
   U1465 : OAI22_X1 port map( A1 => n4671, A2 => n4865, B1 => n3703, B2 => 
                           n4861, ZN => n1931);
   U1466 : OAI22_X1 port map( A1 => n4674, A2 => n4865, B1 => n3704, B2 => 
                           n4861, ZN => n1932);
   U1467 : OAI22_X1 port map( A1 => n4677, A2 => n4865, B1 => n3705, B2 => 
                           n4861, ZN => n1933);
   U1468 : OAI22_X1 port map( A1 => n4680, A2 => n4866, B1 => n3706, B2 => 
                           n4861, ZN => n1934);
   U1469 : OAI22_X1 port map( A1 => n4683, A2 => n4866, B1 => n3707, B2 => 
                           n4862, ZN => n1935);
   U1470 : OAI22_X1 port map( A1 => n4686, A2 => n4866, B1 => n3708, B2 => 
                           n4862, ZN => n1936);
   U1471 : OAI22_X1 port map( A1 => n4689, A2 => n4866, B1 => n3709, B2 => 
                           n4862, ZN => n1937);
   U1472 : OAI22_X1 port map( A1 => n4692, A2 => n4866, B1 => n3710, B2 => 
                           n4862, ZN => n1938);
   U1473 : OAI22_X1 port map( A1 => n4695, A2 => n4866, B1 => n3711, B2 => 
                           n4862, ZN => n1939);
   U1474 : OAI22_X1 port map( A1 => n4698, A2 => n4866, B1 => n3712, B2 => 
                           n4862, ZN => n1940);
   U1475 : OAI22_X1 port map( A1 => n4701, A2 => n4866, B1 => n3713, B2 => 
                           n4862, ZN => n1941);
   U1476 : OAI22_X1 port map( A1 => n4611, A2 => n4888, B1 => n3779, B2 => 
                           n4884, ZN => n2007);
   U1477 : OAI22_X1 port map( A1 => n4614, A2 => n4888, B1 => n3780, B2 => 
                           n4884, ZN => n2008);
   U1478 : OAI22_X1 port map( A1 => n4617, A2 => n4888, B1 => n3781, B2 => 
                           n4884, ZN => n2009);
   U1479 : OAI22_X1 port map( A1 => n4641, A2 => n4888, B1 => n3789, B2 => 
                           n4884, ZN => n2017);
   U1480 : OAI22_X1 port map( A1 => n4644, A2 => n4889, B1 => n3790, B2 => 
                           n4884, ZN => n2018);
   U1481 : OAI22_X1 port map( A1 => n4647, A2 => n4889, B1 => n3791, B2 => 
                           n4885, ZN => n2019);
   U1482 : OAI22_X1 port map( A1 => n4650, A2 => n4889, B1 => n3792, B2 => 
                           n4885, ZN => n2020);
   U1483 : OAI22_X1 port map( A1 => n4653, A2 => n4889, B1 => n3793, B2 => 
                           n4885, ZN => n2021);
   U1484 : OAI22_X1 port map( A1 => n4656, A2 => n4889, B1 => n3794, B2 => 
                           n4885, ZN => n2022);
   U1485 : OAI22_X1 port map( A1 => n4659, A2 => n4889, B1 => n3795, B2 => 
                           n4885, ZN => n2023);
   U1486 : OAI22_X1 port map( A1 => n4662, A2 => n4889, B1 => n3796, B2 => 
                           n4885, ZN => n2024);
   U1487 : OAI22_X1 port map( A1 => n4665, A2 => n4889, B1 => n3797, B2 => 
                           n4885, ZN => n2025);
   U1488 : OAI22_X1 port map( A1 => n4668, A2 => n4889, B1 => n3798, B2 => 
                           n4885, ZN => n2026);
   U1489 : OAI22_X1 port map( A1 => n4671, A2 => n4889, B1 => n3799, B2 => 
                           n4885, ZN => n2027);
   U1490 : OAI22_X1 port map( A1 => n4674, A2 => n4889, B1 => n3800, B2 => 
                           n4885, ZN => n2028);
   U1491 : OAI22_X1 port map( A1 => n4677, A2 => n4889, B1 => n3801, B2 => 
                           n4885, ZN => n2029);
   U1492 : OAI22_X1 port map( A1 => n4680, A2 => n4890, B1 => n3802, B2 => 
                           n4885, ZN => n2030);
   U1493 : OAI22_X1 port map( A1 => n4683, A2 => n4890, B1 => n3803, B2 => 
                           n4886, ZN => n2031);
   U1494 : OAI22_X1 port map( A1 => n4686, A2 => n4890, B1 => n3804, B2 => 
                           n4886, ZN => n2032);
   U1495 : OAI22_X1 port map( A1 => n4689, A2 => n4890, B1 => n3805, B2 => 
                           n4886, ZN => n2033);
   U1496 : OAI22_X1 port map( A1 => n4692, A2 => n4890, B1 => n3806, B2 => 
                           n4886, ZN => n2034);
   U1497 : OAI22_X1 port map( A1 => n4695, A2 => n4890, B1 => n3807, B2 => 
                           n4886, ZN => n2035);
   U1498 : OAI22_X1 port map( A1 => n4698, A2 => n4890, B1 => n3808, B2 => 
                           n4886, ZN => n2036);
   U1499 : OAI22_X1 port map( A1 => n4701, A2 => n4890, B1 => n3809, B2 => 
                           n4886, ZN => n2037);
   U1500 : OAI22_X1 port map( A1 => n4611, A2 => n4896, B1 => n3811, B2 => 
                           n4892, ZN => n2039);
   U1501 : OAI22_X1 port map( A1 => n4614, A2 => n4896, B1 => n3812, B2 => 
                           n4892, ZN => n2040);
   U1502 : OAI22_X1 port map( A1 => n4617, A2 => n4896, B1 => n3813, B2 => 
                           n4892, ZN => n2041);
   U1503 : OAI22_X1 port map( A1 => n4641, A2 => n4896, B1 => n3821, B2 => 
                           n4892, ZN => n2049);
   U1504 : OAI22_X1 port map( A1 => n4644, A2 => n4897, B1 => n3822, B2 => 
                           n4892, ZN => n2050);
   U1505 : OAI22_X1 port map( A1 => n4647, A2 => n4897, B1 => n3823, B2 => 
                           n4893, ZN => n2051);
   U1506 : OAI22_X1 port map( A1 => n4650, A2 => n4897, B1 => n3824, B2 => 
                           n4893, ZN => n2052);
   U1507 : OAI22_X1 port map( A1 => n4653, A2 => n4897, B1 => n3825, B2 => 
                           n4893, ZN => n2053);
   U1508 : OAI22_X1 port map( A1 => n4656, A2 => n4897, B1 => n3826, B2 => 
                           n4893, ZN => n2054);
   U1509 : OAI22_X1 port map( A1 => n4659, A2 => n4897, B1 => n3827, B2 => 
                           n4893, ZN => n2055);
   U1510 : OAI22_X1 port map( A1 => n4662, A2 => n4897, B1 => n3828, B2 => 
                           n4893, ZN => n2056);
   U1511 : OAI22_X1 port map( A1 => n4665, A2 => n4897, B1 => n3829, B2 => 
                           n4893, ZN => n2057);
   U1512 : OAI22_X1 port map( A1 => n4668, A2 => n4897, B1 => n3830, B2 => 
                           n4893, ZN => n2058);
   U1513 : OAI22_X1 port map( A1 => n4671, A2 => n4897, B1 => n3831, B2 => 
                           n4893, ZN => n2059);
   U1514 : OAI22_X1 port map( A1 => n4674, A2 => n4897, B1 => n3832, B2 => 
                           n4893, ZN => n2060);
   U1515 : OAI22_X1 port map( A1 => n4677, A2 => n4897, B1 => n3833, B2 => 
                           n4893, ZN => n2061);
   U1516 : OAI22_X1 port map( A1 => n4680, A2 => n4898, B1 => n3834, B2 => 
                           n4893, ZN => n2062);
   U1517 : OAI22_X1 port map( A1 => n4683, A2 => n4898, B1 => n3835, B2 => 
                           n4894, ZN => n2063);
   U1518 : OAI22_X1 port map( A1 => n4686, A2 => n4898, B1 => n3836, B2 => 
                           n4894, ZN => n2064);
   U1519 : OAI22_X1 port map( A1 => n4689, A2 => n4898, B1 => n3837, B2 => 
                           n4894, ZN => n2065);
   U1520 : OAI22_X1 port map( A1 => n4692, A2 => n4898, B1 => n3838, B2 => 
                           n4894, ZN => n2066);
   U1521 : OAI22_X1 port map( A1 => n4695, A2 => n4898, B1 => n3839, B2 => 
                           n4894, ZN => n2067);
   U1522 : OAI22_X1 port map( A1 => n4698, A2 => n4898, B1 => n3840, B2 => 
                           n4894, ZN => n2068);
   U1523 : OAI22_X1 port map( A1 => n4701, A2 => n4898, B1 => n3841, B2 => 
                           n4894, ZN => n2069);
   U1524 : OAI22_X1 port map( A1 => n4611, A2 => n4920, B1 => n3907, B2 => 
                           n4916, ZN => n2135);
   U1525 : OAI22_X1 port map( A1 => n4614, A2 => n4920, B1 => n3908, B2 => 
                           n4916, ZN => n2136);
   U1526 : OAI22_X1 port map( A1 => n4617, A2 => n4920, B1 => n3909, B2 => 
                           n4916, ZN => n2137);
   U1527 : OAI22_X1 port map( A1 => n4641, A2 => n4920, B1 => n3917, B2 => 
                           n4916, ZN => n2145);
   U1528 : OAI22_X1 port map( A1 => n4644, A2 => n4921, B1 => n3918, B2 => 
                           n4916, ZN => n2146);
   U1529 : OAI22_X1 port map( A1 => n4647, A2 => n4921, B1 => n3919, B2 => 
                           n4917, ZN => n2147);
   U1530 : OAI22_X1 port map( A1 => n4650, A2 => n4921, B1 => n3920, B2 => 
                           n4917, ZN => n2148);
   U1531 : OAI22_X1 port map( A1 => n4653, A2 => n4921, B1 => n3921, B2 => 
                           n4917, ZN => n2149);
   U1532 : OAI22_X1 port map( A1 => n4656, A2 => n4921, B1 => n3922, B2 => 
                           n4917, ZN => n2150);
   U1533 : OAI22_X1 port map( A1 => n4659, A2 => n4921, B1 => n3923, B2 => 
                           n4917, ZN => n2151);
   U1534 : OAI22_X1 port map( A1 => n4662, A2 => n4921, B1 => n3924, B2 => 
                           n4917, ZN => n2152);
   U1535 : OAI22_X1 port map( A1 => n4665, A2 => n4921, B1 => n3925, B2 => 
                           n4917, ZN => n2153);
   U1536 : OAI22_X1 port map( A1 => n4668, A2 => n4921, B1 => n3926, B2 => 
                           n4917, ZN => n2154);
   U1537 : OAI22_X1 port map( A1 => n4671, A2 => n4921, B1 => n3927, B2 => 
                           n4917, ZN => n2155);
   U1538 : OAI22_X1 port map( A1 => n4674, A2 => n4921, B1 => n3928, B2 => 
                           n4917, ZN => n2156);
   U1539 : OAI22_X1 port map( A1 => n4677, A2 => n4921, B1 => n3929, B2 => 
                           n4917, ZN => n2157);
   U1540 : OAI22_X1 port map( A1 => n4680, A2 => n4922, B1 => n3930, B2 => 
                           n4917, ZN => n2158);
   U1541 : OAI22_X1 port map( A1 => n4683, A2 => n4922, B1 => n3931, B2 => 
                           n4918, ZN => n2159);
   U1542 : OAI22_X1 port map( A1 => n4686, A2 => n4922, B1 => n3932, B2 => 
                           n4918, ZN => n2160);
   U1543 : OAI22_X1 port map( A1 => n4689, A2 => n4922, B1 => n3933, B2 => 
                           n4918, ZN => n2161);
   U1544 : OAI22_X1 port map( A1 => n4692, A2 => n4922, B1 => n3934, B2 => 
                           n4918, ZN => n2162);
   U1545 : OAI22_X1 port map( A1 => n4695, A2 => n4922, B1 => n3935, B2 => 
                           n4918, ZN => n2163);
   U1546 : OAI22_X1 port map( A1 => n4698, A2 => n4922, B1 => n3936, B2 => 
                           n4918, ZN => n2164);
   U1547 : OAI22_X1 port map( A1 => n4701, A2 => n4922, B1 => n3937, B2 => 
                           n4918, ZN => n2165);
   U1548 : OAI22_X1 port map( A1 => n4611, A2 => n4928, B1 => n3939, B2 => 
                           n4924, ZN => n2167);
   U1549 : OAI22_X1 port map( A1 => n4614, A2 => n4928, B1 => n3940, B2 => 
                           n4924, ZN => n2168);
   U1550 : OAI22_X1 port map( A1 => n4617, A2 => n4928, B1 => n3941, B2 => 
                           n4924, ZN => n2169);
   U1551 : OAI22_X1 port map( A1 => n4641, A2 => n4928, B1 => n3949, B2 => 
                           n4924, ZN => n2177);
   U1552 : OAI22_X1 port map( A1 => n4644, A2 => n4929, B1 => n3950, B2 => 
                           n4924, ZN => n2178);
   U1553 : OAI22_X1 port map( A1 => n4647, A2 => n4929, B1 => n3951, B2 => 
                           n4925, ZN => n2179);
   U1554 : OAI22_X1 port map( A1 => n4650, A2 => n4929, B1 => n3952, B2 => 
                           n4925, ZN => n2180);
   U1555 : OAI22_X1 port map( A1 => n4653, A2 => n4929, B1 => n3953, B2 => 
                           n4925, ZN => n2181);
   U1556 : OAI22_X1 port map( A1 => n4656, A2 => n4929, B1 => n3954, B2 => 
                           n4925, ZN => n2182);
   U1557 : OAI22_X1 port map( A1 => n4659, A2 => n4929, B1 => n3955, B2 => 
                           n4925, ZN => n2183);
   U1558 : OAI22_X1 port map( A1 => n4662, A2 => n4929, B1 => n3956, B2 => 
                           n4925, ZN => n2184);
   U1559 : OAI22_X1 port map( A1 => n4665, A2 => n4929, B1 => n3957, B2 => 
                           n4925, ZN => n2185);
   U1560 : OAI22_X1 port map( A1 => n4668, A2 => n4929, B1 => n3958, B2 => 
                           n4925, ZN => n2186);
   U1561 : OAI22_X1 port map( A1 => n4671, A2 => n4929, B1 => n3959, B2 => 
                           n4925, ZN => n2187);
   U1562 : OAI22_X1 port map( A1 => n4674, A2 => n4929, B1 => n3960, B2 => 
                           n4925, ZN => n2188);
   U1563 : OAI22_X1 port map( A1 => n4677, A2 => n4929, B1 => n3961, B2 => 
                           n4925, ZN => n2189);
   U1564 : OAI22_X1 port map( A1 => n4680, A2 => n4930, B1 => n3962, B2 => 
                           n4925, ZN => n2190);
   U1565 : OAI22_X1 port map( A1 => n4683, A2 => n4930, B1 => n3963, B2 => 
                           n4926, ZN => n2191);
   U1566 : OAI22_X1 port map( A1 => n4686, A2 => n4930, B1 => n3964, B2 => 
                           n4926, ZN => n2192);
   U1567 : OAI22_X1 port map( A1 => n4689, A2 => n4930, B1 => n3965, B2 => 
                           n4926, ZN => n2193);
   U1568 : OAI22_X1 port map( A1 => n4692, A2 => n4930, B1 => n3966, B2 => 
                           n4926, ZN => n2194);
   U1569 : OAI22_X1 port map( A1 => n4695, A2 => n4930, B1 => n3967, B2 => 
                           n4926, ZN => n2195);
   U1570 : OAI22_X1 port map( A1 => n4698, A2 => n4930, B1 => n3968, B2 => 
                           n4926, ZN => n2196);
   U1571 : OAI22_X1 port map( A1 => n4701, A2 => n4930, B1 => n3969, B2 => 
                           n4926, ZN => n2197);
   U1572 : OAI22_X1 port map( A1 => n4611, A2 => n4952, B1 => n4035, B2 => 
                           n4948, ZN => n2263);
   U1573 : OAI22_X1 port map( A1 => n4614, A2 => n4952, B1 => n4036, B2 => 
                           n4948, ZN => n2264);
   U1574 : OAI22_X1 port map( A1 => n4617, A2 => n4952, B1 => n4037, B2 => 
                           n4948, ZN => n2265);
   U1575 : OAI22_X1 port map( A1 => n4641, A2 => n4952, B1 => n4045, B2 => 
                           n4948, ZN => n2273);
   U1576 : OAI22_X1 port map( A1 => n4644, A2 => n4953, B1 => n4046, B2 => 
                           n4948, ZN => n2274);
   U1577 : OAI22_X1 port map( A1 => n4647, A2 => n4953, B1 => n4047, B2 => 
                           n4949, ZN => n2275);
   U1578 : OAI22_X1 port map( A1 => n4650, A2 => n4953, B1 => n4048, B2 => 
                           n4949, ZN => n2276);
   U1579 : OAI22_X1 port map( A1 => n4653, A2 => n4953, B1 => n4049, B2 => 
                           n4949, ZN => n2277);
   U1580 : OAI22_X1 port map( A1 => n4656, A2 => n4953, B1 => n4050, B2 => 
                           n4949, ZN => n2278);
   U1581 : OAI22_X1 port map( A1 => n4659, A2 => n4953, B1 => n4051, B2 => 
                           n4949, ZN => n2279);
   U1582 : OAI22_X1 port map( A1 => n4662, A2 => n4953, B1 => n4052, B2 => 
                           n4949, ZN => n2280);
   U1583 : OAI22_X1 port map( A1 => n4665, A2 => n4953, B1 => n4053, B2 => 
                           n4949, ZN => n2281);
   U1584 : OAI22_X1 port map( A1 => n4668, A2 => n4953, B1 => n4054, B2 => 
                           n4949, ZN => n2282);
   U1585 : OAI22_X1 port map( A1 => n4671, A2 => n4953, B1 => n4055, B2 => 
                           n4949, ZN => n2283);
   U1586 : OAI22_X1 port map( A1 => n4674, A2 => n4953, B1 => n4056, B2 => 
                           n4949, ZN => n2284);
   U1587 : OAI22_X1 port map( A1 => n4677, A2 => n4953, B1 => n4057, B2 => 
                           n4949, ZN => n2285);
   U1588 : OAI22_X1 port map( A1 => n4680, A2 => n4954, B1 => n4058, B2 => 
                           n4949, ZN => n2286);
   U1589 : OAI22_X1 port map( A1 => n4683, A2 => n4954, B1 => n4059, B2 => 
                           n4950, ZN => n2287);
   U1590 : OAI22_X1 port map( A1 => n4686, A2 => n4954, B1 => n4060, B2 => 
                           n4950, ZN => n2288);
   U1591 : OAI22_X1 port map( A1 => n4689, A2 => n4954, B1 => n4061, B2 => 
                           n4950, ZN => n2289);
   U1592 : OAI22_X1 port map( A1 => n4692, A2 => n4954, B1 => n4062, B2 => 
                           n4950, ZN => n2290);
   U1593 : OAI22_X1 port map( A1 => n4695, A2 => n4954, B1 => n4063, B2 => 
                           n4950, ZN => n2291);
   U1594 : OAI22_X1 port map( A1 => n4698, A2 => n4954, B1 => n4064, B2 => 
                           n4950, ZN => n2292);
   U1595 : OAI22_X1 port map( A1 => n4701, A2 => n4954, B1 => n4065, B2 => 
                           n4950, ZN => n2293);
   U1596 : OAI22_X1 port map( A1 => n4611, A2 => n4872, B1 => n3715, B2 => 
                           n4868, ZN => n1943);
   U1597 : OAI22_X1 port map( A1 => n4614, A2 => n4872, B1 => n3716, B2 => 
                           n4868, ZN => n1944);
   U1598 : OAI22_X1 port map( A1 => n4617, A2 => n4872, B1 => n3717, B2 => 
                           n4868, ZN => n1945);
   U1599 : OAI22_X1 port map( A1 => n4641, A2 => n4872, B1 => n3725, B2 => 
                           n4868, ZN => n1953);
   U1600 : OAI22_X1 port map( A1 => n4644, A2 => n4873, B1 => n3726, B2 => 
                           n4868, ZN => n1954);
   U1601 : OAI22_X1 port map( A1 => n4647, A2 => n4873, B1 => n3727, B2 => 
                           n4869, ZN => n1955);
   U1602 : OAI22_X1 port map( A1 => n4650, A2 => n4873, B1 => n3728, B2 => 
                           n4869, ZN => n1956);
   U1603 : OAI22_X1 port map( A1 => n4653, A2 => n4873, B1 => n3729, B2 => 
                           n4869, ZN => n1957);
   U1604 : OAI22_X1 port map( A1 => n4656, A2 => n4873, B1 => n3730, B2 => 
                           n4869, ZN => n1958);
   U1605 : OAI22_X1 port map( A1 => n4659, A2 => n4873, B1 => n3731, B2 => 
                           n4869, ZN => n1959);
   U1606 : OAI22_X1 port map( A1 => n4662, A2 => n4873, B1 => n3732, B2 => 
                           n4869, ZN => n1960);
   U1607 : OAI22_X1 port map( A1 => n4665, A2 => n4873, B1 => n3733, B2 => 
                           n4869, ZN => n1961);
   U1608 : OAI22_X1 port map( A1 => n4668, A2 => n4873, B1 => n3734, B2 => 
                           n4869, ZN => n1962);
   U1609 : OAI22_X1 port map( A1 => n4671, A2 => n4873, B1 => n3735, B2 => 
                           n4869, ZN => n1963);
   U1610 : OAI22_X1 port map( A1 => n4674, A2 => n4873, B1 => n3736, B2 => 
                           n4869, ZN => n1964);
   U1611 : OAI22_X1 port map( A1 => n4677, A2 => n4873, B1 => n3737, B2 => 
                           n4869, ZN => n1965);
   U1612 : OAI22_X1 port map( A1 => n4680, A2 => n4874, B1 => n3738, B2 => 
                           n4869, ZN => n1966);
   U1613 : OAI22_X1 port map( A1 => n4683, A2 => n4874, B1 => n3739, B2 => 
                           n4870, ZN => n1967);
   U1614 : OAI22_X1 port map( A1 => n4686, A2 => n4874, B1 => n3740, B2 => 
                           n4870, ZN => n1968);
   U1615 : OAI22_X1 port map( A1 => n4689, A2 => n4874, B1 => n3741, B2 => 
                           n4870, ZN => n1969);
   U1616 : OAI22_X1 port map( A1 => n4692, A2 => n4874, B1 => n3742, B2 => 
                           n4870, ZN => n1970);
   U1617 : OAI22_X1 port map( A1 => n4695, A2 => n4874, B1 => n3743, B2 => 
                           n4870, ZN => n1971);
   U1618 : OAI22_X1 port map( A1 => n4698, A2 => n4874, B1 => n3744, B2 => 
                           n4870, ZN => n1972);
   U1619 : OAI22_X1 port map( A1 => n4701, A2 => n4874, B1 => n3745, B2 => 
                           n4870, ZN => n1973);
   U1620 : OAI22_X1 port map( A1 => n4611, A2 => n4880, B1 => n3747, B2 => 
                           n4876, ZN => n1975);
   U1621 : OAI22_X1 port map( A1 => n4614, A2 => n4880, B1 => n3748, B2 => 
                           n4876, ZN => n1976);
   U1622 : OAI22_X1 port map( A1 => n4617, A2 => n4880, B1 => n3749, B2 => 
                           n4876, ZN => n1977);
   U1623 : OAI22_X1 port map( A1 => n4641, A2 => n4880, B1 => n3757, B2 => 
                           n4876, ZN => n1985);
   U1624 : OAI22_X1 port map( A1 => n4644, A2 => n4881, B1 => n3758, B2 => 
                           n4876, ZN => n1986);
   U1625 : OAI22_X1 port map( A1 => n4647, A2 => n4881, B1 => n3759, B2 => 
                           n4877, ZN => n1987);
   U1626 : OAI22_X1 port map( A1 => n4650, A2 => n4881, B1 => n3760, B2 => 
                           n4877, ZN => n1988);
   U1627 : OAI22_X1 port map( A1 => n4653, A2 => n4881, B1 => n3761, B2 => 
                           n4877, ZN => n1989);
   U1628 : OAI22_X1 port map( A1 => n4656, A2 => n4881, B1 => n3762, B2 => 
                           n4877, ZN => n1990);
   U1629 : OAI22_X1 port map( A1 => n4659, A2 => n4881, B1 => n3763, B2 => 
                           n4877, ZN => n1991);
   U1630 : OAI22_X1 port map( A1 => n4662, A2 => n4881, B1 => n3764, B2 => 
                           n4877, ZN => n1992);
   U1631 : OAI22_X1 port map( A1 => n4665, A2 => n4881, B1 => n3765, B2 => 
                           n4877, ZN => n1993);
   U1632 : OAI22_X1 port map( A1 => n4668, A2 => n4881, B1 => n3766, B2 => 
                           n4877, ZN => n1994);
   U1633 : OAI22_X1 port map( A1 => n4671, A2 => n4881, B1 => n3767, B2 => 
                           n4877, ZN => n1995);
   U1634 : OAI22_X1 port map( A1 => n4674, A2 => n4881, B1 => n3768, B2 => 
                           n4877, ZN => n1996);
   U1635 : OAI22_X1 port map( A1 => n4677, A2 => n4881, B1 => n3769, B2 => 
                           n4877, ZN => n1997);
   U1636 : OAI22_X1 port map( A1 => n4680, A2 => n4882, B1 => n3770, B2 => 
                           n4877, ZN => n1998);
   U1637 : OAI22_X1 port map( A1 => n4683, A2 => n4882, B1 => n3771, B2 => 
                           n4878, ZN => n1999);
   U1638 : OAI22_X1 port map( A1 => n4686, A2 => n4882, B1 => n3772, B2 => 
                           n4878, ZN => n2000);
   U1639 : OAI22_X1 port map( A1 => n4689, A2 => n4882, B1 => n3773, B2 => 
                           n4878, ZN => n2001);
   U1640 : OAI22_X1 port map( A1 => n4692, A2 => n4882, B1 => n3774, B2 => 
                           n4878, ZN => n2002);
   U1641 : OAI22_X1 port map( A1 => n4695, A2 => n4882, B1 => n3775, B2 => 
                           n4878, ZN => n2003);
   U1642 : OAI22_X1 port map( A1 => n4698, A2 => n4882, B1 => n3776, B2 => 
                           n4878, ZN => n2004);
   U1643 : OAI22_X1 port map( A1 => n4701, A2 => n4882, B1 => n3777, B2 => 
                           n4878, ZN => n2005);
   U1644 : OAI22_X1 port map( A1 => n4611, A2 => n4904, B1 => n3843, B2 => 
                           n4900, ZN => n2071);
   U1645 : OAI22_X1 port map( A1 => n4614, A2 => n4904, B1 => n3844, B2 => 
                           n4900, ZN => n2072);
   U1646 : OAI22_X1 port map( A1 => n4617, A2 => n4904, B1 => n3845, B2 => 
                           n4900, ZN => n2073);
   U1647 : OAI22_X1 port map( A1 => n4641, A2 => n4904, B1 => n3853, B2 => 
                           n4900, ZN => n2081);
   U1648 : OAI22_X1 port map( A1 => n4644, A2 => n4905, B1 => n3854, B2 => 
                           n4900, ZN => n2082);
   U1649 : OAI22_X1 port map( A1 => n4647, A2 => n4905, B1 => n3855, B2 => 
                           n4901, ZN => n2083);
   U1650 : OAI22_X1 port map( A1 => n4650, A2 => n4905, B1 => n3856, B2 => 
                           n4901, ZN => n2084);
   U1651 : OAI22_X1 port map( A1 => n4653, A2 => n4905, B1 => n3857, B2 => 
                           n4901, ZN => n2085);
   U1652 : OAI22_X1 port map( A1 => n4656, A2 => n4905, B1 => n3858, B2 => 
                           n4901, ZN => n2086);
   U1653 : OAI22_X1 port map( A1 => n4659, A2 => n4905, B1 => n3859, B2 => 
                           n4901, ZN => n2087);
   U1654 : OAI22_X1 port map( A1 => n4662, A2 => n4905, B1 => n3860, B2 => 
                           n4901, ZN => n2088);
   U1655 : OAI22_X1 port map( A1 => n4665, A2 => n4905, B1 => n3861, B2 => 
                           n4901, ZN => n2089);
   U1656 : OAI22_X1 port map( A1 => n4668, A2 => n4905, B1 => n3862, B2 => 
                           n4901, ZN => n2090);
   U1657 : OAI22_X1 port map( A1 => n4671, A2 => n4905, B1 => n3863, B2 => 
                           n4901, ZN => n2091);
   U1658 : OAI22_X1 port map( A1 => n4674, A2 => n4905, B1 => n3864, B2 => 
                           n4901, ZN => n2092);
   U1659 : OAI22_X1 port map( A1 => n4677, A2 => n4905, B1 => n3865, B2 => 
                           n4901, ZN => n2093);
   U1660 : OAI22_X1 port map( A1 => n4680, A2 => n4906, B1 => n3866, B2 => 
                           n4901, ZN => n2094);
   U1661 : OAI22_X1 port map( A1 => n4683, A2 => n4906, B1 => n3867, B2 => 
                           n4902, ZN => n2095);
   U1662 : OAI22_X1 port map( A1 => n4686, A2 => n4906, B1 => n3868, B2 => 
                           n4902, ZN => n2096);
   U1663 : OAI22_X1 port map( A1 => n4689, A2 => n4906, B1 => n3869, B2 => 
                           n4902, ZN => n2097);
   U1664 : OAI22_X1 port map( A1 => n4692, A2 => n4906, B1 => n3870, B2 => 
                           n4902, ZN => n2098);
   U1665 : OAI22_X1 port map( A1 => n4695, A2 => n4906, B1 => n3871, B2 => 
                           n4902, ZN => n2099);
   U1666 : OAI22_X1 port map( A1 => n4698, A2 => n4906, B1 => n3872, B2 => 
                           n4902, ZN => n2100);
   U1667 : OAI22_X1 port map( A1 => n4701, A2 => n4906, B1 => n3873, B2 => 
                           n4902, ZN => n2101);
   U1668 : OAI22_X1 port map( A1 => n4611, A2 => n4912, B1 => n3875, B2 => 
                           n4908, ZN => n2103);
   U1669 : OAI22_X1 port map( A1 => n4614, A2 => n4912, B1 => n3876, B2 => 
                           n4908, ZN => n2104);
   U1670 : OAI22_X1 port map( A1 => n4617, A2 => n4912, B1 => n3877, B2 => 
                           n4908, ZN => n2105);
   U1671 : OAI22_X1 port map( A1 => n4641, A2 => n4912, B1 => n3885, B2 => 
                           n4908, ZN => n2113);
   U1672 : OAI22_X1 port map( A1 => n4644, A2 => n4913, B1 => n3886, B2 => 
                           n4908, ZN => n2114);
   U1673 : OAI22_X1 port map( A1 => n4647, A2 => n4913, B1 => n3887, B2 => 
                           n4909, ZN => n2115);
   U1674 : OAI22_X1 port map( A1 => n4650, A2 => n4913, B1 => n3888, B2 => 
                           n4909, ZN => n2116);
   U1675 : OAI22_X1 port map( A1 => n4653, A2 => n4913, B1 => n3889, B2 => 
                           n4909, ZN => n2117);
   U1676 : OAI22_X1 port map( A1 => n4656, A2 => n4913, B1 => n3890, B2 => 
                           n4909, ZN => n2118);
   U1677 : OAI22_X1 port map( A1 => n4659, A2 => n4913, B1 => n3891, B2 => 
                           n4909, ZN => n2119);
   U1678 : OAI22_X1 port map( A1 => n4662, A2 => n4913, B1 => n3892, B2 => 
                           n4909, ZN => n2120);
   U1679 : OAI22_X1 port map( A1 => n4665, A2 => n4913, B1 => n3893, B2 => 
                           n4909, ZN => n2121);
   U1680 : OAI22_X1 port map( A1 => n4668, A2 => n4913, B1 => n3894, B2 => 
                           n4909, ZN => n2122);
   U1681 : OAI22_X1 port map( A1 => n4671, A2 => n4913, B1 => n3895, B2 => 
                           n4909, ZN => n2123);
   U1682 : OAI22_X1 port map( A1 => n4674, A2 => n4913, B1 => n3896, B2 => 
                           n4909, ZN => n2124);
   U1683 : OAI22_X1 port map( A1 => n4677, A2 => n4913, B1 => n3897, B2 => 
                           n4909, ZN => n2125);
   U1684 : OAI22_X1 port map( A1 => n4680, A2 => n4914, B1 => n3898, B2 => 
                           n4909, ZN => n2126);
   U1685 : OAI22_X1 port map( A1 => n4683, A2 => n4914, B1 => n3899, B2 => 
                           n4910, ZN => n2127);
   U1686 : OAI22_X1 port map( A1 => n4686, A2 => n4914, B1 => n3900, B2 => 
                           n4910, ZN => n2128);
   U1687 : OAI22_X1 port map( A1 => n4689, A2 => n4914, B1 => n3901, B2 => 
                           n4910, ZN => n2129);
   U1688 : OAI22_X1 port map( A1 => n4692, A2 => n4914, B1 => n3902, B2 => 
                           n4910, ZN => n2130);
   U1689 : OAI22_X1 port map( A1 => n4695, A2 => n4914, B1 => n3903, B2 => 
                           n4910, ZN => n2131);
   U1690 : OAI22_X1 port map( A1 => n4698, A2 => n4914, B1 => n3904, B2 => 
                           n4910, ZN => n2132);
   U1691 : OAI22_X1 port map( A1 => n4701, A2 => n4914, B1 => n3905, B2 => 
                           n4910, ZN => n2133);
   U1692 : OAI22_X1 port map( A1 => n4611, A2 => n4936, B1 => n3971, B2 => 
                           n4932, ZN => n2199);
   U1693 : OAI22_X1 port map( A1 => n4614, A2 => n4936, B1 => n3972, B2 => 
                           n4932, ZN => n2200);
   U1694 : OAI22_X1 port map( A1 => n4617, A2 => n4936, B1 => n3973, B2 => 
                           n4932, ZN => n2201);
   U1695 : OAI22_X1 port map( A1 => n4641, A2 => n4936, B1 => n3981, B2 => 
                           n4932, ZN => n2209);
   U1696 : OAI22_X1 port map( A1 => n4644, A2 => n4937, B1 => n3982, B2 => 
                           n4932, ZN => n2210);
   U1697 : OAI22_X1 port map( A1 => n4647, A2 => n4937, B1 => n3983, B2 => 
                           n4933, ZN => n2211);
   U1698 : OAI22_X1 port map( A1 => n4650, A2 => n4937, B1 => n3984, B2 => 
                           n4933, ZN => n2212);
   U1699 : OAI22_X1 port map( A1 => n4653, A2 => n4937, B1 => n3985, B2 => 
                           n4933, ZN => n2213);
   U1700 : OAI22_X1 port map( A1 => n4656, A2 => n4937, B1 => n3986, B2 => 
                           n4933, ZN => n2214);
   U1701 : OAI22_X1 port map( A1 => n4659, A2 => n4937, B1 => n3987, B2 => 
                           n4933, ZN => n2215);
   U1702 : OAI22_X1 port map( A1 => n4662, A2 => n4937, B1 => n3988, B2 => 
                           n4933, ZN => n2216);
   U1703 : OAI22_X1 port map( A1 => n4665, A2 => n4937, B1 => n3989, B2 => 
                           n4933, ZN => n2217);
   U1704 : OAI22_X1 port map( A1 => n4668, A2 => n4937, B1 => n3990, B2 => 
                           n4933, ZN => n2218);
   U1705 : OAI22_X1 port map( A1 => n4671, A2 => n4937, B1 => n3991, B2 => 
                           n4933, ZN => n2219);
   U1706 : OAI22_X1 port map( A1 => n4674, A2 => n4937, B1 => n3992, B2 => 
                           n4933, ZN => n2220);
   U1707 : OAI22_X1 port map( A1 => n4677, A2 => n4937, B1 => n3993, B2 => 
                           n4933, ZN => n2221);
   U1708 : OAI22_X1 port map( A1 => n4680, A2 => n4938, B1 => n3994, B2 => 
                           n4933, ZN => n2222);
   U1709 : OAI22_X1 port map( A1 => n4683, A2 => n4938, B1 => n3995, B2 => 
                           n4934, ZN => n2223);
   U1710 : OAI22_X1 port map( A1 => n4686, A2 => n4938, B1 => n3996, B2 => 
                           n4934, ZN => n2224);
   U1711 : OAI22_X1 port map( A1 => n4689, A2 => n4938, B1 => n3997, B2 => 
                           n4934, ZN => n2225);
   U1712 : OAI22_X1 port map( A1 => n4692, A2 => n4938, B1 => n3998, B2 => 
                           n4934, ZN => n2226);
   U1713 : OAI22_X1 port map( A1 => n4695, A2 => n4938, B1 => n3999, B2 => 
                           n4934, ZN => n2227);
   U1714 : OAI22_X1 port map( A1 => n4698, A2 => n4938, B1 => n4000, B2 => 
                           n4934, ZN => n2228);
   U1715 : OAI22_X1 port map( A1 => n4701, A2 => n4938, B1 => n4001, B2 => 
                           n4934, ZN => n2229);
   U1716 : OAI22_X1 port map( A1 => n4611, A2 => n4944, B1 => n4003, B2 => 
                           n4940, ZN => n2231);
   U1717 : OAI22_X1 port map( A1 => n4614, A2 => n4944, B1 => n4004, B2 => 
                           n4940, ZN => n2232);
   U1718 : OAI22_X1 port map( A1 => n4617, A2 => n4944, B1 => n4005, B2 => 
                           n4940, ZN => n2233);
   U1719 : OAI22_X1 port map( A1 => n4641, A2 => n4944, B1 => n4013, B2 => 
                           n4940, ZN => n2241);
   U1720 : OAI22_X1 port map( A1 => n4644, A2 => n4945, B1 => n4014, B2 => 
                           n4940, ZN => n2242);
   U1721 : OAI22_X1 port map( A1 => n4647, A2 => n4945, B1 => n4015, B2 => 
                           n4941, ZN => n2243);
   U1722 : OAI22_X1 port map( A1 => n4650, A2 => n4945, B1 => n4016, B2 => 
                           n4941, ZN => n2244);
   U1723 : OAI22_X1 port map( A1 => n4653, A2 => n4945, B1 => n4017, B2 => 
                           n4941, ZN => n2245);
   U1724 : OAI22_X1 port map( A1 => n4656, A2 => n4945, B1 => n4018, B2 => 
                           n4941, ZN => n2246);
   U1725 : OAI22_X1 port map( A1 => n4659, A2 => n4945, B1 => n4019, B2 => 
                           n4941, ZN => n2247);
   U1726 : OAI22_X1 port map( A1 => n4662, A2 => n4945, B1 => n4020, B2 => 
                           n4941, ZN => n2248);
   U1727 : OAI22_X1 port map( A1 => n4665, A2 => n4945, B1 => n4021, B2 => 
                           n4941, ZN => n2249);
   U1728 : OAI22_X1 port map( A1 => n4668, A2 => n4945, B1 => n4022, B2 => 
                           n4941, ZN => n2250);
   U1729 : OAI22_X1 port map( A1 => n4671, A2 => n4945, B1 => n4023, B2 => 
                           n4941, ZN => n2251);
   U1730 : OAI22_X1 port map( A1 => n4674, A2 => n4945, B1 => n4024, B2 => 
                           n4941, ZN => n2252);
   U1731 : OAI22_X1 port map( A1 => n4677, A2 => n4945, B1 => n4025, B2 => 
                           n4941, ZN => n2253);
   U1732 : OAI22_X1 port map( A1 => n4680, A2 => n4946, B1 => n4026, B2 => 
                           n4941, ZN => n2254);
   U1733 : OAI22_X1 port map( A1 => n4683, A2 => n4946, B1 => n4027, B2 => 
                           n4942, ZN => n2255);
   U1734 : OAI22_X1 port map( A1 => n4686, A2 => n4946, B1 => n4028, B2 => 
                           n4942, ZN => n2256);
   U1735 : OAI22_X1 port map( A1 => n4689, A2 => n4946, B1 => n4029, B2 => 
                           n4942, ZN => n2257);
   U1736 : OAI22_X1 port map( A1 => n4692, A2 => n4946, B1 => n4030, B2 => 
                           n4942, ZN => n2258);
   U1737 : OAI22_X1 port map( A1 => n4695, A2 => n4946, B1 => n4031, B2 => 
                           n4942, ZN => n2259);
   U1738 : OAI22_X1 port map( A1 => n4698, A2 => n4946, B1 => n4032, B2 => 
                           n4942, ZN => n2260);
   U1739 : OAI22_X1 port map( A1 => n4701, A2 => n4946, B1 => n4033, B2 => 
                           n4942, ZN => n2261);
   U1740 : OAI22_X1 port map( A1 => n4612, A2 => n4824, B1 => n3523, B2 => 
                           n4820, ZN => n1751);
   U1741 : OAI22_X1 port map( A1 => n4615, A2 => n4824, B1 => n3524, B2 => 
                           n4820, ZN => n1752);
   U1742 : OAI22_X1 port map( A1 => n4618, A2 => n4824, B1 => n3525, B2 => 
                           n4820, ZN => n1753);
   U1743 : OAI22_X1 port map( A1 => n4642, A2 => n4824, B1 => n3533, B2 => 
                           n4820, ZN => n1761);
   U1744 : OAI22_X1 port map( A1 => n4645, A2 => n4825, B1 => n3534, B2 => 
                           n4820, ZN => n1762);
   U1745 : OAI22_X1 port map( A1 => n4648, A2 => n4825, B1 => n3535, B2 => 
                           n4821, ZN => n1763);
   U1746 : OAI22_X1 port map( A1 => n4651, A2 => n4825, B1 => n3536, B2 => 
                           n4821, ZN => n1764);
   U1747 : OAI22_X1 port map( A1 => n4654, A2 => n4825, B1 => n3537, B2 => 
                           n4821, ZN => n1765);
   U1748 : OAI22_X1 port map( A1 => n4657, A2 => n4825, B1 => n3538, B2 => 
                           n4821, ZN => n1766);
   U1749 : OAI22_X1 port map( A1 => n4660, A2 => n4825, B1 => n3539, B2 => 
                           n4821, ZN => n1767);
   U1750 : OAI22_X1 port map( A1 => n4663, A2 => n4825, B1 => n3540, B2 => 
                           n4821, ZN => n1768);
   U1751 : OAI22_X1 port map( A1 => n4666, A2 => n4825, B1 => n3541, B2 => 
                           n4821, ZN => n1769);
   U1752 : OAI22_X1 port map( A1 => n4669, A2 => n4825, B1 => n3542, B2 => 
                           n4821, ZN => n1770);
   U1753 : OAI22_X1 port map( A1 => n4672, A2 => n4825, B1 => n3543, B2 => 
                           n4821, ZN => n1771);
   U1754 : OAI22_X1 port map( A1 => n4675, A2 => n4825, B1 => n3544, B2 => 
                           n4821, ZN => n1772);
   U1755 : OAI22_X1 port map( A1 => n4678, A2 => n4825, B1 => n3545, B2 => 
                           n4821, ZN => n1773);
   U1756 : OAI22_X1 port map( A1 => n4612, A2 => n4856, B1 => n3651, B2 => 
                           n4852, ZN => n1879);
   U1757 : OAI22_X1 port map( A1 => n4615, A2 => n4856, B1 => n3652, B2 => 
                           n4852, ZN => n1880);
   U1758 : OAI22_X1 port map( A1 => n4618, A2 => n4856, B1 => n3653, B2 => 
                           n4852, ZN => n1881);
   U1759 : OAI22_X1 port map( A1 => n4642, A2 => n4856, B1 => n3661, B2 => 
                           n4852, ZN => n1889);
   U1760 : OAI22_X1 port map( A1 => n4645, A2 => n4857, B1 => n3662, B2 => 
                           n4852, ZN => n1890);
   U1761 : OAI22_X1 port map( A1 => n4648, A2 => n4857, B1 => n3663, B2 => 
                           n4853, ZN => n1891);
   U1762 : OAI22_X1 port map( A1 => n4651, A2 => n4857, B1 => n3664, B2 => 
                           n4853, ZN => n1892);
   U1763 : OAI22_X1 port map( A1 => n4654, A2 => n4857, B1 => n3665, B2 => 
                           n4853, ZN => n1893);
   U1764 : OAI22_X1 port map( A1 => n4657, A2 => n4857, B1 => n3666, B2 => 
                           n4853, ZN => n1894);
   U1765 : OAI22_X1 port map( A1 => n4660, A2 => n4857, B1 => n3667, B2 => 
                           n4853, ZN => n1895);
   U1766 : OAI22_X1 port map( A1 => n4663, A2 => n4857, B1 => n3668, B2 => 
                           n4853, ZN => n1896);
   U1767 : OAI22_X1 port map( A1 => n4666, A2 => n4857, B1 => n3669, B2 => 
                           n4853, ZN => n1897);
   U1768 : OAI22_X1 port map( A1 => n4669, A2 => n4857, B1 => n3670, B2 => 
                           n4853, ZN => n1898);
   U1769 : OAI22_X1 port map( A1 => n4672, A2 => n4857, B1 => n3671, B2 => 
                           n4853, ZN => n1899);
   U1770 : OAI22_X1 port map( A1 => n4675, A2 => n4857, B1 => n3672, B2 => 
                           n4853, ZN => n1900);
   U1771 : OAI22_X1 port map( A1 => n4678, A2 => n4857, B1 => n3673, B2 => 
                           n4853, ZN => n1901);
   U1772 : OAI22_X1 port map( A1 => n4681, A2 => n4858, B1 => n3674, B2 => 
                           n4853, ZN => n1902);
   U1773 : OAI22_X1 port map( A1 => n4684, A2 => n4858, B1 => n3675, B2 => 
                           n4854, ZN => n1903);
   U1774 : OAI22_X1 port map( A1 => n4687, A2 => n4858, B1 => n3676, B2 => 
                           n4854, ZN => n1904);
   U1775 : OAI22_X1 port map( A1 => n4690, A2 => n4858, B1 => n3677, B2 => 
                           n4854, ZN => n1905);
   U1776 : OAI22_X1 port map( A1 => n4693, A2 => n4858, B1 => n3678, B2 => 
                           n4854, ZN => n1906);
   U1777 : OAI22_X1 port map( A1 => n4696, A2 => n4858, B1 => n3679, B2 => 
                           n4854, ZN => n1907);
   U1778 : OAI22_X1 port map( A1 => n4699, A2 => n4858, B1 => n3680, B2 => 
                           n4854, ZN => n1908);
   U1779 : OAI22_X1 port map( A1 => n4702, A2 => n4858, B1 => n3681, B2 => 
                           n4854, ZN => n1909);
   U1780 : OAI22_X1 port map( A1 => n4612, A2 => n4840, B1 => n3587, B2 => 
                           n4836, ZN => n1815);
   U1781 : OAI22_X1 port map( A1 => n4615, A2 => n4840, B1 => n3588, B2 => 
                           n4836, ZN => n1816);
   U1782 : OAI22_X1 port map( A1 => n4618, A2 => n4840, B1 => n3589, B2 => 
                           n4836, ZN => n1817);
   U1783 : OAI22_X1 port map( A1 => n4642, A2 => n4840, B1 => n3597, B2 => 
                           n4836, ZN => n1825);
   U1784 : OAI22_X1 port map( A1 => n4645, A2 => n4841, B1 => n3598, B2 => 
                           n4836, ZN => n1826);
   U1785 : OAI22_X1 port map( A1 => n4648, A2 => n4841, B1 => n3599, B2 => 
                           n4837, ZN => n1827);
   U1786 : OAI22_X1 port map( A1 => n4651, A2 => n4841, B1 => n3600, B2 => 
                           n4837, ZN => n1828);
   U1787 : OAI22_X1 port map( A1 => n4654, A2 => n4841, B1 => n3601, B2 => 
                           n4837, ZN => n1829);
   U1788 : OAI22_X1 port map( A1 => n4657, A2 => n4841, B1 => n3602, B2 => 
                           n4837, ZN => n1830);
   U1789 : OAI22_X1 port map( A1 => n4660, A2 => n4841, B1 => n3603, B2 => 
                           n4837, ZN => n1831);
   U1790 : OAI22_X1 port map( A1 => n4663, A2 => n4841, B1 => n3604, B2 => 
                           n4837, ZN => n1832);
   U1791 : OAI22_X1 port map( A1 => n4666, A2 => n4841, B1 => n3605, B2 => 
                           n4837, ZN => n1833);
   U1792 : OAI22_X1 port map( A1 => n4669, A2 => n4841, B1 => n3606, B2 => 
                           n4837, ZN => n1834);
   U1793 : OAI22_X1 port map( A1 => n4672, A2 => n4841, B1 => n3607, B2 => 
                           n4837, ZN => n1835);
   U1794 : OAI22_X1 port map( A1 => n4675, A2 => n4841, B1 => n3608, B2 => 
                           n4837, ZN => n1836);
   U1795 : OAI22_X1 port map( A1 => n4678, A2 => n4841, B1 => n3609, B2 => 
                           n4837, ZN => n1837);
   U1796 : OAI22_X1 port map( A1 => n4681, A2 => n4842, B1 => n3610, B2 => 
                           n4837, ZN => n1838);
   U1797 : OAI22_X1 port map( A1 => n4684, A2 => n4842, B1 => n3611, B2 => 
                           n4838, ZN => n1839);
   U1798 : OAI22_X1 port map( A1 => n4687, A2 => n4842, B1 => n3612, B2 => 
                           n4838, ZN => n1840);
   U1799 : OAI22_X1 port map( A1 => n4690, A2 => n4842, B1 => n3613, B2 => 
                           n4838, ZN => n1841);
   U1800 : OAI22_X1 port map( A1 => n4693, A2 => n4842, B1 => n3614, B2 => 
                           n4838, ZN => n1842);
   U1801 : OAI22_X1 port map( A1 => n4696, A2 => n4842, B1 => n3615, B2 => 
                           n4838, ZN => n1843);
   U1802 : OAI22_X1 port map( A1 => n4699, A2 => n4842, B1 => n3616, B2 => 
                           n4838, ZN => n1844);
   U1803 : OAI22_X1 port map( A1 => n4702, A2 => n4842, B1 => n3617, B2 => 
                           n4838, ZN => n1845);
   U1804 : OAI22_X1 port map( A1 => n4612, A2 => n4848, B1 => n3619, B2 => 
                           n4844, ZN => n1847);
   U1805 : OAI22_X1 port map( A1 => n4615, A2 => n4848, B1 => n3620, B2 => 
                           n4844, ZN => n1848);
   U1806 : OAI22_X1 port map( A1 => n4618, A2 => n4848, B1 => n3621, B2 => 
                           n4844, ZN => n1849);
   U1807 : OAI22_X1 port map( A1 => n4642, A2 => n4848, B1 => n3629, B2 => 
                           n4844, ZN => n1857);
   U1808 : OAI22_X1 port map( A1 => n4645, A2 => n4849, B1 => n3630, B2 => 
                           n4844, ZN => n1858);
   U1809 : OAI22_X1 port map( A1 => n4648, A2 => n4849, B1 => n3631, B2 => 
                           n4845, ZN => n1859);
   U1810 : OAI22_X1 port map( A1 => n4651, A2 => n4849, B1 => n3632, B2 => 
                           n4845, ZN => n1860);
   U1811 : OAI22_X1 port map( A1 => n4654, A2 => n4849, B1 => n3633, B2 => 
                           n4845, ZN => n1861);
   U1812 : OAI22_X1 port map( A1 => n4657, A2 => n4849, B1 => n3634, B2 => 
                           n4845, ZN => n1862);
   U1813 : OAI22_X1 port map( A1 => n4660, A2 => n4849, B1 => n3635, B2 => 
                           n4845, ZN => n1863);
   U1814 : OAI22_X1 port map( A1 => n4663, A2 => n4849, B1 => n3636, B2 => 
                           n4845, ZN => n1864);
   U1815 : OAI22_X1 port map( A1 => n4666, A2 => n4849, B1 => n3637, B2 => 
                           n4845, ZN => n1865);
   U1816 : OAI22_X1 port map( A1 => n4669, A2 => n4849, B1 => n3638, B2 => 
                           n4845, ZN => n1866);
   U1817 : OAI22_X1 port map( A1 => n4672, A2 => n4849, B1 => n3639, B2 => 
                           n4845, ZN => n1867);
   U1818 : OAI22_X1 port map( A1 => n4675, A2 => n4849, B1 => n3640, B2 => 
                           n4845, ZN => n1868);
   U1819 : OAI22_X1 port map( A1 => n4678, A2 => n4849, B1 => n3641, B2 => 
                           n4845, ZN => n1869);
   U1820 : OAI22_X1 port map( A1 => n4681, A2 => n4850, B1 => n3642, B2 => 
                           n4845, ZN => n1870);
   U1821 : OAI22_X1 port map( A1 => n4684, A2 => n4850, B1 => n3643, B2 => 
                           n4846, ZN => n1871);
   U1822 : OAI22_X1 port map( A1 => n4687, A2 => n4850, B1 => n3644, B2 => 
                           n4846, ZN => n1872);
   U1823 : OAI22_X1 port map( A1 => n4690, A2 => n4850, B1 => n3645, B2 => 
                           n4846, ZN => n1873);
   U1824 : OAI22_X1 port map( A1 => n4693, A2 => n4850, B1 => n3646, B2 => 
                           n4846, ZN => n1874);
   U1825 : OAI22_X1 port map( A1 => n4696, A2 => n4850, B1 => n3647, B2 => 
                           n4846, ZN => n1875);
   U1826 : OAI22_X1 port map( A1 => n4699, A2 => n4850, B1 => n3648, B2 => 
                           n4846, ZN => n1876);
   U1827 : OAI22_X1 port map( A1 => n4702, A2 => n4850, B1 => n3649, B2 => 
                           n4846, ZN => n1877);
   U1828 : OAI22_X1 port map( A1 => n4612, A2 => n4768, B1 => n3299, B2 => 
                           n4764, ZN => n1527);
   U1829 : OAI22_X1 port map( A1 => n4615, A2 => n4768, B1 => n3300, B2 => 
                           n4764, ZN => n1528);
   U1830 : OAI22_X1 port map( A1 => n4618, A2 => n4768, B1 => n3301, B2 => 
                           n4764, ZN => n1529);
   U1831 : OAI22_X1 port map( A1 => n4642, A2 => n4768, B1 => n3309, B2 => 
                           n4764, ZN => n1537);
   U1832 : OAI22_X1 port map( A1 => n4645, A2 => n4769, B1 => n3310, B2 => 
                           n4764, ZN => n1538);
   U1833 : OAI22_X1 port map( A1 => n4648, A2 => n4769, B1 => n3311, B2 => 
                           n4765, ZN => n1539);
   U1834 : OAI22_X1 port map( A1 => n4651, A2 => n4769, B1 => n3312, B2 => 
                           n4765, ZN => n1540);
   U1835 : OAI22_X1 port map( A1 => n4654, A2 => n4769, B1 => n3313, B2 => 
                           n4765, ZN => n1541);
   U1836 : OAI22_X1 port map( A1 => n4657, A2 => n4769, B1 => n3314, B2 => 
                           n4765, ZN => n1542);
   U1837 : OAI22_X1 port map( A1 => n4660, A2 => n4769, B1 => n3315, B2 => 
                           n4765, ZN => n1543);
   U1838 : OAI22_X1 port map( A1 => n4663, A2 => n4769, B1 => n3316, B2 => 
                           n4765, ZN => n1544);
   U1839 : OAI22_X1 port map( A1 => n4666, A2 => n4769, B1 => n3317, B2 => 
                           n4765, ZN => n1545);
   U1840 : OAI22_X1 port map( A1 => n4669, A2 => n4769, B1 => n3318, B2 => 
                           n4765, ZN => n1546);
   U1841 : OAI22_X1 port map( A1 => n4672, A2 => n4769, B1 => n3319, B2 => 
                           n4765, ZN => n1547);
   U1842 : OAI22_X1 port map( A1 => n4675, A2 => n4769, B1 => n3320, B2 => 
                           n4765, ZN => n1548);
   U1843 : OAI22_X1 port map( A1 => n4678, A2 => n4769, B1 => n3321, B2 => 
                           n4765, ZN => n1549);
   U1844 : OAI22_X1 port map( A1 => n4612, A2 => n4776, B1 => n3331, B2 => 
                           n4772, ZN => n1559);
   U1845 : OAI22_X1 port map( A1 => n4615, A2 => n4776, B1 => n3332, B2 => 
                           n4772, ZN => n1560);
   U1846 : OAI22_X1 port map( A1 => n4618, A2 => n4776, B1 => n3333, B2 => 
                           n4772, ZN => n1561);
   U1847 : OAI22_X1 port map( A1 => n4642, A2 => n4776, B1 => n3341, B2 => 
                           n4772, ZN => n1569);
   U1848 : OAI22_X1 port map( A1 => n4645, A2 => n4777, B1 => n3342, B2 => 
                           n4772, ZN => n1570);
   U1849 : OAI22_X1 port map( A1 => n4648, A2 => n4777, B1 => n3343, B2 => 
                           n4773, ZN => n1571);
   U1850 : OAI22_X1 port map( A1 => n4651, A2 => n4777, B1 => n3344, B2 => 
                           n4773, ZN => n1572);
   U1851 : OAI22_X1 port map( A1 => n4654, A2 => n4777, B1 => n3345, B2 => 
                           n4773, ZN => n1573);
   U1852 : OAI22_X1 port map( A1 => n4657, A2 => n4777, B1 => n3346, B2 => 
                           n4773, ZN => n1574);
   U1853 : OAI22_X1 port map( A1 => n4660, A2 => n4777, B1 => n3347, B2 => 
                           n4773, ZN => n1575);
   U1854 : OAI22_X1 port map( A1 => n4663, A2 => n4777, B1 => n3348, B2 => 
                           n4773, ZN => n1576);
   U1855 : OAI22_X1 port map( A1 => n4666, A2 => n4777, B1 => n3349, B2 => 
                           n4773, ZN => n1577);
   U1856 : OAI22_X1 port map( A1 => n4669, A2 => n4777, B1 => n3350, B2 => 
                           n4773, ZN => n1578);
   U1857 : OAI22_X1 port map( A1 => n4672, A2 => n4777, B1 => n3351, B2 => 
                           n4773, ZN => n1579);
   U1858 : OAI22_X1 port map( A1 => n4675, A2 => n4777, B1 => n3352, B2 => 
                           n4773, ZN => n1580);
   U1859 : OAI22_X1 port map( A1 => n4678, A2 => n4777, B1 => n3353, B2 => 
                           n4773, ZN => n1581);
   U1860 : OAI22_X1 port map( A1 => n4612, A2 => n4784, B1 => n3363, B2 => 
                           n4780, ZN => n1591);
   U1861 : OAI22_X1 port map( A1 => n4615, A2 => n4784, B1 => n3364, B2 => 
                           n4780, ZN => n1592);
   U1862 : OAI22_X1 port map( A1 => n4618, A2 => n4784, B1 => n3365, B2 => 
                           n4780, ZN => n1593);
   U1863 : OAI22_X1 port map( A1 => n4642, A2 => n4784, B1 => n3373, B2 => 
                           n4780, ZN => n1601);
   U1864 : OAI22_X1 port map( A1 => n4645, A2 => n4785, B1 => n3374, B2 => 
                           n4780, ZN => n1602);
   U1865 : OAI22_X1 port map( A1 => n4648, A2 => n4785, B1 => n3375, B2 => 
                           n4781, ZN => n1603);
   U1866 : OAI22_X1 port map( A1 => n4651, A2 => n4785, B1 => n3376, B2 => 
                           n4781, ZN => n1604);
   U1867 : OAI22_X1 port map( A1 => n4654, A2 => n4785, B1 => n3377, B2 => 
                           n4781, ZN => n1605);
   U1868 : OAI22_X1 port map( A1 => n4657, A2 => n4785, B1 => n3378, B2 => 
                           n4781, ZN => n1606);
   U1869 : OAI22_X1 port map( A1 => n4660, A2 => n4785, B1 => n3379, B2 => 
                           n4781, ZN => n1607);
   U1870 : OAI22_X1 port map( A1 => n4663, A2 => n4785, B1 => n3380, B2 => 
                           n4781, ZN => n1608);
   U1871 : OAI22_X1 port map( A1 => n4666, A2 => n4785, B1 => n3381, B2 => 
                           n4781, ZN => n1609);
   U1872 : OAI22_X1 port map( A1 => n4669, A2 => n4785, B1 => n3382, B2 => 
                           n4781, ZN => n1610);
   U1873 : OAI22_X1 port map( A1 => n4672, A2 => n4785, B1 => n3383, B2 => 
                           n4781, ZN => n1611);
   U1874 : OAI22_X1 port map( A1 => n4675, A2 => n4785, B1 => n3384, B2 => 
                           n4781, ZN => n1612);
   U1875 : OAI22_X1 port map( A1 => n4678, A2 => n4785, B1 => n3385, B2 => 
                           n4781, ZN => n1613);
   U1876 : OAI22_X1 port map( A1 => n4612, A2 => n4792, B1 => n3395, B2 => 
                           n4788, ZN => n1623);
   U1877 : OAI22_X1 port map( A1 => n4615, A2 => n4792, B1 => n3396, B2 => 
                           n4788, ZN => n1624);
   U1878 : OAI22_X1 port map( A1 => n4618, A2 => n4792, B1 => n3397, B2 => 
                           n4788, ZN => n1625);
   U1879 : OAI22_X1 port map( A1 => n4642, A2 => n4792, B1 => n3405, B2 => 
                           n4788, ZN => n1633);
   U1880 : OAI22_X1 port map( A1 => n4645, A2 => n4793, B1 => n3406, B2 => 
                           n4788, ZN => n1634);
   U1881 : OAI22_X1 port map( A1 => n4648, A2 => n4793, B1 => n3407, B2 => 
                           n4789, ZN => n1635);
   U1882 : OAI22_X1 port map( A1 => n4651, A2 => n4793, B1 => n3408, B2 => 
                           n4789, ZN => n1636);
   U1883 : OAI22_X1 port map( A1 => n4654, A2 => n4793, B1 => n3409, B2 => 
                           n4789, ZN => n1637);
   U1884 : OAI22_X1 port map( A1 => n4657, A2 => n4793, B1 => n3410, B2 => 
                           n4789, ZN => n1638);
   U1885 : OAI22_X1 port map( A1 => n4660, A2 => n4793, B1 => n3411, B2 => 
                           n4789, ZN => n1639);
   U1886 : OAI22_X1 port map( A1 => n4663, A2 => n4793, B1 => n3412, B2 => 
                           n4789, ZN => n1640);
   U1887 : OAI22_X1 port map( A1 => n4666, A2 => n4793, B1 => n3413, B2 => 
                           n4789, ZN => n1641);
   U1888 : OAI22_X1 port map( A1 => n4669, A2 => n4793, B1 => n3414, B2 => 
                           n4789, ZN => n1642);
   U1889 : OAI22_X1 port map( A1 => n4672, A2 => n4793, B1 => n3415, B2 => 
                           n4789, ZN => n1643);
   U1890 : OAI22_X1 port map( A1 => n4675, A2 => n4793, B1 => n3416, B2 => 
                           n4789, ZN => n1644);
   U1891 : OAI22_X1 port map( A1 => n4678, A2 => n4793, B1 => n3417, B2 => 
                           n4789, ZN => n1645);
   U1892 : OAI22_X1 port map( A1 => n4612, A2 => n4800, B1 => n3427, B2 => 
                           n4796, ZN => n1655);
   U1893 : OAI22_X1 port map( A1 => n4615, A2 => n4800, B1 => n3428, B2 => 
                           n4796, ZN => n1656);
   U1894 : OAI22_X1 port map( A1 => n4618, A2 => n4800, B1 => n3429, B2 => 
                           n4796, ZN => n1657);
   U1895 : OAI22_X1 port map( A1 => n4642, A2 => n4800, B1 => n3437, B2 => 
                           n4796, ZN => n1665);
   U1896 : OAI22_X1 port map( A1 => n4645, A2 => n4801, B1 => n3438, B2 => 
                           n4796, ZN => n1666);
   U1897 : OAI22_X1 port map( A1 => n4648, A2 => n4801, B1 => n3439, B2 => 
                           n4797, ZN => n1667);
   U1898 : OAI22_X1 port map( A1 => n4651, A2 => n4801, B1 => n3440, B2 => 
                           n4797, ZN => n1668);
   U1899 : OAI22_X1 port map( A1 => n4654, A2 => n4801, B1 => n3441, B2 => 
                           n4797, ZN => n1669);
   U1900 : OAI22_X1 port map( A1 => n4657, A2 => n4801, B1 => n3442, B2 => 
                           n4797, ZN => n1670);
   U1901 : OAI22_X1 port map( A1 => n4660, A2 => n4801, B1 => n3443, B2 => 
                           n4797, ZN => n1671);
   U1902 : OAI22_X1 port map( A1 => n4663, A2 => n4801, B1 => n3444, B2 => 
                           n4797, ZN => n1672);
   U1903 : OAI22_X1 port map( A1 => n4666, A2 => n4801, B1 => n3445, B2 => 
                           n4797, ZN => n1673);
   U1904 : OAI22_X1 port map( A1 => n4669, A2 => n4801, B1 => n3446, B2 => 
                           n4797, ZN => n1674);
   U1905 : OAI22_X1 port map( A1 => n4672, A2 => n4801, B1 => n3447, B2 => 
                           n4797, ZN => n1675);
   U1906 : OAI22_X1 port map( A1 => n4675, A2 => n4801, B1 => n3448, B2 => 
                           n4797, ZN => n1676);
   U1907 : OAI22_X1 port map( A1 => n4678, A2 => n4801, B1 => n3449, B2 => 
                           n4797, ZN => n1677);
   U1908 : OAI22_X1 port map( A1 => n4612, A2 => n4816, B1 => n3491, B2 => 
                           n4812, ZN => n1719);
   U1909 : OAI22_X1 port map( A1 => n4615, A2 => n4816, B1 => n3492, B2 => 
                           n4812, ZN => n1720);
   U1910 : OAI22_X1 port map( A1 => n4618, A2 => n4816, B1 => n3493, B2 => 
                           n4812, ZN => n1721);
   U1911 : OAI22_X1 port map( A1 => n4642, A2 => n4816, B1 => n3501, B2 => 
                           n4812, ZN => n1729);
   U1912 : OAI22_X1 port map( A1 => n4645, A2 => n4817, B1 => n3502, B2 => 
                           n4812, ZN => n1730);
   U1913 : OAI22_X1 port map( A1 => n4648, A2 => n4817, B1 => n3503, B2 => 
                           n4813, ZN => n1731);
   U1914 : OAI22_X1 port map( A1 => n4651, A2 => n4817, B1 => n3504, B2 => 
                           n4813, ZN => n1732);
   U1915 : OAI22_X1 port map( A1 => n4654, A2 => n4817, B1 => n3505, B2 => 
                           n4813, ZN => n1733);
   U1916 : OAI22_X1 port map( A1 => n4657, A2 => n4817, B1 => n3506, B2 => 
                           n4813, ZN => n1734);
   U1917 : OAI22_X1 port map( A1 => n4660, A2 => n4817, B1 => n3507, B2 => 
                           n4813, ZN => n1735);
   U1918 : OAI22_X1 port map( A1 => n4663, A2 => n4817, B1 => n3508, B2 => 
                           n4813, ZN => n1736);
   U1919 : OAI22_X1 port map( A1 => n4666, A2 => n4817, B1 => n3509, B2 => 
                           n4813, ZN => n1737);
   U1920 : OAI22_X1 port map( A1 => n4669, A2 => n4817, B1 => n3510, B2 => 
                           n4813, ZN => n1738);
   U1921 : OAI22_X1 port map( A1 => n4672, A2 => n4817, B1 => n3511, B2 => 
                           n4813, ZN => n1739);
   U1922 : OAI22_X1 port map( A1 => n4675, A2 => n4817, B1 => n3512, B2 => 
                           n4813, ZN => n1740);
   U1923 : OAI22_X1 port map( A1 => n4678, A2 => n4817, B1 => n3513, B2 => 
                           n4813, ZN => n1741);
   U1924 : OAI22_X1 port map( A1 => n4612, A2 => n4832, B1 => n3555, B2 => 
                           n4828, ZN => n1783);
   U1925 : OAI22_X1 port map( A1 => n4615, A2 => n4832, B1 => n3556, B2 => 
                           n4828, ZN => n1784);
   U1926 : OAI22_X1 port map( A1 => n4618, A2 => n4832, B1 => n3557, B2 => 
                           n4828, ZN => n1785);
   U1927 : OAI22_X1 port map( A1 => n4642, A2 => n4832, B1 => n3565, B2 => 
                           n4828, ZN => n1793);
   U1928 : OAI22_X1 port map( A1 => n4645, A2 => n4833, B1 => n3566, B2 => 
                           n4828, ZN => n1794);
   U1929 : OAI22_X1 port map( A1 => n4648, A2 => n4833, B1 => n3567, B2 => 
                           n4829, ZN => n1795);
   U1930 : OAI22_X1 port map( A1 => n4651, A2 => n4833, B1 => n3568, B2 => 
                           n4829, ZN => n1796);
   U1931 : OAI22_X1 port map( A1 => n4654, A2 => n4833, B1 => n3569, B2 => 
                           n4829, ZN => n1797);
   U1932 : OAI22_X1 port map( A1 => n4657, A2 => n4833, B1 => n3570, B2 => 
                           n4829, ZN => n1798);
   U1933 : OAI22_X1 port map( A1 => n4660, A2 => n4833, B1 => n3571, B2 => 
                           n4829, ZN => n1799);
   U1934 : OAI22_X1 port map( A1 => n4663, A2 => n4833, B1 => n3572, B2 => 
                           n4829, ZN => n1800);
   U1935 : OAI22_X1 port map( A1 => n4666, A2 => n4833, B1 => n3573, B2 => 
                           n4829, ZN => n1801);
   U1936 : OAI22_X1 port map( A1 => n4669, A2 => n4833, B1 => n3574, B2 => 
                           n4829, ZN => n1802);
   U1937 : OAI22_X1 port map( A1 => n4672, A2 => n4833, B1 => n3575, B2 => 
                           n4829, ZN => n1803);
   U1938 : OAI22_X1 port map( A1 => n4675, A2 => n4833, B1 => n3576, B2 => 
                           n4829, ZN => n1804);
   U1939 : OAI22_X1 port map( A1 => n4678, A2 => n4833, B1 => n3577, B2 => 
                           n4829, ZN => n1805);
   U1940 : OAI22_X1 port map( A1 => n4681, A2 => n4826, B1 => n3546, B2 => 
                           n4821, ZN => n1774);
   U1941 : OAI22_X1 port map( A1 => n4684, A2 => n4826, B1 => n3547, B2 => 
                           n4822, ZN => n1775);
   U1942 : OAI22_X1 port map( A1 => n4687, A2 => n4826, B1 => n3548, B2 => 
                           n4822, ZN => n1776);
   U1943 : OAI22_X1 port map( A1 => n4690, A2 => n4826, B1 => n3549, B2 => 
                           n4822, ZN => n1777);
   U1944 : OAI22_X1 port map( A1 => n4693, A2 => n4826, B1 => n3550, B2 => 
                           n4822, ZN => n1778);
   U1945 : OAI22_X1 port map( A1 => n4696, A2 => n4826, B1 => n3551, B2 => 
                           n4822, ZN => n1779);
   U1946 : OAI22_X1 port map( A1 => n4699, A2 => n4826, B1 => n3552, B2 => 
                           n4822, ZN => n1780);
   U1947 : OAI22_X1 port map( A1 => n4702, A2 => n4826, B1 => n3553, B2 => 
                           n4822, ZN => n1781);
   U1948 : OAI22_X1 port map( A1 => n4681, A2 => n4770, B1 => n3322, B2 => 
                           n4765, ZN => n1550);
   U1949 : OAI22_X1 port map( A1 => n4684, A2 => n4770, B1 => n3323, B2 => 
                           n4766, ZN => n1551);
   U1950 : OAI22_X1 port map( A1 => n4687, A2 => n4770, B1 => n3324, B2 => 
                           n4766, ZN => n1552);
   U1951 : OAI22_X1 port map( A1 => n4690, A2 => n4770, B1 => n3325, B2 => 
                           n4766, ZN => n1553);
   U1952 : OAI22_X1 port map( A1 => n4693, A2 => n4770, B1 => n3326, B2 => 
                           n4766, ZN => n1554);
   U1953 : OAI22_X1 port map( A1 => n4696, A2 => n4770, B1 => n3327, B2 => 
                           n4766, ZN => n1555);
   U1954 : OAI22_X1 port map( A1 => n4699, A2 => n4770, B1 => n3328, B2 => 
                           n4766, ZN => n1556);
   U1955 : OAI22_X1 port map( A1 => n4702, A2 => n4770, B1 => n3329, B2 => 
                           n4766, ZN => n1557);
   U1956 : OAI22_X1 port map( A1 => n4681, A2 => n4778, B1 => n3354, B2 => 
                           n4773, ZN => n1582);
   U1957 : OAI22_X1 port map( A1 => n4684, A2 => n4778, B1 => n3355, B2 => 
                           n4774, ZN => n1583);
   U1958 : OAI22_X1 port map( A1 => n4687, A2 => n4778, B1 => n3356, B2 => 
                           n4774, ZN => n1584);
   U1959 : OAI22_X1 port map( A1 => n4690, A2 => n4778, B1 => n3357, B2 => 
                           n4774, ZN => n1585);
   U1960 : OAI22_X1 port map( A1 => n4693, A2 => n4778, B1 => n3358, B2 => 
                           n4774, ZN => n1586);
   U1961 : OAI22_X1 port map( A1 => n4696, A2 => n4778, B1 => n3359, B2 => 
                           n4774, ZN => n1587);
   U1962 : OAI22_X1 port map( A1 => n4699, A2 => n4778, B1 => n3360, B2 => 
                           n4774, ZN => n1588);
   U1963 : OAI22_X1 port map( A1 => n4702, A2 => n4778, B1 => n3361, B2 => 
                           n4774, ZN => n1589);
   U1964 : OAI22_X1 port map( A1 => n4681, A2 => n4786, B1 => n3386, B2 => 
                           n4781, ZN => n1614);
   U1965 : OAI22_X1 port map( A1 => n4684, A2 => n4786, B1 => n3387, B2 => 
                           n4782, ZN => n1615);
   U1966 : OAI22_X1 port map( A1 => n4687, A2 => n4786, B1 => n3388, B2 => 
                           n4782, ZN => n1616);
   U1967 : OAI22_X1 port map( A1 => n4690, A2 => n4786, B1 => n3389, B2 => 
                           n4782, ZN => n1617);
   U1968 : OAI22_X1 port map( A1 => n4693, A2 => n4786, B1 => n3390, B2 => 
                           n4782, ZN => n1618);
   U1969 : OAI22_X1 port map( A1 => n4696, A2 => n4786, B1 => n3391, B2 => 
                           n4782, ZN => n1619);
   U1970 : OAI22_X1 port map( A1 => n4699, A2 => n4786, B1 => n3392, B2 => 
                           n4782, ZN => n1620);
   U1971 : OAI22_X1 port map( A1 => n4702, A2 => n4786, B1 => n3393, B2 => 
                           n4782, ZN => n1621);
   U1972 : OAI22_X1 port map( A1 => n4681, A2 => n4794, B1 => n3418, B2 => 
                           n4789, ZN => n1646);
   U1973 : OAI22_X1 port map( A1 => n4684, A2 => n4794, B1 => n3419, B2 => 
                           n4790, ZN => n1647);
   U1974 : OAI22_X1 port map( A1 => n4687, A2 => n4794, B1 => n3420, B2 => 
                           n4790, ZN => n1648);
   U1975 : OAI22_X1 port map( A1 => n4690, A2 => n4794, B1 => n3421, B2 => 
                           n4790, ZN => n1649);
   U1976 : OAI22_X1 port map( A1 => n4693, A2 => n4794, B1 => n3422, B2 => 
                           n4790, ZN => n1650);
   U1977 : OAI22_X1 port map( A1 => n4696, A2 => n4794, B1 => n3423, B2 => 
                           n4790, ZN => n1651);
   U1978 : OAI22_X1 port map( A1 => n4699, A2 => n4794, B1 => n3424, B2 => 
                           n4790, ZN => n1652);
   U1979 : OAI22_X1 port map( A1 => n4702, A2 => n4794, B1 => n3425, B2 => 
                           n4790, ZN => n1653);
   U1980 : OAI22_X1 port map( A1 => n4681, A2 => n4802, B1 => n3450, B2 => 
                           n4797, ZN => n1678);
   U1981 : OAI22_X1 port map( A1 => n4684, A2 => n4802, B1 => n3451, B2 => 
                           n4798, ZN => n1679);
   U1982 : OAI22_X1 port map( A1 => n4687, A2 => n4802, B1 => n3452, B2 => 
                           n4798, ZN => n1680);
   U1983 : OAI22_X1 port map( A1 => n4690, A2 => n4802, B1 => n3453, B2 => 
                           n4798, ZN => n1681);
   U1984 : OAI22_X1 port map( A1 => n4693, A2 => n4802, B1 => n3454, B2 => 
                           n4798, ZN => n1682);
   U1985 : OAI22_X1 port map( A1 => n4696, A2 => n4802, B1 => n3455, B2 => 
                           n4798, ZN => n1683);
   U1986 : OAI22_X1 port map( A1 => n4699, A2 => n4802, B1 => n3456, B2 => 
                           n4798, ZN => n1684);
   U1987 : OAI22_X1 port map( A1 => n4702, A2 => n4802, B1 => n3457, B2 => 
                           n4798, ZN => n1685);
   U1988 : OAI22_X1 port map( A1 => n4681, A2 => n4818, B1 => n3514, B2 => 
                           n4813, ZN => n1742);
   U1989 : OAI22_X1 port map( A1 => n4684, A2 => n4818, B1 => n3515, B2 => 
                           n4814, ZN => n1743);
   U1990 : OAI22_X1 port map( A1 => n4687, A2 => n4818, B1 => n3516, B2 => 
                           n4814, ZN => n1744);
   U1991 : OAI22_X1 port map( A1 => n4690, A2 => n4818, B1 => n3517, B2 => 
                           n4814, ZN => n1745);
   U1992 : OAI22_X1 port map( A1 => n4693, A2 => n4818, B1 => n3518, B2 => 
                           n4814, ZN => n1746);
   U1993 : OAI22_X1 port map( A1 => n4696, A2 => n4818, B1 => n3519, B2 => 
                           n4814, ZN => n1747);
   U1994 : OAI22_X1 port map( A1 => n4699, A2 => n4818, B1 => n3520, B2 => 
                           n4814, ZN => n1748);
   U1995 : OAI22_X1 port map( A1 => n4702, A2 => n4818, B1 => n3521, B2 => 
                           n4814, ZN => n1749);
   U1996 : OAI22_X1 port map( A1 => n4681, A2 => n4834, B1 => n3578, B2 => 
                           n4829, ZN => n1806);
   U1997 : OAI22_X1 port map( A1 => n4684, A2 => n4834, B1 => n3579, B2 => 
                           n4830, ZN => n1807);
   U1998 : OAI22_X1 port map( A1 => n4687, A2 => n4834, B1 => n3580, B2 => 
                           n4830, ZN => n1808);
   U1999 : OAI22_X1 port map( A1 => n4690, A2 => n4834, B1 => n3581, B2 => 
                           n4830, ZN => n1809);
   U2000 : OAI22_X1 port map( A1 => n4693, A2 => n4834, B1 => n3582, B2 => 
                           n4830, ZN => n1810);
   U2001 : OAI22_X1 port map( A1 => n4696, A2 => n4834, B1 => n3583, B2 => 
                           n4830, ZN => n1811);
   U2002 : OAI22_X1 port map( A1 => n4699, A2 => n4834, B1 => n3584, B2 => 
                           n4830, ZN => n1812);
   U2003 : OAI22_X1 port map( A1 => n4702, A2 => n4834, B1 => n3585, B2 => 
                           n4830, ZN => n1813);
   U2004 : OAI22_X1 port map( A1 => n4960, A2 => n4638, B1 => n4076, B2 => 
                           n4956, ZN => n2304);
   U2005 : INV_X1 port map( A => DATAIN(9), ZN => n5162);
   U2006 : OAI22_X1 port map( A1 => n4639, A2 => n4760, B1 => n3276, B2 => 
                           n4756, ZN => n1504);
   U2007 : OAI22_X1 port map( A1 => n4639, A2 => n4808, B1 => n3468, B2 => 
                           n4804, ZN => n1696);
   U2008 : OAI22_X1 port map( A1 => n4638, A2 => n4864, B1 => n3692, B2 => 
                           n4860, ZN => n1920);
   U2009 : OAI22_X1 port map( A1 => n4638, A2 => n4888, B1 => n3788, B2 => 
                           n4884, ZN => n2016);
   U2010 : OAI22_X1 port map( A1 => n4638, A2 => n4896, B1 => n3820, B2 => 
                           n4892, ZN => n2048);
   U2011 : OAI22_X1 port map( A1 => n4638, A2 => n4920, B1 => n3916, B2 => 
                           n4916, ZN => n2144);
   U2012 : OAI22_X1 port map( A1 => n4638, A2 => n4928, B1 => n3948, B2 => 
                           n4924, ZN => n2176);
   U2013 : OAI22_X1 port map( A1 => n4638, A2 => n4952, B1 => n4044, B2 => 
                           n4948, ZN => n2272);
   U2014 : OAI22_X1 port map( A1 => n4638, A2 => n4872, B1 => n3724, B2 => 
                           n4868, ZN => n1952);
   U2015 : OAI22_X1 port map( A1 => n4638, A2 => n4880, B1 => n3756, B2 => 
                           n4876, ZN => n1984);
   U2016 : OAI22_X1 port map( A1 => n4638, A2 => n4904, B1 => n3852, B2 => 
                           n4900, ZN => n2080);
   U2017 : OAI22_X1 port map( A1 => n4638, A2 => n4912, B1 => n3884, B2 => 
                           n4908, ZN => n2112);
   U2018 : OAI22_X1 port map( A1 => n4638, A2 => n4936, B1 => n3980, B2 => 
                           n4932, ZN => n2208);
   U2019 : OAI22_X1 port map( A1 => n4638, A2 => n4944, B1 => n4012, B2 => 
                           n4940, ZN => n2240);
   U2020 : OAI22_X1 port map( A1 => n4639, A2 => n4824, B1 => n3532, B2 => 
                           n4820, ZN => n1760);
   U2021 : OAI22_X1 port map( A1 => n4639, A2 => n4856, B1 => n3660, B2 => 
                           n4852, ZN => n1888);
   U2022 : OAI22_X1 port map( A1 => n4639, A2 => n4840, B1 => n3596, B2 => 
                           n4836, ZN => n1824);
   U2023 : OAI22_X1 port map( A1 => n4639, A2 => n4848, B1 => n3628, B2 => 
                           n4844, ZN => n1856);
   U2024 : OAI22_X1 port map( A1 => n4639, A2 => n4768, B1 => n3308, B2 => 
                           n4764, ZN => n1536);
   U2025 : OAI22_X1 port map( A1 => n4639, A2 => n4776, B1 => n3340, B2 => 
                           n4772, ZN => n1568);
   U2026 : OAI22_X1 port map( A1 => n4639, A2 => n4784, B1 => n3372, B2 => 
                           n4780, ZN => n1600);
   U2027 : OAI22_X1 port map( A1 => n4639, A2 => n4792, B1 => n3404, B2 => 
                           n4788, ZN => n1632);
   U2028 : OAI22_X1 port map( A1 => n4639, A2 => n4800, B1 => n3436, B2 => 
                           n4796, ZN => n1664);
   U2029 : OAI22_X1 port map( A1 => n4639, A2 => n4816, B1 => n3500, B2 => 
                           n4812, ZN => n1728);
   U2030 : OAI22_X1 port map( A1 => n4639, A2 => n4832, B1 => n3564, B2 => 
                           n4828, ZN => n1792);
   U2031 : OAI22_X1 port map( A1 => n4622, A2 => n4736, B1 => n3174, B2 => 
                           n4732, ZN => n1402);
   U2032 : OAI22_X1 port map( A1 => n4625, A2 => n4736, B1 => n3175, B2 => 
                           n4732, ZN => n1403);
   U2033 : OAI22_X1 port map( A1 => n4628, A2 => n4736, B1 => n3176, B2 => 
                           n4732, ZN => n1404);
   U2034 : OAI22_X1 port map( A1 => n4631, A2 => n4736, B1 => n3177, B2 => 
                           n4732, ZN => n1405);
   U2035 : OAI22_X1 port map( A1 => n4634, A2 => n4736, B1 => n3178, B2 => 
                           n4732, ZN => n1406);
   U2036 : OAI22_X1 port map( A1 => n4637, A2 => n4736, B1 => n3179, B2 => 
                           n4732, ZN => n1407);
   U2037 : OAI22_X1 port map( A1 => n4706, A2 => n4738, B1 => n3202, B2 => 
                           n4734, ZN => n1430);
   U2038 : OAI22_X1 port map( A1 => n4622, A2 => n4712, B1 => n3078, B2 => 
                           n4708, ZN => n1306);
   U2039 : OAI22_X1 port map( A1 => n4625, A2 => n4712, B1 => n3079, B2 => 
                           n4708, ZN => n1307);
   U2040 : OAI22_X1 port map( A1 => n4628, A2 => n4712, B1 => n3080, B2 => 
                           n4708, ZN => n1308);
   U2041 : OAI22_X1 port map( A1 => n4631, A2 => n4712, B1 => n3081, B2 => 
                           n4708, ZN => n1309);
   U2042 : OAI22_X1 port map( A1 => n4634, A2 => n4712, B1 => n3082, B2 => 
                           n4708, ZN => n1310);
   U2043 : OAI22_X1 port map( A1 => n4637, A2 => n4712, B1 => n3083, B2 => 
                           n4708, ZN => n1311);
   U2044 : OAI22_X1 port map( A1 => n4622, A2 => n4744, B1 => n3206, B2 => 
                           n4740, ZN => n1434);
   U2045 : OAI22_X1 port map( A1 => n4625, A2 => n4744, B1 => n3207, B2 => 
                           n4740, ZN => n1435);
   U2046 : OAI22_X1 port map( A1 => n4628, A2 => n4744, B1 => n3208, B2 => 
                           n4740, ZN => n1436);
   U2047 : OAI22_X1 port map( A1 => n4631, A2 => n4744, B1 => n3209, B2 => 
                           n4740, ZN => n1437);
   U2048 : OAI22_X1 port map( A1 => n4634, A2 => n4744, B1 => n3210, B2 => 
                           n4740, ZN => n1438);
   U2049 : OAI22_X1 port map( A1 => n4637, A2 => n4744, B1 => n3211, B2 => 
                           n4740, ZN => n1439);
   U2050 : OAI22_X1 port map( A1 => n4622, A2 => n4720, B1 => n3110, B2 => 
                           n4716, ZN => n1338);
   U2051 : OAI22_X1 port map( A1 => n4625, A2 => n4720, B1 => n3111, B2 => 
                           n4716, ZN => n1339);
   U2052 : OAI22_X1 port map( A1 => n4628, A2 => n4720, B1 => n3112, B2 => 
                           n4716, ZN => n1340);
   U2053 : OAI22_X1 port map( A1 => n4631, A2 => n4720, B1 => n3113, B2 => 
                           n4716, ZN => n1341);
   U2054 : OAI22_X1 port map( A1 => n4634, A2 => n4720, B1 => n3114, B2 => 
                           n4716, ZN => n1342);
   U2055 : OAI22_X1 port map( A1 => n4637, A2 => n4720, B1 => n3115, B2 => 
                           n4716, ZN => n1343);
   U2056 : OAI22_X1 port map( A1 => n4622, A2 => n4728, B1 => n3142, B2 => 
                           n4724, ZN => n1370);
   U2057 : OAI22_X1 port map( A1 => n4625, A2 => n4728, B1 => n3143, B2 => 
                           n4724, ZN => n1371);
   U2058 : OAI22_X1 port map( A1 => n4628, A2 => n4728, B1 => n3144, B2 => 
                           n4724, ZN => n1372);
   U2059 : OAI22_X1 port map( A1 => n4631, A2 => n4728, B1 => n3145, B2 => 
                           n4724, ZN => n1373);
   U2060 : OAI22_X1 port map( A1 => n4634, A2 => n4728, B1 => n3146, B2 => 
                           n4724, ZN => n1374);
   U2061 : OAI22_X1 port map( A1 => n4637, A2 => n4728, B1 => n3147, B2 => 
                           n4724, ZN => n1375);
   U2062 : OAI22_X1 port map( A1 => n4622, A2 => n4752, B1 => n3238, B2 => 
                           n4748, ZN => n1466);
   U2063 : OAI22_X1 port map( A1 => n4625, A2 => n4752, B1 => n3239, B2 => 
                           n4748, ZN => n1467);
   U2064 : OAI22_X1 port map( A1 => n4628, A2 => n4752, B1 => n3240, B2 => 
                           n4748, ZN => n1468);
   U2065 : OAI22_X1 port map( A1 => n4631, A2 => n4752, B1 => n3241, B2 => 
                           n4748, ZN => n1469);
   U2066 : OAI22_X1 port map( A1 => n4634, A2 => n4752, B1 => n3242, B2 => 
                           n4748, ZN => n1470);
   U2067 : OAI22_X1 port map( A1 => n4637, A2 => n4752, B1 => n3243, B2 => 
                           n4748, ZN => n1471);
   U2068 : OAI22_X1 port map( A1 => n4706, A2 => n4714, B1 => n3106, B2 => 
                           n4710, ZN => n1334);
   U2069 : OAI22_X1 port map( A1 => n4706, A2 => n4746, B1 => n3234, B2 => 
                           n4742, ZN => n1462);
   U2070 : OAI22_X1 port map( A1 => n4706, A2 => n4722, B1 => n3138, B2 => 
                           n4718, ZN => n1366);
   U2071 : OAI22_X1 port map( A1 => n4706, A2 => n4730, B1 => n3170, B2 => 
                           n4726, ZN => n1398);
   U2072 : OAI22_X1 port map( A1 => n4706, A2 => n4754, B1 => n3266, B2 => 
                           n4750, ZN => n1494);
   U2073 : OAI22_X1 port map( A1 => n4613, A2 => n4736, B1 => n3171, B2 => 
                           n4732, ZN => n1399);
   U2074 : OAI22_X1 port map( A1 => n4616, A2 => n4736, B1 => n3172, B2 => 
                           n4732, ZN => n1400);
   U2075 : OAI22_X1 port map( A1 => n4619, A2 => n4736, B1 => n3173, B2 => 
                           n4732, ZN => n1401);
   U2076 : OAI22_X1 port map( A1 => n4643, A2 => n4736, B1 => n3181, B2 => 
                           n4732, ZN => n1409);
   U2077 : OAI22_X1 port map( A1 => n4646, A2 => n4737, B1 => n3182, B2 => 
                           n4732, ZN => n1410);
   U2078 : OAI22_X1 port map( A1 => n4649, A2 => n4737, B1 => n3183, B2 => 
                           n4733, ZN => n1411);
   U2079 : OAI22_X1 port map( A1 => n4652, A2 => n4737, B1 => n3184, B2 => 
                           n4733, ZN => n1412);
   U2080 : OAI22_X1 port map( A1 => n4655, A2 => n4737, B1 => n3185, B2 => 
                           n4733, ZN => n1413);
   U2081 : OAI22_X1 port map( A1 => n4658, A2 => n4737, B1 => n3186, B2 => 
                           n4733, ZN => n1414);
   U2082 : OAI22_X1 port map( A1 => n4661, A2 => n4737, B1 => n3187, B2 => 
                           n4733, ZN => n1415);
   U2083 : OAI22_X1 port map( A1 => n4664, A2 => n4737, B1 => n3188, B2 => 
                           n4733, ZN => n1416);
   U2084 : OAI22_X1 port map( A1 => n4667, A2 => n4737, B1 => n3189, B2 => 
                           n4733, ZN => n1417);
   U2085 : OAI22_X1 port map( A1 => n4670, A2 => n4737, B1 => n3190, B2 => 
                           n4733, ZN => n1418);
   U2086 : OAI22_X1 port map( A1 => n4673, A2 => n4737, B1 => n3191, B2 => 
                           n4733, ZN => n1419);
   U2087 : OAI22_X1 port map( A1 => n4676, A2 => n4737, B1 => n3192, B2 => 
                           n4733, ZN => n1420);
   U2088 : OAI22_X1 port map( A1 => n4679, A2 => n4737, B1 => n3193, B2 => 
                           n4733, ZN => n1421);
   U2089 : OAI22_X1 port map( A1 => n4682, A2 => n4738, B1 => n3194, B2 => 
                           n4733, ZN => n1422);
   U2090 : OAI22_X1 port map( A1 => n4685, A2 => n4738, B1 => n3195, B2 => 
                           n4734, ZN => n1423);
   U2091 : OAI22_X1 port map( A1 => n4688, A2 => n4738, B1 => n3196, B2 => 
                           n4734, ZN => n1424);
   U2092 : OAI22_X1 port map( A1 => n4691, A2 => n4738, B1 => n3197, B2 => 
                           n4734, ZN => n1425);
   U2093 : OAI22_X1 port map( A1 => n4694, A2 => n4738, B1 => n3198, B2 => 
                           n4734, ZN => n1426);
   U2094 : OAI22_X1 port map( A1 => n4697, A2 => n4738, B1 => n3199, B2 => 
                           n4734, ZN => n1427);
   U2095 : OAI22_X1 port map( A1 => n4700, A2 => n4738, B1 => n3200, B2 => 
                           n4734, ZN => n1428);
   U2096 : OAI22_X1 port map( A1 => n4703, A2 => n4738, B1 => n3201, B2 => 
                           n4734, ZN => n1429);
   U2097 : OAI22_X1 port map( A1 => n4613, A2 => n4712, B1 => n3075, B2 => 
                           n4708, ZN => n1303);
   U2098 : OAI22_X1 port map( A1 => n4616, A2 => n4712, B1 => n3076, B2 => 
                           n4708, ZN => n1304);
   U2099 : OAI22_X1 port map( A1 => n4619, A2 => n4712, B1 => n3077, B2 => 
                           n4708, ZN => n1305);
   U2100 : OAI22_X1 port map( A1 => n4643, A2 => n4712, B1 => n3085, B2 => 
                           n4708, ZN => n1313);
   U2101 : OAI22_X1 port map( A1 => n4646, A2 => n4713, B1 => n3086, B2 => 
                           n4708, ZN => n1314);
   U2102 : OAI22_X1 port map( A1 => n4649, A2 => n4713, B1 => n3087, B2 => 
                           n4709, ZN => n1315);
   U2103 : OAI22_X1 port map( A1 => n4652, A2 => n4713, B1 => n3088, B2 => 
                           n4709, ZN => n1316);
   U2104 : OAI22_X1 port map( A1 => n4655, A2 => n4713, B1 => n3089, B2 => 
                           n4709, ZN => n1317);
   U2105 : OAI22_X1 port map( A1 => n4658, A2 => n4713, B1 => n3090, B2 => 
                           n4709, ZN => n1318);
   U2106 : OAI22_X1 port map( A1 => n4661, A2 => n4713, B1 => n3091, B2 => 
                           n4709, ZN => n1319);
   U2107 : OAI22_X1 port map( A1 => n4664, A2 => n4713, B1 => n3092, B2 => 
                           n4709, ZN => n1320);
   U2108 : OAI22_X1 port map( A1 => n4667, A2 => n4713, B1 => n3093, B2 => 
                           n4709, ZN => n1321);
   U2109 : OAI22_X1 port map( A1 => n4670, A2 => n4713, B1 => n3094, B2 => 
                           n4709, ZN => n1322);
   U2110 : OAI22_X1 port map( A1 => n4673, A2 => n4713, B1 => n3095, B2 => 
                           n4709, ZN => n1323);
   U2111 : OAI22_X1 port map( A1 => n4676, A2 => n4713, B1 => n3096, B2 => 
                           n4709, ZN => n1324);
   U2112 : OAI22_X1 port map( A1 => n4679, A2 => n4713, B1 => n3097, B2 => 
                           n4709, ZN => n1325);
   U2113 : OAI22_X1 port map( A1 => n4613, A2 => n4744, B1 => n3203, B2 => 
                           n4740, ZN => n1431);
   U2114 : OAI22_X1 port map( A1 => n4616, A2 => n4744, B1 => n3204, B2 => 
                           n4740, ZN => n1432);
   U2115 : OAI22_X1 port map( A1 => n4619, A2 => n4744, B1 => n3205, B2 => 
                           n4740, ZN => n1433);
   U2116 : OAI22_X1 port map( A1 => n4643, A2 => n4744, B1 => n3213, B2 => 
                           n4740, ZN => n1441);
   U2117 : OAI22_X1 port map( A1 => n4646, A2 => n4745, B1 => n3214, B2 => 
                           n4740, ZN => n1442);
   U2118 : OAI22_X1 port map( A1 => n4649, A2 => n4745, B1 => n3215, B2 => 
                           n4741, ZN => n1443);
   U2119 : OAI22_X1 port map( A1 => n4652, A2 => n4745, B1 => n3216, B2 => 
                           n4741, ZN => n1444);
   U2120 : OAI22_X1 port map( A1 => n4655, A2 => n4745, B1 => n3217, B2 => 
                           n4741, ZN => n1445);
   U2121 : OAI22_X1 port map( A1 => n4658, A2 => n4745, B1 => n3218, B2 => 
                           n4741, ZN => n1446);
   U2122 : OAI22_X1 port map( A1 => n4661, A2 => n4745, B1 => n3219, B2 => 
                           n4741, ZN => n1447);
   U2123 : OAI22_X1 port map( A1 => n4664, A2 => n4745, B1 => n3220, B2 => 
                           n4741, ZN => n1448);
   U2124 : OAI22_X1 port map( A1 => n4667, A2 => n4745, B1 => n3221, B2 => 
                           n4741, ZN => n1449);
   U2125 : OAI22_X1 port map( A1 => n4670, A2 => n4745, B1 => n3222, B2 => 
                           n4741, ZN => n1450);
   U2126 : OAI22_X1 port map( A1 => n4673, A2 => n4745, B1 => n3223, B2 => 
                           n4741, ZN => n1451);
   U2127 : OAI22_X1 port map( A1 => n4676, A2 => n4745, B1 => n3224, B2 => 
                           n4741, ZN => n1452);
   U2128 : OAI22_X1 port map( A1 => n4679, A2 => n4745, B1 => n3225, B2 => 
                           n4741, ZN => n1453);
   U2129 : OAI22_X1 port map( A1 => n4613, A2 => n4720, B1 => n3107, B2 => 
                           n4716, ZN => n1335);
   U2130 : OAI22_X1 port map( A1 => n4616, A2 => n4720, B1 => n3108, B2 => 
                           n4716, ZN => n1336);
   U2131 : OAI22_X1 port map( A1 => n4619, A2 => n4720, B1 => n3109, B2 => 
                           n4716, ZN => n1337);
   U2132 : OAI22_X1 port map( A1 => n4643, A2 => n4720, B1 => n3117, B2 => 
                           n4716, ZN => n1345);
   U2133 : OAI22_X1 port map( A1 => n4646, A2 => n4721, B1 => n3118, B2 => 
                           n4716, ZN => n1346);
   U2134 : OAI22_X1 port map( A1 => n4649, A2 => n4721, B1 => n3119, B2 => 
                           n4717, ZN => n1347);
   U2135 : OAI22_X1 port map( A1 => n4652, A2 => n4721, B1 => n3120, B2 => 
                           n4717, ZN => n1348);
   U2136 : OAI22_X1 port map( A1 => n4655, A2 => n4721, B1 => n3121, B2 => 
                           n4717, ZN => n1349);
   U2137 : OAI22_X1 port map( A1 => n4658, A2 => n4721, B1 => n3122, B2 => 
                           n4717, ZN => n1350);
   U2138 : OAI22_X1 port map( A1 => n4661, A2 => n4721, B1 => n3123, B2 => 
                           n4717, ZN => n1351);
   U2139 : OAI22_X1 port map( A1 => n4664, A2 => n4721, B1 => n3124, B2 => 
                           n4717, ZN => n1352);
   U2140 : OAI22_X1 port map( A1 => n4667, A2 => n4721, B1 => n3125, B2 => 
                           n4717, ZN => n1353);
   U2141 : OAI22_X1 port map( A1 => n4670, A2 => n4721, B1 => n3126, B2 => 
                           n4717, ZN => n1354);
   U2142 : OAI22_X1 port map( A1 => n4673, A2 => n4721, B1 => n3127, B2 => 
                           n4717, ZN => n1355);
   U2143 : OAI22_X1 port map( A1 => n4676, A2 => n4721, B1 => n3128, B2 => 
                           n4717, ZN => n1356);
   U2144 : OAI22_X1 port map( A1 => n4679, A2 => n4721, B1 => n3129, B2 => 
                           n4717, ZN => n1357);
   U2145 : OAI22_X1 port map( A1 => n4613, A2 => n4728, B1 => n3139, B2 => 
                           n4724, ZN => n1367);
   U2146 : OAI22_X1 port map( A1 => n4616, A2 => n4728, B1 => n3140, B2 => 
                           n4724, ZN => n1368);
   U2147 : OAI22_X1 port map( A1 => n4619, A2 => n4728, B1 => n3141, B2 => 
                           n4724, ZN => n1369);
   U2148 : OAI22_X1 port map( A1 => n4643, A2 => n4728, B1 => n3149, B2 => 
                           n4724, ZN => n1377);
   U2149 : OAI22_X1 port map( A1 => n4646, A2 => n4729, B1 => n3150, B2 => 
                           n4724, ZN => n1378);
   U2150 : OAI22_X1 port map( A1 => n4649, A2 => n4729, B1 => n3151, B2 => 
                           n4725, ZN => n1379);
   U2151 : OAI22_X1 port map( A1 => n4652, A2 => n4729, B1 => n3152, B2 => 
                           n4725, ZN => n1380);
   U2152 : OAI22_X1 port map( A1 => n4655, A2 => n4729, B1 => n3153, B2 => 
                           n4725, ZN => n1381);
   U2153 : OAI22_X1 port map( A1 => n4658, A2 => n4729, B1 => n3154, B2 => 
                           n4725, ZN => n1382);
   U2154 : OAI22_X1 port map( A1 => n4661, A2 => n4729, B1 => n3155, B2 => 
                           n4725, ZN => n1383);
   U2155 : OAI22_X1 port map( A1 => n4664, A2 => n4729, B1 => n3156, B2 => 
                           n4725, ZN => n1384);
   U2156 : OAI22_X1 port map( A1 => n4667, A2 => n4729, B1 => n3157, B2 => 
                           n4725, ZN => n1385);
   U2157 : OAI22_X1 port map( A1 => n4670, A2 => n4729, B1 => n3158, B2 => 
                           n4725, ZN => n1386);
   U2158 : OAI22_X1 port map( A1 => n4673, A2 => n4729, B1 => n3159, B2 => 
                           n4725, ZN => n1387);
   U2159 : OAI22_X1 port map( A1 => n4676, A2 => n4729, B1 => n3160, B2 => 
                           n4725, ZN => n1388);
   U2160 : OAI22_X1 port map( A1 => n4679, A2 => n4729, B1 => n3161, B2 => 
                           n4725, ZN => n1389);
   U2161 : OAI22_X1 port map( A1 => n4613, A2 => n4752, B1 => n3235, B2 => 
                           n4748, ZN => n1463);
   U2162 : OAI22_X1 port map( A1 => n4616, A2 => n4752, B1 => n3236, B2 => 
                           n4748, ZN => n1464);
   U2163 : OAI22_X1 port map( A1 => n4619, A2 => n4752, B1 => n3237, B2 => 
                           n4748, ZN => n1465);
   U2164 : OAI22_X1 port map( A1 => n4643, A2 => n4752, B1 => n3245, B2 => 
                           n4748, ZN => n1473);
   U2165 : OAI22_X1 port map( A1 => n4646, A2 => n4753, B1 => n3246, B2 => 
                           n4748, ZN => n1474);
   U2166 : OAI22_X1 port map( A1 => n4649, A2 => n4753, B1 => n3247, B2 => 
                           n4749, ZN => n1475);
   U2167 : OAI22_X1 port map( A1 => n4652, A2 => n4753, B1 => n3248, B2 => 
                           n4749, ZN => n1476);
   U2168 : OAI22_X1 port map( A1 => n4655, A2 => n4753, B1 => n3249, B2 => 
                           n4749, ZN => n1477);
   U2169 : OAI22_X1 port map( A1 => n4658, A2 => n4753, B1 => n3250, B2 => 
                           n4749, ZN => n1478);
   U2170 : OAI22_X1 port map( A1 => n4661, A2 => n4753, B1 => n3251, B2 => 
                           n4749, ZN => n1479);
   U2171 : OAI22_X1 port map( A1 => n4664, A2 => n4753, B1 => n3252, B2 => 
                           n4749, ZN => n1480);
   U2172 : OAI22_X1 port map( A1 => n4667, A2 => n4753, B1 => n3253, B2 => 
                           n4749, ZN => n1481);
   U2173 : OAI22_X1 port map( A1 => n4670, A2 => n4753, B1 => n3254, B2 => 
                           n4749, ZN => n1482);
   U2174 : OAI22_X1 port map( A1 => n4673, A2 => n4753, B1 => n3255, B2 => 
                           n4749, ZN => n1483);
   U2175 : OAI22_X1 port map( A1 => n4676, A2 => n4753, B1 => n3256, B2 => 
                           n4749, ZN => n1484);
   U2176 : OAI22_X1 port map( A1 => n4679, A2 => n4753, B1 => n3257, B2 => 
                           n4749, ZN => n1485);
   U2177 : OAI22_X1 port map( A1 => n4682, A2 => n4714, B1 => n3098, B2 => 
                           n4709, ZN => n1326);
   U2178 : OAI22_X1 port map( A1 => n4685, A2 => n4714, B1 => n3099, B2 => 
                           n4710, ZN => n1327);
   U2179 : OAI22_X1 port map( A1 => n4688, A2 => n4714, B1 => n3100, B2 => 
                           n4710, ZN => n1328);
   U2180 : OAI22_X1 port map( A1 => n4691, A2 => n4714, B1 => n3101, B2 => 
                           n4710, ZN => n1329);
   U2181 : OAI22_X1 port map( A1 => n4694, A2 => n4714, B1 => n3102, B2 => 
                           n4710, ZN => n1330);
   U2182 : OAI22_X1 port map( A1 => n4697, A2 => n4714, B1 => n3103, B2 => 
                           n4710, ZN => n1331);
   U2183 : OAI22_X1 port map( A1 => n4700, A2 => n4714, B1 => n3104, B2 => 
                           n4710, ZN => n1332);
   U2184 : OAI22_X1 port map( A1 => n4703, A2 => n4714, B1 => n3105, B2 => 
                           n4710, ZN => n1333);
   U2185 : OAI22_X1 port map( A1 => n4682, A2 => n4746, B1 => n3226, B2 => 
                           n4741, ZN => n1454);
   U2186 : OAI22_X1 port map( A1 => n4685, A2 => n4746, B1 => n3227, B2 => 
                           n4742, ZN => n1455);
   U2187 : OAI22_X1 port map( A1 => n4688, A2 => n4746, B1 => n3228, B2 => 
                           n4742, ZN => n1456);
   U2188 : OAI22_X1 port map( A1 => n4691, A2 => n4746, B1 => n3229, B2 => 
                           n4742, ZN => n1457);
   U2189 : OAI22_X1 port map( A1 => n4694, A2 => n4746, B1 => n3230, B2 => 
                           n4742, ZN => n1458);
   U2190 : OAI22_X1 port map( A1 => n4697, A2 => n4746, B1 => n3231, B2 => 
                           n4742, ZN => n1459);
   U2191 : OAI22_X1 port map( A1 => n4700, A2 => n4746, B1 => n3232, B2 => 
                           n4742, ZN => n1460);
   U2192 : OAI22_X1 port map( A1 => n4703, A2 => n4746, B1 => n3233, B2 => 
                           n4742, ZN => n1461);
   U2193 : OAI22_X1 port map( A1 => n4682, A2 => n4722, B1 => n3130, B2 => 
                           n4717, ZN => n1358);
   U2194 : OAI22_X1 port map( A1 => n4685, A2 => n4722, B1 => n3131, B2 => 
                           n4718, ZN => n1359);
   U2195 : OAI22_X1 port map( A1 => n4688, A2 => n4722, B1 => n3132, B2 => 
                           n4718, ZN => n1360);
   U2196 : OAI22_X1 port map( A1 => n4691, A2 => n4722, B1 => n3133, B2 => 
                           n4718, ZN => n1361);
   U2197 : OAI22_X1 port map( A1 => n4694, A2 => n4722, B1 => n3134, B2 => 
                           n4718, ZN => n1362);
   U2198 : OAI22_X1 port map( A1 => n4697, A2 => n4722, B1 => n3135, B2 => 
                           n4718, ZN => n1363);
   U2199 : OAI22_X1 port map( A1 => n4700, A2 => n4722, B1 => n3136, B2 => 
                           n4718, ZN => n1364);
   U2200 : OAI22_X1 port map( A1 => n4703, A2 => n4722, B1 => n3137, B2 => 
                           n4718, ZN => n1365);
   U2201 : OAI22_X1 port map( A1 => n4682, A2 => n4730, B1 => n3162, B2 => 
                           n4725, ZN => n1390);
   U2202 : OAI22_X1 port map( A1 => n4685, A2 => n4730, B1 => n3163, B2 => 
                           n4726, ZN => n1391);
   U2203 : OAI22_X1 port map( A1 => n4688, A2 => n4730, B1 => n3164, B2 => 
                           n4726, ZN => n1392);
   U2204 : OAI22_X1 port map( A1 => n4691, A2 => n4730, B1 => n3165, B2 => 
                           n4726, ZN => n1393);
   U2205 : OAI22_X1 port map( A1 => n4694, A2 => n4730, B1 => n3166, B2 => 
                           n4726, ZN => n1394);
   U2206 : OAI22_X1 port map( A1 => n4697, A2 => n4730, B1 => n3167, B2 => 
                           n4726, ZN => n1395);
   U2207 : OAI22_X1 port map( A1 => n4700, A2 => n4730, B1 => n3168, B2 => 
                           n4726, ZN => n1396);
   U2208 : OAI22_X1 port map( A1 => n4703, A2 => n4730, B1 => n3169, B2 => 
                           n4726, ZN => n1397);
   U2209 : OAI22_X1 port map( A1 => n4682, A2 => n4754, B1 => n3258, B2 => 
                           n4749, ZN => n1486);
   U2210 : OAI22_X1 port map( A1 => n4685, A2 => n4754, B1 => n3259, B2 => 
                           n4750, ZN => n1487);
   U2211 : OAI22_X1 port map( A1 => n4688, A2 => n4754, B1 => n3260, B2 => 
                           n4750, ZN => n1488);
   U2212 : OAI22_X1 port map( A1 => n4691, A2 => n4754, B1 => n3261, B2 => 
                           n4750, ZN => n1489);
   U2213 : OAI22_X1 port map( A1 => n4694, A2 => n4754, B1 => n3262, B2 => 
                           n4750, ZN => n1490);
   U2214 : OAI22_X1 port map( A1 => n4697, A2 => n4754, B1 => n3263, B2 => 
                           n4750, ZN => n1491);
   U2215 : OAI22_X1 port map( A1 => n4700, A2 => n4754, B1 => n3264, B2 => 
                           n4750, ZN => n1492);
   U2216 : OAI22_X1 port map( A1 => n4703, A2 => n4754, B1 => n3265, B2 => 
                           n4750, ZN => n1493);
   U2217 : OAI22_X1 port map( A1 => n4640, A2 => n4736, B1 => n3180, B2 => 
                           n4732, ZN => n1408);
   U2218 : OAI22_X1 port map( A1 => n4640, A2 => n4712, B1 => n3084, B2 => 
                           n4708, ZN => n1312);
   U2219 : OAI22_X1 port map( A1 => n4640, A2 => n4744, B1 => n3212, B2 => 
                           n4740, ZN => n1440);
   U2220 : OAI22_X1 port map( A1 => n4640, A2 => n4720, B1 => n3116, B2 => 
                           n4716, ZN => n1344);
   U2221 : OAI22_X1 port map( A1 => n4640, A2 => n4728, B1 => n3148, B2 => 
                           n4724, ZN => n1376);
   U2222 : OAI22_X1 port map( A1 => n4640, A2 => n4752, B1 => n3244, B2 => 
                           n4748, ZN => n1472);
   U2223 : NOR3_X1 port map( A1 => n5137, A2 => ADD_RD2(1), A3 => n5131, ZN => 
                           n2664);
   U2224 : OAI22_X1 port map( A1 => n3043, A2 => n5040, B1 => n2655, B2 => 
                           n5036, ZN => n4099);
   U2225 : NOR4_X1 port map( A1 => n2656, A2 => n2657, A3 => n2658, A4 => n2659
                           , ZN => n2655);
   U2226 : OAI221_X1 port map( B1 => n3267, B2 => n4996, C1 => n3075, C2 => 
                           n4992, A => n2681, ZN => n2657);
   U2227 : OAI221_X1 port map( B1 => n3171, B2 => n4980, C1 => n3203, C2 => 
                           n4976, A => n2683, ZN => n2656);
   U2228 : OAI22_X1 port map( A1 => n3044, A2 => n5040, B1 => n2636, B2 => 
                           n5036, ZN => n4100);
   U2229 : NOR4_X1 port map( A1 => n2637, A2 => n2638, A3 => n2639, A4 => n2640
                           , ZN => n2636);
   U2230 : OAI221_X1 port map( B1 => n3268, B2 => n4996, C1 => n3076, C2 => 
                           n4992, A => n2653, ZN => n2638);
   U2231 : OAI221_X1 port map( B1 => n3172, B2 => n4980, C1 => n3204, C2 => 
                           n4976, A => n2654, ZN => n2637);
   U2232 : OAI22_X1 port map( A1 => n3045, A2 => n5040, B1 => n2617, B2 => 
                           n5036, ZN => n4101);
   U2233 : NOR4_X1 port map( A1 => n2618, A2 => n2619, A3 => n2620, A4 => n2621
                           , ZN => n2617);
   U2234 : OAI221_X1 port map( B1 => n3269, B2 => n4996, C1 => n3077, C2 => 
                           n4992, A => n2634, ZN => n2619);
   U2235 : OAI221_X1 port map( B1 => n3173, B2 => n4980, C1 => n3205, C2 => 
                           n4976, A => n2635, ZN => n2618);
   U2236 : OAI22_X1 port map( A1 => n3046, A2 => n5040, B1 => n2598, B2 => 
                           n5036, ZN => n4102);
   U2237 : NOR4_X1 port map( A1 => n2599, A2 => n2600, A3 => n2601, A4 => n2602
                           , ZN => n2598);
   U2238 : OAI221_X1 port map( B1 => n3270, B2 => n4996, C1 => n3078, C2 => 
                           n4992, A => n2615, ZN => n2600);
   U2239 : OAI221_X1 port map( B1 => n3174, B2 => n4980, C1 => n3206, C2 => 
                           n4976, A => n2616, ZN => n2599);
   U2240 : OAI22_X1 port map( A1 => n3047, A2 => n5040, B1 => n2579, B2 => 
                           n5036, ZN => n4103);
   U2241 : NOR4_X1 port map( A1 => n2580, A2 => n2581, A3 => n2582, A4 => n2583
                           , ZN => n2579);
   U2242 : OAI221_X1 port map( B1 => n3271, B2 => n4996, C1 => n3079, C2 => 
                           n4992, A => n2596, ZN => n2581);
   U2243 : OAI221_X1 port map( B1 => n3175, B2 => n4980, C1 => n3207, C2 => 
                           n4976, A => n2597, ZN => n2580);
   U2244 : OAI22_X1 port map( A1 => n3048, A2 => n5040, B1 => n2560, B2 => 
                           n5036, ZN => n4104);
   U2245 : NOR4_X1 port map( A1 => n2561, A2 => n2562, A3 => n2563, A4 => n2564
                           , ZN => n2560);
   U2246 : OAI221_X1 port map( B1 => n3272, B2 => n4996, C1 => n3080, C2 => 
                           n4992, A => n2577, ZN => n2562);
   U2247 : OAI221_X1 port map( B1 => n3176, B2 => n4980, C1 => n3208, C2 => 
                           n4976, A => n2578, ZN => n2561);
   U2248 : OAI22_X1 port map( A1 => n3049, A2 => n5040, B1 => n2541, B2 => 
                           n5036, ZN => n4105);
   U2249 : NOR4_X1 port map( A1 => n2542, A2 => n2543, A3 => n2544, A4 => n2545
                           , ZN => n2541);
   U2250 : OAI221_X1 port map( B1 => n3273, B2 => n4996, C1 => n3081, C2 => 
                           n4992, A => n2558, ZN => n2543);
   U2251 : OAI221_X1 port map( B1 => n3177, B2 => n4980, C1 => n3209, C2 => 
                           n4976, A => n2559, ZN => n2542);
   U2252 : OAI22_X1 port map( A1 => n3050, A2 => n5040, B1 => n2522, B2 => 
                           n5036, ZN => n4106);
   U2253 : NOR4_X1 port map( A1 => n2523, A2 => n2524, A3 => n2525, A4 => n2526
                           , ZN => n2522);
   U2254 : OAI221_X1 port map( B1 => n3274, B2 => n4996, C1 => n3082, C2 => 
                           n4992, A => n2539, ZN => n2524);
   U2255 : OAI221_X1 port map( B1 => n3178, B2 => n4980, C1 => n3210, C2 => 
                           n4976, A => n2540, ZN => n2523);
   U2256 : OAI22_X1 port map( A1 => n3051, A2 => n5040, B1 => n2503, B2 => 
                           n5036, ZN => n4107);
   U2257 : NOR4_X1 port map( A1 => n2504, A2 => n2505, A3 => n2506, A4 => n2507
                           , ZN => n2503);
   U2258 : OAI221_X1 port map( B1 => n3275, B2 => n4996, C1 => n3083, C2 => 
                           n4992, A => n2520, ZN => n2505);
   U2259 : OAI221_X1 port map( B1 => n3179, B2 => n4980, C1 => n3211, C2 => 
                           n4976, A => n2521, ZN => n2504);
   U2260 : OAI22_X1 port map( A1 => n3052, A2 => n5040, B1 => n2484, B2 => 
                           n5036, ZN => n4108);
   U2261 : NOR4_X1 port map( A1 => n2485, A2 => n2486, A3 => n2487, A4 => n2488
                           , ZN => n2484);
   U2262 : OAI221_X1 port map( B1 => n3276, B2 => n4996, C1 => n3084, C2 => 
                           n4992, A => n2501, ZN => n2486);
   U2263 : OAI221_X1 port map( B1 => n3180, B2 => n4980, C1 => n3212, C2 => 
                           n4976, A => n2502, ZN => n2485);
   U2264 : OAI22_X1 port map( A1 => n3053, A2 => n5040, B1 => n2465, B2 => 
                           n5036, ZN => n4109);
   U2265 : NOR4_X1 port map( A1 => n2466, A2 => n2467, A3 => n2468, A4 => n2469
                           , ZN => n2465);
   U2266 : OAI221_X1 port map( B1 => n3277, B2 => n4996, C1 => n3085, C2 => 
                           n4992, A => n2482, ZN => n2467);
   U2267 : OAI221_X1 port map( B1 => n3181, B2 => n4980, C1 => n3213, C2 => 
                           n4976, A => n2483, ZN => n2466);
   U2268 : OAI22_X1 port map( A1 => n3054, A2 => n5040, B1 => n2446, B2 => 
                           n5037, ZN => n4110);
   U2269 : NOR4_X1 port map( A1 => n2447, A2 => n2448, A3 => n2449, A4 => n2450
                           , ZN => n2446);
   U2270 : OAI221_X1 port map( B1 => n3278, B2 => n4996, C1 => n3086, C2 => 
                           n4992, A => n2463, ZN => n2448);
   U2271 : OAI221_X1 port map( B1 => n3182, B2 => n4980, C1 => n3214, C2 => 
                           n4976, A => n2464, ZN => n2447);
   U2272 : OAI22_X1 port map( A1 => n3055, A2 => n5041, B1 => n2427, B2 => 
                           n5037, ZN => n4111);
   U2273 : NOR4_X1 port map( A1 => n2428, A2 => n2429, A3 => n2430, A4 => n2431
                           , ZN => n2427);
   U2274 : OAI221_X1 port map( B1 => n3279, B2 => n4997, C1 => n3087, C2 => 
                           n4993, A => n2444, ZN => n2429);
   U2275 : OAI221_X1 port map( B1 => n3183, B2 => n4981, C1 => n3215, C2 => 
                           n4977, A => n2445, ZN => n2428);
   U2276 : OAI22_X1 port map( A1 => n3056, A2 => n5041, B1 => n2408, B2 => 
                           n5037, ZN => n4112);
   U2277 : NOR4_X1 port map( A1 => n2409, A2 => n2410, A3 => n2411, A4 => n2412
                           , ZN => n2408);
   U2278 : OAI221_X1 port map( B1 => n3280, B2 => n4997, C1 => n3088, C2 => 
                           n4993, A => n2425, ZN => n2410);
   U2279 : OAI221_X1 port map( B1 => n3184, B2 => n4981, C1 => n3216, C2 => 
                           n4977, A => n2426, ZN => n2409);
   U2280 : OAI22_X1 port map( A1 => n3057, A2 => n5041, B1 => n2389, B2 => 
                           n5037, ZN => n4113);
   U2281 : NOR4_X1 port map( A1 => n2390, A2 => n2391, A3 => n2392, A4 => n2393
                           , ZN => n2389);
   U2282 : OAI221_X1 port map( B1 => n3281, B2 => n4997, C1 => n3089, C2 => 
                           n4993, A => n2406, ZN => n2391);
   U2283 : OAI221_X1 port map( B1 => n3185, B2 => n4981, C1 => n3217, C2 => 
                           n4977, A => n2407, ZN => n2390);
   U2284 : OAI22_X1 port map( A1 => n3058, A2 => n5041, B1 => n2370, B2 => 
                           n5037, ZN => n4114);
   U2285 : NOR4_X1 port map( A1 => n2371, A2 => n2372, A3 => n2373, A4 => n2374
                           , ZN => n2370);
   U2286 : OAI221_X1 port map( B1 => n3282, B2 => n4997, C1 => n3090, C2 => 
                           n4993, A => n2387, ZN => n2372);
   U2287 : OAI221_X1 port map( B1 => n3186, B2 => n4981, C1 => n3218, C2 => 
                           n4977, A => n2388, ZN => n2371);
   U2288 : OAI22_X1 port map( A1 => n3059, A2 => n5041, B1 => n2351, B2 => 
                           n5037, ZN => n4115);
   U2289 : NOR4_X1 port map( A1 => n2352, A2 => n2353, A3 => n2354, A4 => n2355
                           , ZN => n2351);
   U2290 : OAI221_X1 port map( B1 => n3283, B2 => n4997, C1 => n3091, C2 => 
                           n4993, A => n2368, ZN => n2353);
   U2291 : OAI221_X1 port map( B1 => n3187, B2 => n4981, C1 => n3219, C2 => 
                           n4977, A => n2369, ZN => n2352);
   U2292 : OAI22_X1 port map( A1 => n3060, A2 => n5041, B1 => n2332, B2 => 
                           n5037, ZN => n4116);
   U2293 : NOR4_X1 port map( A1 => n2333, A2 => n2334, A3 => n2335, A4 => n2336
                           , ZN => n2332);
   U2294 : OAI221_X1 port map( B1 => n3284, B2 => n4997, C1 => n3092, C2 => 
                           n4993, A => n2349, ZN => n2334);
   U2295 : OAI221_X1 port map( B1 => n3188, B2 => n4981, C1 => n3220, C2 => 
                           n4977, A => n2350, ZN => n2333);
   U2296 : OAI22_X1 port map( A1 => n3061, A2 => n5041, B1 => n1289, B2 => 
                           n5037, ZN => n4117);
   U2297 : NOR4_X1 port map( A1 => n1290, A2 => n1291, A3 => n1292, A4 => n1293
                           , ZN => n1289);
   U2298 : OAI221_X1 port map( B1 => n3285, B2 => n4997, C1 => n3093, C2 => 
                           n4993, A => n2330, ZN => n1291);
   U2299 : OAI221_X1 port map( B1 => n3189, B2 => n4981, C1 => n3221, C2 => 
                           n4977, A => n2331, ZN => n1290);
   U2300 : OAI22_X1 port map( A1 => n3062, A2 => n5041, B1 => n1270, B2 => 
                           n5037, ZN => n4118);
   U2301 : NOR4_X1 port map( A1 => n1271, A2 => n1272, A3 => n1273, A4 => n1274
                           , ZN => n1270);
   U2302 : OAI221_X1 port map( B1 => n3286, B2 => n4997, C1 => n3094, C2 => 
                           n4993, A => n1287, ZN => n1272);
   U2303 : OAI221_X1 port map( B1 => n3190, B2 => n4981, C1 => n3222, C2 => 
                           n4977, A => n1288, ZN => n1271);
   U2304 : OAI22_X1 port map( A1 => n3063, A2 => n5041, B1 => n1251, B2 => 
                           n5037, ZN => n4119);
   U2305 : NOR4_X1 port map( A1 => n1252, A2 => n1253, A3 => n1254, A4 => n1255
                           , ZN => n1251);
   U2306 : OAI221_X1 port map( B1 => n3287, B2 => n4997, C1 => n3095, C2 => 
                           n4993, A => n1268, ZN => n1253);
   U2307 : OAI221_X1 port map( B1 => n3191, B2 => n4981, C1 => n3223, C2 => 
                           n4977, A => n1269, ZN => n1252);
   U2308 : OAI22_X1 port map( A1 => n3064, A2 => n5041, B1 => n1232, B2 => 
                           n5037, ZN => n4120);
   U2309 : NOR4_X1 port map( A1 => n1233, A2 => n1234, A3 => n1235, A4 => n1236
                           , ZN => n1232);
   U2310 : OAI221_X1 port map( B1 => n3288, B2 => n4997, C1 => n3096, C2 => 
                           n4993, A => n1249, ZN => n1234);
   U2311 : OAI221_X1 port map( B1 => n3192, B2 => n4981, C1 => n3224, C2 => 
                           n4977, A => n1250, ZN => n1233);
   U2312 : OAI22_X1 port map( A1 => n3065, A2 => n5041, B1 => n1213, B2 => 
                           n5037, ZN => n4121);
   U2313 : NOR4_X1 port map( A1 => n1214, A2 => n1215, A3 => n1216, A4 => n1217
                           , ZN => n1213);
   U2314 : OAI221_X1 port map( B1 => n3289, B2 => n4997, C1 => n3097, C2 => 
                           n4993, A => n1230, ZN => n1215);
   U2315 : OAI221_X1 port map( B1 => n3193, B2 => n4981, C1 => n3225, C2 => 
                           n4977, A => n1231, ZN => n1214);
   U2316 : OAI22_X1 port map( A1 => n3066, A2 => n5041, B1 => n1194, B2 => 
                           n5038, ZN => n4122);
   U2317 : NOR4_X1 port map( A1 => n1195, A2 => n1196, A3 => n1197, A4 => n1198
                           , ZN => n1194);
   U2318 : OAI221_X1 port map( B1 => n3290, B2 => n4997, C1 => n3098, C2 => 
                           n4993, A => n1211, ZN => n1196);
   U2319 : OAI221_X1 port map( B1 => n3194, B2 => n4981, C1 => n3226, C2 => 
                           n4977, A => n1212, ZN => n1195);
   U2320 : OAI22_X1 port map( A1 => n3067, A2 => n5042, B1 => n1175, B2 => 
                           n5038, ZN => n4123);
   U2321 : NOR4_X1 port map( A1 => n1176, A2 => n1177, A3 => n1178, A4 => n1179
                           , ZN => n1175);
   U2322 : OAI221_X1 port map( B1 => n3291, B2 => n4998, C1 => n3099, C2 => 
                           n4994, A => n1192, ZN => n1177);
   U2323 : OAI221_X1 port map( B1 => n3195, B2 => n4982, C1 => n3227, C2 => 
                           n4978, A => n1193, ZN => n1176);
   U2324 : OAI22_X1 port map( A1 => n3068, A2 => n5042, B1 => n1156, B2 => 
                           n5038, ZN => n4124);
   U2325 : NOR4_X1 port map( A1 => n1157, A2 => n1158, A3 => n1159, A4 => n1160
                           , ZN => n1156);
   U2326 : OAI221_X1 port map( B1 => n3292, B2 => n4998, C1 => n3100, C2 => 
                           n4994, A => n1173, ZN => n1158);
   U2327 : OAI221_X1 port map( B1 => n3196, B2 => n4982, C1 => n3228, C2 => 
                           n4978, A => n1174, ZN => n1157);
   U2328 : OAI22_X1 port map( A1 => n3069, A2 => n5042, B1 => n1137, B2 => 
                           n5038, ZN => n4125);
   U2329 : NOR4_X1 port map( A1 => n1138, A2 => n1139, A3 => n1140, A4 => n1141
                           , ZN => n1137);
   U2330 : OAI221_X1 port map( B1 => n3293, B2 => n4998, C1 => n3101, C2 => 
                           n4994, A => n1154, ZN => n1139);
   U2331 : OAI221_X1 port map( B1 => n3197, B2 => n4982, C1 => n3229, C2 => 
                           n4978, A => n1155, ZN => n1138);
   U2332 : OAI22_X1 port map( A1 => n3070, A2 => n5042, B1 => n1118, B2 => 
                           n5038, ZN => n4126);
   U2333 : NOR4_X1 port map( A1 => n1119, A2 => n1120, A3 => n1121, A4 => n1122
                           , ZN => n1118);
   U2334 : OAI221_X1 port map( B1 => n3294, B2 => n4998, C1 => n3102, C2 => 
                           n4994, A => n1135, ZN => n1120);
   U2335 : OAI221_X1 port map( B1 => n3198, B2 => n4982, C1 => n3230, C2 => 
                           n4978, A => n1136, ZN => n1119);
   U2336 : OAI22_X1 port map( A1 => n3071, A2 => n5042, B1 => n1099, B2 => 
                           n5038, ZN => n4127);
   U2337 : NOR4_X1 port map( A1 => n1100, A2 => n1101, A3 => n1102, A4 => n1103
                           , ZN => n1099);
   U2338 : OAI221_X1 port map( B1 => n3295, B2 => n4998, C1 => n3103, C2 => 
                           n4994, A => n1116, ZN => n1101);
   U2339 : OAI221_X1 port map( B1 => n3199, B2 => n4982, C1 => n3231, C2 => 
                           n4978, A => n1117, ZN => n1100);
   U2340 : OAI22_X1 port map( A1 => n3072, A2 => n5042, B1 => n1080, B2 => 
                           n5038, ZN => n4128);
   U2341 : NOR4_X1 port map( A1 => n1081, A2 => n1082, A3 => n1083, A4 => n1084
                           , ZN => n1080);
   U2342 : OAI221_X1 port map( B1 => n3296, B2 => n4998, C1 => n3104, C2 => 
                           n4994, A => n1097, ZN => n1082);
   U2343 : OAI221_X1 port map( B1 => n3200, B2 => n4982, C1 => n3232, C2 => 
                           n4978, A => n1098, ZN => n1081);
   U2344 : OAI22_X1 port map( A1 => n3651, A2 => n4483, B1 => n3587, B2 => 
                           n4491, ZN => n2673);
   U2345 : OAI22_X1 port map( A1 => n3652, A2 => n4483, B1 => n3588, B2 => 
                           n4491, ZN => n2651);
   U2346 : OAI22_X1 port map( A1 => n3653, A2 => n4483, B1 => n3589, B2 => 
                           n4491, ZN => n2632);
   U2347 : OAI22_X1 port map( A1 => n3654, A2 => n4483, B1 => n3590, B2 => 
                           n4491, ZN => n2613);
   U2348 : OAI22_X1 port map( A1 => n3655, A2 => n4483, B1 => n3591, B2 => 
                           n4491, ZN => n2594);
   U2349 : OAI22_X1 port map( A1 => n3656, A2 => n4483, B1 => n3592, B2 => 
                           n4491, ZN => n2575);
   U2350 : OAI22_X1 port map( A1 => n3657, A2 => n4484, B1 => n3593, B2 => 
                           n4492, ZN => n2556);
   U2351 : OAI22_X1 port map( A1 => n3658, A2 => n4484, B1 => n3594, B2 => 
                           n4492, ZN => n2537);
   U2352 : OAI22_X1 port map( A1 => n3659, A2 => n4484, B1 => n3595, B2 => 
                           n4492, ZN => n2518);
   U2353 : OAI22_X1 port map( A1 => n3660, A2 => n4484, B1 => n3596, B2 => 
                           n4492, ZN => n2499);
   U2354 : OAI22_X1 port map( A1 => n3661, A2 => n4484, B1 => n3597, B2 => 
                           n4492, ZN => n2480);
   U2355 : OAI22_X1 port map( A1 => n3662, A2 => n4484, B1 => n3598, B2 => 
                           n4492, ZN => n2461);
   U2356 : OAI22_X1 port map( A1 => n3663, A2 => n4485, B1 => n3599, B2 => 
                           n4493, ZN => n2442);
   U2357 : OAI22_X1 port map( A1 => n3664, A2 => n4485, B1 => n3600, B2 => 
                           n4493, ZN => n2423);
   U2358 : OAI22_X1 port map( A1 => n3665, A2 => n4485, B1 => n3601, B2 => 
                           n4493, ZN => n2404);
   U2359 : OAI22_X1 port map( A1 => n3666, A2 => n4485, B1 => n3602, B2 => 
                           n4493, ZN => n2385);
   U2360 : OAI22_X1 port map( A1 => n3667, A2 => n4485, B1 => n3603, B2 => 
                           n4493, ZN => n2366);
   U2361 : OAI22_X1 port map( A1 => n3668, A2 => n4485, B1 => n3604, B2 => 
                           n4493, ZN => n2347);
   U2362 : OAI22_X1 port map( A1 => n3669, A2 => n4486, B1 => n3605, B2 => 
                           n4494, ZN => n2328);
   U2363 : OAI22_X1 port map( A1 => n3670, A2 => n4486, B1 => n3606, B2 => 
                           n4494, ZN => n1285);
   U2364 : OAI22_X1 port map( A1 => n3671, A2 => n4486, B1 => n3607, B2 => 
                           n4494, ZN => n1266);
   U2365 : OAI22_X1 port map( A1 => n3672, A2 => n4486, B1 => n3608, B2 => 
                           n4494, ZN => n1247);
   U2366 : OAI22_X1 port map( A1 => n3673, A2 => n4486, B1 => n3609, B2 => 
                           n4494, ZN => n1228);
   U2367 : OAI22_X1 port map( A1 => n3674, A2 => n4486, B1 => n3610, B2 => 
                           n4494, ZN => n1209);
   U2368 : OAI22_X1 port map( A1 => n3675, A2 => n4487, B1 => n3611, B2 => 
                           n4495, ZN => n1190);
   U2369 : OAI22_X1 port map( A1 => n3676, A2 => n4487, B1 => n3612, B2 => 
                           n4495, ZN => n1171);
   U2370 : OAI22_X1 port map( A1 => n3677, A2 => n4487, B1 => n3613, B2 => 
                           n4495, ZN => n1152);
   U2371 : OAI22_X1 port map( A1 => n3678, A2 => n4487, B1 => n3614, B2 => 
                           n4495, ZN => n1133);
   U2372 : OAI22_X1 port map( A1 => n3679, A2 => n4487, B1 => n3615, B2 => 
                           n4495, ZN => n1114);
   U2373 : OAI22_X1 port map( A1 => n3680, A2 => n4487, B1 => n3616, B2 => 
                           n4495, ZN => n1095);
   U2374 : INV_X1 port map( A => ADD_RD2(0), ZN => n5131);
   U2375 : NOR3_X1 port map( A1 => n5150, A2 => ADD_RD1(1), A3 => n5144, ZN => 
                           n1002);
   U2376 : OAI22_X1 port map( A1 => n3011, A2 => n5120, B1 => n993, B2 => n5116
                           , ZN => n4131);
   U2377 : NOR4_X1 port map( A1 => n994, A2 => n995, A3 => n996, A4 => n997, ZN
                           => n993);
   U2378 : OAI221_X1 port map( B1 => n3171, B2 => n5060, C1 => n3203, C2 => 
                           n5056, A => n1021, ZN => n994);
   U2379 : OAI221_X1 port map( B1 => n3267, B2 => n5076, C1 => n3075, C2 => 
                           n5072, A => n1019, ZN => n995);
   U2380 : OAI22_X1 port map( A1 => n3012, A2 => n5120, B1 => n974, B2 => n5116
                           , ZN => n4132);
   U2381 : NOR4_X1 port map( A1 => n975, A2 => n976, A3 => n977, A4 => n978, ZN
                           => n974);
   U2382 : OAI221_X1 port map( B1 => n3172, B2 => n5060, C1 => n3204, C2 => 
                           n5056, A => n992, ZN => n975);
   U2383 : OAI221_X1 port map( B1 => n3268, B2 => n5076, C1 => n3076, C2 => 
                           n5072, A => n991, ZN => n976);
   U2384 : OAI22_X1 port map( A1 => n3013, A2 => n5120, B1 => n955, B2 => n5116
                           , ZN => n4133);
   U2385 : NOR4_X1 port map( A1 => n956, A2 => n957, A3 => n958, A4 => n959, ZN
                           => n955);
   U2386 : OAI221_X1 port map( B1 => n3173, B2 => n5060, C1 => n3205, C2 => 
                           n5056, A => n973, ZN => n956);
   U2387 : OAI221_X1 port map( B1 => n3269, B2 => n5076, C1 => n3077, C2 => 
                           n5072, A => n972, ZN => n957);
   U2388 : OAI22_X1 port map( A1 => n3014, A2 => n5120, B1 => n936, B2 => n5116
                           , ZN => n4134);
   U2389 : NOR4_X1 port map( A1 => n937, A2 => n938, A3 => n939, A4 => n940, ZN
                           => n936);
   U2390 : OAI221_X1 port map( B1 => n3174, B2 => n5060, C1 => n3206, C2 => 
                           n5056, A => n954, ZN => n937);
   U2391 : OAI221_X1 port map( B1 => n3270, B2 => n5076, C1 => n3078, C2 => 
                           n5072, A => n953, ZN => n938);
   U2392 : OAI22_X1 port map( A1 => n3015, A2 => n5120, B1 => n917, B2 => n5116
                           , ZN => n4135);
   U2393 : NOR4_X1 port map( A1 => n918, A2 => n919, A3 => n920, A4 => n921, ZN
                           => n917);
   U2394 : OAI221_X1 port map( B1 => n3175, B2 => n5060, C1 => n3207, C2 => 
                           n5056, A => n935, ZN => n918);
   U2395 : OAI221_X1 port map( B1 => n3271, B2 => n5076, C1 => n3079, C2 => 
                           n5072, A => n934, ZN => n919);
   U2396 : OAI22_X1 port map( A1 => n3016, A2 => n5120, B1 => n898, B2 => n5116
                           , ZN => n4136);
   U2397 : NOR4_X1 port map( A1 => n899, A2 => n900, A3 => n901, A4 => n902, ZN
                           => n898);
   U2398 : OAI221_X1 port map( B1 => n3176, B2 => n5060, C1 => n3208, C2 => 
                           n5056, A => n916, ZN => n899);
   U2399 : OAI221_X1 port map( B1 => n3272, B2 => n5076, C1 => n3080, C2 => 
                           n5072, A => n915, ZN => n900);
   U2400 : OAI22_X1 port map( A1 => n3017, A2 => n5120, B1 => n879, B2 => n5116
                           , ZN => n4137);
   U2401 : NOR4_X1 port map( A1 => n880, A2 => n881, A3 => n882, A4 => n883, ZN
                           => n879);
   U2402 : OAI221_X1 port map( B1 => n3177, B2 => n5060, C1 => n3209, C2 => 
                           n5056, A => n897, ZN => n880);
   U2403 : OAI221_X1 port map( B1 => n3273, B2 => n5076, C1 => n3081, C2 => 
                           n5072, A => n896, ZN => n881);
   U2404 : OAI22_X1 port map( A1 => n3018, A2 => n5120, B1 => n860, B2 => n5116
                           , ZN => n4138);
   U2405 : NOR4_X1 port map( A1 => n861, A2 => n862, A3 => n863, A4 => n864, ZN
                           => n860);
   U2406 : OAI221_X1 port map( B1 => n3178, B2 => n5060, C1 => n3210, C2 => 
                           n5056, A => n878, ZN => n861);
   U2407 : OAI221_X1 port map( B1 => n3274, B2 => n5076, C1 => n3082, C2 => 
                           n5072, A => n877, ZN => n862);
   U2408 : OAI22_X1 port map( A1 => n3019, A2 => n5120, B1 => n841, B2 => n5116
                           , ZN => n4139);
   U2409 : NOR4_X1 port map( A1 => n842, A2 => n843, A3 => n844, A4 => n845, ZN
                           => n841);
   U2410 : OAI221_X1 port map( B1 => n3179, B2 => n5060, C1 => n3211, C2 => 
                           n5056, A => n859, ZN => n842);
   U2411 : OAI221_X1 port map( B1 => n3275, B2 => n5076, C1 => n3083, C2 => 
                           n5072, A => n858, ZN => n843);
   U2412 : OAI22_X1 port map( A1 => n3020, A2 => n5120, B1 => n822, B2 => n5116
                           , ZN => n4140);
   U2413 : NOR4_X1 port map( A1 => n823, A2 => n824, A3 => n825, A4 => n826, ZN
                           => n822);
   U2414 : OAI221_X1 port map( B1 => n3180, B2 => n5060, C1 => n3212, C2 => 
                           n5056, A => n840, ZN => n823);
   U2415 : OAI221_X1 port map( B1 => n3276, B2 => n5076, C1 => n3084, C2 => 
                           n5072, A => n839, ZN => n824);
   U2416 : OAI22_X1 port map( A1 => n3021, A2 => n5120, B1 => n803, B2 => n5116
                           , ZN => n4141);
   U2417 : NOR4_X1 port map( A1 => n804, A2 => n805, A3 => n806, A4 => n807, ZN
                           => n803);
   U2418 : OAI221_X1 port map( B1 => n3181, B2 => n5060, C1 => n3213, C2 => 
                           n5056, A => n821, ZN => n804);
   U2419 : OAI221_X1 port map( B1 => n3277, B2 => n5076, C1 => n3085, C2 => 
                           n5072, A => n820, ZN => n805);
   U2420 : OAI22_X1 port map( A1 => n3022, A2 => n5120, B1 => n784, B2 => n5117
                           , ZN => n4142);
   U2421 : NOR4_X1 port map( A1 => n785, A2 => n786, A3 => n787, A4 => n788, ZN
                           => n784);
   U2422 : OAI221_X1 port map( B1 => n3182, B2 => n5060, C1 => n3214, C2 => 
                           n5056, A => n802, ZN => n785);
   U2423 : OAI221_X1 port map( B1 => n3278, B2 => n5076, C1 => n3086, C2 => 
                           n5072, A => n801, ZN => n786);
   U2424 : OAI22_X1 port map( A1 => n3023, A2 => n5121, B1 => n765, B2 => n5117
                           , ZN => n4143);
   U2425 : NOR4_X1 port map( A1 => n766, A2 => n767, A3 => n768, A4 => n769, ZN
                           => n765);
   U2426 : OAI221_X1 port map( B1 => n3183, B2 => n5061, C1 => n3215, C2 => 
                           n5057, A => n783, ZN => n766);
   U2427 : OAI221_X1 port map( B1 => n3279, B2 => n5077, C1 => n3087, C2 => 
                           n5073, A => n782, ZN => n767);
   U2428 : OAI22_X1 port map( A1 => n3024, A2 => n5121, B1 => n746, B2 => n5117
                           , ZN => n4144);
   U2429 : NOR4_X1 port map( A1 => n747, A2 => n748, A3 => n749, A4 => n750, ZN
                           => n746);
   U2430 : OAI221_X1 port map( B1 => n3184, B2 => n5061, C1 => n3216, C2 => 
                           n5057, A => n764, ZN => n747);
   U2431 : OAI221_X1 port map( B1 => n3280, B2 => n5077, C1 => n3088, C2 => 
                           n5073, A => n763, ZN => n748);
   U2432 : OAI22_X1 port map( A1 => n3025, A2 => n5121, B1 => n727, B2 => n5117
                           , ZN => n4145);
   U2433 : NOR4_X1 port map( A1 => n728, A2 => n729, A3 => n730, A4 => n731, ZN
                           => n727);
   U2434 : OAI221_X1 port map( B1 => n3185, B2 => n5061, C1 => n3217, C2 => 
                           n5057, A => n745, ZN => n728);
   U2435 : OAI221_X1 port map( B1 => n3281, B2 => n5077, C1 => n3089, C2 => 
                           n5073, A => n744, ZN => n729);
   U2436 : OAI22_X1 port map( A1 => n3026, A2 => n5121, B1 => n708, B2 => n5117
                           , ZN => n4146);
   U2437 : NOR4_X1 port map( A1 => n709, A2 => n710, A3 => n711, A4 => n712, ZN
                           => n708);
   U2438 : OAI221_X1 port map( B1 => n3186, B2 => n5061, C1 => n3218, C2 => 
                           n5057, A => n726, ZN => n709);
   U2439 : OAI221_X1 port map( B1 => n3282, B2 => n5077, C1 => n3090, C2 => 
                           n5073, A => n725, ZN => n710);
   U2440 : OAI22_X1 port map( A1 => n3027, A2 => n5121, B1 => n689, B2 => n5117
                           , ZN => n4147);
   U2441 : NOR4_X1 port map( A1 => n690, A2 => n691, A3 => n692, A4 => n693, ZN
                           => n689);
   U2442 : OAI221_X1 port map( B1 => n3187, B2 => n5061, C1 => n3219, C2 => 
                           n5057, A => n707, ZN => n690);
   U2443 : OAI221_X1 port map( B1 => n3283, B2 => n5077, C1 => n3091, C2 => 
                           n5073, A => n706, ZN => n691);
   U2444 : OAI22_X1 port map( A1 => n3028, A2 => n5121, B1 => n670, B2 => n5117
                           , ZN => n4148);
   U2445 : NOR4_X1 port map( A1 => n671, A2 => n672, A3 => n673, A4 => n674, ZN
                           => n670);
   U2446 : OAI221_X1 port map( B1 => n3188, B2 => n5061, C1 => n3220, C2 => 
                           n5057, A => n688, ZN => n671);
   U2447 : OAI221_X1 port map( B1 => n3284, B2 => n5077, C1 => n3092, C2 => 
                           n5073, A => n687, ZN => n672);
   U2448 : OAI22_X1 port map( A1 => n3029, A2 => n5121, B1 => n651, B2 => n5117
                           , ZN => n4149);
   U2449 : NOR4_X1 port map( A1 => n652, A2 => n653, A3 => n654, A4 => n655, ZN
                           => n651);
   U2450 : OAI221_X1 port map( B1 => n3189, B2 => n5061, C1 => n3221, C2 => 
                           n5057, A => n669, ZN => n652);
   U2451 : OAI221_X1 port map( B1 => n3285, B2 => n5077, C1 => n3093, C2 => 
                           n5073, A => n668, ZN => n653);
   U2452 : OAI22_X1 port map( A1 => n3030, A2 => n5121, B1 => n632, B2 => n5117
                           , ZN => n4150);
   U2453 : NOR4_X1 port map( A1 => n633, A2 => n634, A3 => n635, A4 => n636, ZN
                           => n632);
   U2454 : OAI221_X1 port map( B1 => n3190, B2 => n5061, C1 => n3222, C2 => 
                           n5057, A => n650, ZN => n633);
   U2455 : OAI221_X1 port map( B1 => n3286, B2 => n5077, C1 => n3094, C2 => 
                           n5073, A => n649, ZN => n634);
   U2456 : OAI22_X1 port map( A1 => n3031, A2 => n5121, B1 => n613, B2 => n5117
                           , ZN => n4151);
   U2457 : NOR4_X1 port map( A1 => n614, A2 => n615, A3 => n616, A4 => n617, ZN
                           => n613);
   U2458 : OAI221_X1 port map( B1 => n3191, B2 => n5061, C1 => n3223, C2 => 
                           n5057, A => n631, ZN => n614);
   U2459 : OAI221_X1 port map( B1 => n3287, B2 => n5077, C1 => n3095, C2 => 
                           n5073, A => n630, ZN => n615);
   U2460 : OAI22_X1 port map( A1 => n3032, A2 => n5121, B1 => n594, B2 => n5117
                           , ZN => n4152);
   U2461 : NOR4_X1 port map( A1 => n595, A2 => n596, A3 => n597, A4 => n598, ZN
                           => n594);
   U2462 : OAI221_X1 port map( B1 => n3192, B2 => n5061, C1 => n3224, C2 => 
                           n5057, A => n612, ZN => n595);
   U2463 : OAI221_X1 port map( B1 => n3288, B2 => n5077, C1 => n3096, C2 => 
                           n5073, A => n611, ZN => n596);
   U2464 : OAI22_X1 port map( A1 => n3033, A2 => n5121, B1 => n575, B2 => n5117
                           , ZN => n4153);
   U2465 : NOR4_X1 port map( A1 => n576, A2 => n577, A3 => n578, A4 => n579, ZN
                           => n575);
   U2466 : OAI221_X1 port map( B1 => n3193, B2 => n5061, C1 => n3225, C2 => 
                           n5057, A => n593, ZN => n576);
   U2467 : OAI221_X1 port map( B1 => n3289, B2 => n5077, C1 => n3097, C2 => 
                           n5073, A => n592, ZN => n577);
   U2468 : OAI22_X1 port map( A1 => n3034, A2 => n5121, B1 => n556, B2 => n5118
                           , ZN => n4154);
   U2469 : NOR4_X1 port map( A1 => n557, A2 => n558, A3 => n559, A4 => n560, ZN
                           => n556);
   U2470 : OAI221_X1 port map( B1 => n3194, B2 => n5061, C1 => n3226, C2 => 
                           n5057, A => n574, ZN => n557);
   U2471 : OAI221_X1 port map( B1 => n3290, B2 => n5077, C1 => n3098, C2 => 
                           n5073, A => n573, ZN => n558);
   U2472 : OAI22_X1 port map( A1 => n3035, A2 => n5122, B1 => n537, B2 => n5118
                           , ZN => n4155);
   U2473 : NOR4_X1 port map( A1 => n538, A2 => n539, A3 => n540, A4 => n541, ZN
                           => n537);
   U2474 : OAI221_X1 port map( B1 => n3195, B2 => n5062, C1 => n3227, C2 => 
                           n5058, A => n555, ZN => n538);
   U2475 : OAI221_X1 port map( B1 => n3291, B2 => n5078, C1 => n3099, C2 => 
                           n5074, A => n554, ZN => n539);
   U2476 : OAI22_X1 port map( A1 => n3036, A2 => n5122, B1 => n518, B2 => n5118
                           , ZN => n4156);
   U2477 : NOR4_X1 port map( A1 => n519, A2 => n520, A3 => n521, A4 => n522, ZN
                           => n518);
   U2478 : OAI221_X1 port map( B1 => n3196, B2 => n5062, C1 => n3228, C2 => 
                           n5058, A => n536, ZN => n519);
   U2479 : OAI221_X1 port map( B1 => n3292, B2 => n5078, C1 => n3100, C2 => 
                           n5074, A => n535, ZN => n520);
   U2480 : OAI22_X1 port map( A1 => n3037, A2 => n5122, B1 => n499, B2 => n5118
                           , ZN => n4157);
   U2481 : NOR4_X1 port map( A1 => n500, A2 => n501, A3 => n502, A4 => n503, ZN
                           => n499);
   U2482 : OAI221_X1 port map( B1 => n3197, B2 => n5062, C1 => n3229, C2 => 
                           n5058, A => n517, ZN => n500);
   U2483 : OAI221_X1 port map( B1 => n3293, B2 => n5078, C1 => n3101, C2 => 
                           n5074, A => n516, ZN => n501);
   U2484 : OAI22_X1 port map( A1 => n3038, A2 => n5122, B1 => n480, B2 => n5118
                           , ZN => n4158);
   U2485 : NOR4_X1 port map( A1 => n481, A2 => n482, A3 => n483, A4 => n484, ZN
                           => n480);
   U2486 : OAI221_X1 port map( B1 => n3198, B2 => n5062, C1 => n3230, C2 => 
                           n5058, A => n498, ZN => n481);
   U2487 : OAI221_X1 port map( B1 => n3294, B2 => n5078, C1 => n3102, C2 => 
                           n5074, A => n497, ZN => n482);
   U2488 : OAI22_X1 port map( A1 => n3039, A2 => n5122, B1 => n461, B2 => n5118
                           , ZN => n4159);
   U2489 : NOR4_X1 port map( A1 => n462, A2 => n463, A3 => n464, A4 => n465, ZN
                           => n461);
   U2490 : OAI221_X1 port map( B1 => n3199, B2 => n5062, C1 => n3231, C2 => 
                           n5058, A => n479, ZN => n462);
   U2491 : OAI221_X1 port map( B1 => n3295, B2 => n5078, C1 => n3103, C2 => 
                           n5074, A => n478, ZN => n463);
   U2492 : OAI22_X1 port map( A1 => n3040, A2 => n5122, B1 => n442, B2 => n5118
                           , ZN => n4160);
   U2493 : NOR4_X1 port map( A1 => n443, A2 => n444, A3 => n445, A4 => n446, ZN
                           => n442);
   U2494 : OAI221_X1 port map( B1 => n3200, B2 => n5062, C1 => n3232, C2 => 
                           n5058, A => n460, ZN => n443);
   U2495 : OAI221_X1 port map( B1 => n3296, B2 => n5078, C1 => n3104, C2 => 
                           n5074, A => n459, ZN => n444);
   U2496 : OAI22_X1 port map( A1 => n3651, A2 => n4547, B1 => n3587, B2 => 
                           n4555, ZN => n1011);
   U2497 : OAI22_X1 port map( A1 => n3652, A2 => n4547, B1 => n3588, B2 => 
                           n4555, ZN => n989);
   U2498 : OAI22_X1 port map( A1 => n3653, A2 => n4547, B1 => n3589, B2 => 
                           n4555, ZN => n970);
   U2499 : OAI22_X1 port map( A1 => n3654, A2 => n4547, B1 => n3590, B2 => 
                           n4555, ZN => n951);
   U2500 : OAI22_X1 port map( A1 => n3655, A2 => n4547, B1 => n3591, B2 => 
                           n4555, ZN => n932);
   U2501 : OAI22_X1 port map( A1 => n3656, A2 => n4547, B1 => n3592, B2 => 
                           n4555, ZN => n913);
   U2502 : OAI22_X1 port map( A1 => n3657, A2 => n4548, B1 => n3593, B2 => 
                           n4556, ZN => n894);
   U2503 : OAI22_X1 port map( A1 => n3658, A2 => n4548, B1 => n3594, B2 => 
                           n4556, ZN => n875);
   U2504 : OAI22_X1 port map( A1 => n3659, A2 => n4548, B1 => n3595, B2 => 
                           n4556, ZN => n856);
   U2505 : OAI22_X1 port map( A1 => n3660, A2 => n4548, B1 => n3596, B2 => 
                           n4556, ZN => n837);
   U2506 : OAI22_X1 port map( A1 => n3661, A2 => n4548, B1 => n3597, B2 => 
                           n4556, ZN => n818);
   U2507 : OAI22_X1 port map( A1 => n3662, A2 => n4548, B1 => n3598, B2 => 
                           n4556, ZN => n799);
   U2508 : OAI22_X1 port map( A1 => n3663, A2 => n4549, B1 => n3599, B2 => 
                           n4557, ZN => n780);
   U2509 : OAI22_X1 port map( A1 => n3664, A2 => n4549, B1 => n3600, B2 => 
                           n4557, ZN => n761);
   U2510 : OAI22_X1 port map( A1 => n3665, A2 => n4549, B1 => n3601, B2 => 
                           n4557, ZN => n742);
   U2511 : OAI22_X1 port map( A1 => n3666, A2 => n4549, B1 => n3602, B2 => 
                           n4557, ZN => n723);
   U2512 : OAI22_X1 port map( A1 => n3667, A2 => n4549, B1 => n3603, B2 => 
                           n4557, ZN => n704);
   U2513 : OAI22_X1 port map( A1 => n3668, A2 => n4549, B1 => n3604, B2 => 
                           n4557, ZN => n685);
   U2514 : OAI22_X1 port map( A1 => n3669, A2 => n4550, B1 => n3605, B2 => 
                           n4558, ZN => n666);
   U2515 : OAI22_X1 port map( A1 => n3670, A2 => n4550, B1 => n3606, B2 => 
                           n4558, ZN => n647);
   U2516 : OAI22_X1 port map( A1 => n3671, A2 => n4550, B1 => n3607, B2 => 
                           n4558, ZN => n628);
   U2517 : OAI22_X1 port map( A1 => n3672, A2 => n4550, B1 => n3608, B2 => 
                           n4558, ZN => n609);
   U2518 : OAI22_X1 port map( A1 => n3673, A2 => n4550, B1 => n3609, B2 => 
                           n4558, ZN => n590);
   U2519 : OAI22_X1 port map( A1 => n3674, A2 => n4550, B1 => n3610, B2 => 
                           n4558, ZN => n571);
   U2520 : OAI22_X1 port map( A1 => n3675, A2 => n4551, B1 => n3611, B2 => 
                           n4559, ZN => n552);
   U2521 : OAI22_X1 port map( A1 => n3676, A2 => n4551, B1 => n3612, B2 => 
                           n4559, ZN => n533);
   U2522 : OAI22_X1 port map( A1 => n3677, A2 => n4551, B1 => n3613, B2 => 
                           n4559, ZN => n514);
   U2523 : OAI22_X1 port map( A1 => n3678, A2 => n4551, B1 => n3614, B2 => 
                           n4559, ZN => n495);
   U2524 : OAI22_X1 port map( A1 => n3679, A2 => n4551, B1 => n3615, B2 => 
                           n4559, ZN => n476);
   U2525 : OAI22_X1 port map( A1 => n3680, A2 => n4551, B1 => n3616, B2 => 
                           n4559, ZN => n457);
   U2526 : INV_X1 port map( A => ADD_RD1(0), ZN => n5144);
   U2527 : NOR3_X1 port map( A1 => n5136, A2 => ADD_RD2(2), A3 => n5131, ZN => 
                           n2674);
   U2528 : OAI22_X1 port map( A1 => n3779, A2 => n4499, B1 => n3715, B2 => 
                           n4507, ZN => n2672);
   U2529 : OAI22_X1 port map( A1 => n3780, A2 => n4499, B1 => n3716, B2 => 
                           n4507, ZN => n2650);
   U2530 : OAI22_X1 port map( A1 => n3781, A2 => n4499, B1 => n3717, B2 => 
                           n4507, ZN => n2631);
   U2531 : OAI22_X1 port map( A1 => n3782, A2 => n4499, B1 => n3718, B2 => 
                           n4507, ZN => n2612);
   U2532 : OAI22_X1 port map( A1 => n3783, A2 => n4499, B1 => n3719, B2 => 
                           n4507, ZN => n2593);
   U2533 : OAI22_X1 port map( A1 => n3784, A2 => n4499, B1 => n3720, B2 => 
                           n4507, ZN => n2574);
   U2534 : OAI22_X1 port map( A1 => n3785, A2 => n4500, B1 => n3721, B2 => 
                           n4508, ZN => n2555);
   U2535 : OAI22_X1 port map( A1 => n3786, A2 => n4500, B1 => n3722, B2 => 
                           n4508, ZN => n2536);
   U2536 : OAI22_X1 port map( A1 => n3787, A2 => n4500, B1 => n3723, B2 => 
                           n4508, ZN => n2517);
   U2537 : OAI22_X1 port map( A1 => n3788, A2 => n4500, B1 => n3724, B2 => 
                           n4508, ZN => n2498);
   U2538 : OAI22_X1 port map( A1 => n3789, A2 => n4500, B1 => n3725, B2 => 
                           n4508, ZN => n2479);
   U2539 : OAI22_X1 port map( A1 => n3790, A2 => n4500, B1 => n3726, B2 => 
                           n4508, ZN => n2460);
   U2540 : OAI22_X1 port map( A1 => n3791, A2 => n4501, B1 => n3727, B2 => 
                           n4509, ZN => n2441);
   U2541 : OAI22_X1 port map( A1 => n3792, A2 => n4501, B1 => n3728, B2 => 
                           n4509, ZN => n2422);
   U2542 : OAI22_X1 port map( A1 => n3793, A2 => n4501, B1 => n3729, B2 => 
                           n4509, ZN => n2403);
   U2543 : OAI22_X1 port map( A1 => n3794, A2 => n4501, B1 => n3730, B2 => 
                           n4509, ZN => n2384);
   U2544 : OAI22_X1 port map( A1 => n3795, A2 => n4501, B1 => n3731, B2 => 
                           n4509, ZN => n2365);
   U2545 : OAI22_X1 port map( A1 => n3796, A2 => n4501, B1 => n3732, B2 => 
                           n4509, ZN => n2346);
   U2546 : OAI22_X1 port map( A1 => n3797, A2 => n4502, B1 => n3733, B2 => 
                           n4510, ZN => n2327);
   U2547 : OAI22_X1 port map( A1 => n3798, A2 => n4502, B1 => n3734, B2 => 
                           n4510, ZN => n1284);
   U2548 : OAI22_X1 port map( A1 => n3799, A2 => n4502, B1 => n3735, B2 => 
                           n4510, ZN => n1265);
   U2549 : OAI22_X1 port map( A1 => n3800, A2 => n4502, B1 => n3736, B2 => 
                           n4510, ZN => n1246);
   U2550 : OAI22_X1 port map( A1 => n3801, A2 => n4502, B1 => n3737, B2 => 
                           n4510, ZN => n1227);
   U2551 : OAI22_X1 port map( A1 => n3802, A2 => n4502, B1 => n3738, B2 => 
                           n4510, ZN => n1208);
   U2552 : OAI22_X1 port map( A1 => n3803, A2 => n4503, B1 => n3739, B2 => 
                           n4511, ZN => n1189);
   U2553 : OAI22_X1 port map( A1 => n3804, A2 => n4503, B1 => n3740, B2 => 
                           n4511, ZN => n1170);
   U2554 : OAI22_X1 port map( A1 => n3805, A2 => n4503, B1 => n3741, B2 => 
                           n4511, ZN => n1151);
   U2555 : OAI22_X1 port map( A1 => n3806, A2 => n4503, B1 => n3742, B2 => 
                           n4511, ZN => n1132);
   U2556 : OAI22_X1 port map( A1 => n3807, A2 => n4503, B1 => n3743, B2 => 
                           n4511, ZN => n1113);
   U2557 : OAI22_X1 port map( A1 => n3808, A2 => n4503, B1 => n3744, B2 => 
                           n4511, ZN => n1094);
   U2558 : NOR3_X1 port map( A1 => n5149, A2 => ADD_RD1(2), A3 => n5144, ZN => 
                           n1012);
   U2559 : OAI22_X1 port map( A1 => n3779, A2 => n4563, B1 => n3715, B2 => 
                           n4571, ZN => n1010);
   U2560 : OAI22_X1 port map( A1 => n3780, A2 => n4563, B1 => n3716, B2 => 
                           n4571, ZN => n988);
   U2561 : OAI22_X1 port map( A1 => n3781, A2 => n4563, B1 => n3717, B2 => 
                           n4571, ZN => n969);
   U2562 : OAI22_X1 port map( A1 => n3782, A2 => n4563, B1 => n3718, B2 => 
                           n4571, ZN => n950);
   U2563 : OAI22_X1 port map( A1 => n3783, A2 => n4563, B1 => n3719, B2 => 
                           n4571, ZN => n931);
   U2564 : OAI22_X1 port map( A1 => n3784, A2 => n4563, B1 => n3720, B2 => 
                           n4571, ZN => n912);
   U2565 : OAI22_X1 port map( A1 => n3785, A2 => n4564, B1 => n3721, B2 => 
                           n4572, ZN => n893);
   U2566 : OAI22_X1 port map( A1 => n3786, A2 => n4564, B1 => n3722, B2 => 
                           n4572, ZN => n874);
   U2567 : OAI22_X1 port map( A1 => n3787, A2 => n4564, B1 => n3723, B2 => 
                           n4572, ZN => n855);
   U2568 : OAI22_X1 port map( A1 => n3788, A2 => n4564, B1 => n3724, B2 => 
                           n4572, ZN => n836);
   U2569 : OAI22_X1 port map( A1 => n3789, A2 => n4564, B1 => n3725, B2 => 
                           n4572, ZN => n817);
   U2570 : OAI22_X1 port map( A1 => n3790, A2 => n4564, B1 => n3726, B2 => 
                           n4572, ZN => n798);
   U2571 : OAI22_X1 port map( A1 => n3791, A2 => n4565, B1 => n3727, B2 => 
                           n4573, ZN => n779);
   U2572 : OAI22_X1 port map( A1 => n3792, A2 => n4565, B1 => n3728, B2 => 
                           n4573, ZN => n760);
   U2573 : OAI22_X1 port map( A1 => n3793, A2 => n4565, B1 => n3729, B2 => 
                           n4573, ZN => n741);
   U2574 : OAI22_X1 port map( A1 => n3794, A2 => n4565, B1 => n3730, B2 => 
                           n4573, ZN => n722);
   U2575 : OAI22_X1 port map( A1 => n3795, A2 => n4565, B1 => n3731, B2 => 
                           n4573, ZN => n703);
   U2576 : OAI22_X1 port map( A1 => n3796, A2 => n4565, B1 => n3732, B2 => 
                           n4573, ZN => n684);
   U2577 : OAI22_X1 port map( A1 => n3797, A2 => n4566, B1 => n3733, B2 => 
                           n4574, ZN => n665);
   U2578 : OAI22_X1 port map( A1 => n3798, A2 => n4566, B1 => n3734, B2 => 
                           n4574, ZN => n646);
   U2579 : OAI22_X1 port map( A1 => n3799, A2 => n4566, B1 => n3735, B2 => 
                           n4574, ZN => n627);
   U2580 : OAI22_X1 port map( A1 => n3800, A2 => n4566, B1 => n3736, B2 => 
                           n4574, ZN => n608);
   U2581 : OAI22_X1 port map( A1 => n3801, A2 => n4566, B1 => n3737, B2 => 
                           n4574, ZN => n589);
   U2582 : OAI22_X1 port map( A1 => n3802, A2 => n4566, B1 => n3738, B2 => 
                           n4574, ZN => n570);
   U2583 : OAI22_X1 port map( A1 => n3803, A2 => n4567, B1 => n3739, B2 => 
                           n4575, ZN => n551);
   U2584 : OAI22_X1 port map( A1 => n3804, A2 => n4567, B1 => n3740, B2 => 
                           n4575, ZN => n532);
   U2585 : OAI22_X1 port map( A1 => n3805, A2 => n4567, B1 => n3741, B2 => 
                           n4575, ZN => n513);
   U2586 : OAI22_X1 port map( A1 => n3806, A2 => n4567, B1 => n3742, B2 => 
                           n4575, ZN => n494);
   U2587 : OAI22_X1 port map( A1 => n3807, A2 => n4567, B1 => n3743, B2 => 
                           n4575, ZN => n475);
   U2588 : OAI22_X1 port map( A1 => n3808, A2 => n4567, B1 => n3744, B2 => 
                           n4575, ZN => n456);
   U2589 : INV_X1 port map( A => ADD_RD2(2), ZN => n5137);
   U2590 : INV_X1 port map( A => ADD_RD2(1), ZN => n5136);
   U2591 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n5131, 
                           ZN => n2675);
   U2592 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n5144, 
                           ZN => n1013);
   U2593 : INV_X1 port map( A => ADD_RD1(1), ZN => n5149);
   U2594 : INV_X1 port map( A => ADD_RD1(2), ZN => n5150);
   U2595 : OAI22_X1 port map( A1 => n3907, A2 => n4483, B1 => n3843, B2 => 
                           n4491, ZN => n2669);
   U2596 : OAI22_X1 port map( A1 => n3908, A2 => n4483, B1 => n3844, B2 => 
                           n4491, ZN => n2647);
   U2597 : OAI22_X1 port map( A1 => n3909, A2 => n4483, B1 => n3845, B2 => 
                           n4491, ZN => n2628);
   U2598 : OAI22_X1 port map( A1 => n3910, A2 => n4483, B1 => n3846, B2 => 
                           n4491, ZN => n2609);
   U2599 : OAI22_X1 port map( A1 => n3911, A2 => n4483, B1 => n3847, B2 => 
                           n4491, ZN => n2590);
   U2600 : OAI22_X1 port map( A1 => n3912, A2 => n4483, B1 => n3848, B2 => 
                           n4491, ZN => n2571);
   U2601 : OAI22_X1 port map( A1 => n3913, A2 => n4484, B1 => n3849, B2 => 
                           n4492, ZN => n2552);
   U2602 : OAI22_X1 port map( A1 => n3914, A2 => n4484, B1 => n3850, B2 => 
                           n4492, ZN => n2533);
   U2603 : OAI22_X1 port map( A1 => n3915, A2 => n4484, B1 => n3851, B2 => 
                           n4492, ZN => n2514);
   U2604 : OAI22_X1 port map( A1 => n3916, A2 => n4484, B1 => n3852, B2 => 
                           n4492, ZN => n2495);
   U2605 : OAI22_X1 port map( A1 => n3917, A2 => n4484, B1 => n3853, B2 => 
                           n4492, ZN => n2476);
   U2606 : OAI22_X1 port map( A1 => n3918, A2 => n4484, B1 => n3854, B2 => 
                           n4492, ZN => n2457);
   U2607 : OAI22_X1 port map( A1 => n3919, A2 => n4485, B1 => n3855, B2 => 
                           n4493, ZN => n2438);
   U2608 : OAI22_X1 port map( A1 => n3920, A2 => n4485, B1 => n3856, B2 => 
                           n4493, ZN => n2419);
   U2609 : OAI22_X1 port map( A1 => n3921, A2 => n4485, B1 => n3857, B2 => 
                           n4493, ZN => n2400);
   U2610 : OAI22_X1 port map( A1 => n3922, A2 => n4485, B1 => n3858, B2 => 
                           n4493, ZN => n2381);
   U2611 : OAI22_X1 port map( A1 => n3923, A2 => n4485, B1 => n3859, B2 => 
                           n4493, ZN => n2362);
   U2612 : OAI22_X1 port map( A1 => n3924, A2 => n4485, B1 => n3860, B2 => 
                           n4493, ZN => n2343);
   U2613 : OAI22_X1 port map( A1 => n3925, A2 => n4486, B1 => n3861, B2 => 
                           n4494, ZN => n1300);
   U2614 : OAI22_X1 port map( A1 => n3926, A2 => n4486, B1 => n3862, B2 => 
                           n4494, ZN => n1281);
   U2615 : OAI22_X1 port map( A1 => n3927, A2 => n4486, B1 => n3863, B2 => 
                           n4494, ZN => n1262);
   U2616 : OAI22_X1 port map( A1 => n3928, A2 => n4486, B1 => n3864, B2 => 
                           n4494, ZN => n1243);
   U2617 : OAI22_X1 port map( A1 => n3929, A2 => n4486, B1 => n3865, B2 => 
                           n4494, ZN => n1224);
   U2618 : OAI22_X1 port map( A1 => n3930, A2 => n4486, B1 => n3866, B2 => 
                           n4494, ZN => n1205);
   U2619 : OAI22_X1 port map( A1 => n3931, A2 => n4487, B1 => n3867, B2 => 
                           n4495, ZN => n1186);
   U2620 : OAI22_X1 port map( A1 => n3932, A2 => n4487, B1 => n3868, B2 => 
                           n4495, ZN => n1167);
   U2621 : OAI22_X1 port map( A1 => n3933, A2 => n4487, B1 => n3869, B2 => 
                           n4495, ZN => n1148);
   U2622 : OAI22_X1 port map( A1 => n3934, A2 => n4487, B1 => n3870, B2 => 
                           n4495, ZN => n1129);
   U2623 : OAI22_X1 port map( A1 => n3935, A2 => n4487, B1 => n3871, B2 => 
                           n4495, ZN => n1110);
   U2624 : OAI22_X1 port map( A1 => n3936, A2 => n4487, B1 => n3872, B2 => 
                           n4495, ZN => n1091);
   U2625 : OAI22_X1 port map( A1 => n3907, A2 => n4547, B1 => n3843, B2 => 
                           n4555, ZN => n1007);
   U2626 : OAI22_X1 port map( A1 => n3908, A2 => n4547, B1 => n3844, B2 => 
                           n4555, ZN => n985);
   U2627 : OAI22_X1 port map( A1 => n3909, A2 => n4547, B1 => n3845, B2 => 
                           n4555, ZN => n966);
   U2628 : OAI22_X1 port map( A1 => n3910, A2 => n4547, B1 => n3846, B2 => 
                           n4555, ZN => n947);
   U2629 : OAI22_X1 port map( A1 => n3911, A2 => n4547, B1 => n3847, B2 => 
                           n4555, ZN => n928);
   U2630 : OAI22_X1 port map( A1 => n3912, A2 => n4547, B1 => n3848, B2 => 
                           n4555, ZN => n909);
   U2631 : OAI22_X1 port map( A1 => n3913, A2 => n4548, B1 => n3849, B2 => 
                           n4556, ZN => n890);
   U2632 : OAI22_X1 port map( A1 => n3914, A2 => n4548, B1 => n3850, B2 => 
                           n4556, ZN => n871);
   U2633 : OAI22_X1 port map( A1 => n3915, A2 => n4548, B1 => n3851, B2 => 
                           n4556, ZN => n852);
   U2634 : OAI22_X1 port map( A1 => n3916, A2 => n4548, B1 => n3852, B2 => 
                           n4556, ZN => n833);
   U2635 : OAI22_X1 port map( A1 => n3917, A2 => n4548, B1 => n3853, B2 => 
                           n4556, ZN => n814);
   U2636 : OAI22_X1 port map( A1 => n3918, A2 => n4548, B1 => n3854, B2 => 
                           n4556, ZN => n795);
   U2637 : OAI22_X1 port map( A1 => n3919, A2 => n4549, B1 => n3855, B2 => 
                           n4557, ZN => n776);
   U2638 : OAI22_X1 port map( A1 => n3920, A2 => n4549, B1 => n3856, B2 => 
                           n4557, ZN => n757);
   U2639 : OAI22_X1 port map( A1 => n3921, A2 => n4549, B1 => n3857, B2 => 
                           n4557, ZN => n738);
   U2640 : OAI22_X1 port map( A1 => n3922, A2 => n4549, B1 => n3858, B2 => 
                           n4557, ZN => n719);
   U2641 : OAI22_X1 port map( A1 => n3923, A2 => n4549, B1 => n3859, B2 => 
                           n4557, ZN => n700);
   U2642 : OAI22_X1 port map( A1 => n3924, A2 => n4549, B1 => n3860, B2 => 
                           n4557, ZN => n681);
   U2643 : OAI22_X1 port map( A1 => n3925, A2 => n4550, B1 => n3861, B2 => 
                           n4558, ZN => n662);
   U2644 : OAI22_X1 port map( A1 => n3926, A2 => n4550, B1 => n3862, B2 => 
                           n4558, ZN => n643);
   U2645 : OAI22_X1 port map( A1 => n3927, A2 => n4550, B1 => n3863, B2 => 
                           n4558, ZN => n624);
   U2646 : OAI22_X1 port map( A1 => n3928, A2 => n4550, B1 => n3864, B2 => 
                           n4558, ZN => n605);
   U2647 : OAI22_X1 port map( A1 => n3929, A2 => n4550, B1 => n3865, B2 => 
                           n4558, ZN => n586);
   U2648 : OAI22_X1 port map( A1 => n3930, A2 => n4550, B1 => n3866, B2 => 
                           n4558, ZN => n567);
   U2649 : OAI22_X1 port map( A1 => n3931, A2 => n4551, B1 => n3867, B2 => 
                           n4559, ZN => n548);
   U2650 : OAI22_X1 port map( A1 => n3932, A2 => n4551, B1 => n3868, B2 => 
                           n4559, ZN => n529);
   U2651 : OAI22_X1 port map( A1 => n3933, A2 => n4551, B1 => n3869, B2 => 
                           n4559, ZN => n510);
   U2652 : OAI22_X1 port map( A1 => n3934, A2 => n4551, B1 => n3870, B2 => 
                           n4559, ZN => n491);
   U2653 : OAI22_X1 port map( A1 => n3935, A2 => n4551, B1 => n3871, B2 => 
                           n4559, ZN => n472);
   U2654 : OAI22_X1 port map( A1 => n3936, A2 => n4551, B1 => n3872, B2 => 
                           n4559, ZN => n453);
   U2655 : OAI22_X1 port map( A1 => n4035, A2 => n4499, B1 => n3971, B2 => 
                           n4507, ZN => n2668);
   U2656 : OAI22_X1 port map( A1 => n4036, A2 => n4499, B1 => n3972, B2 => 
                           n4507, ZN => n2646);
   U2657 : OAI22_X1 port map( A1 => n4037, A2 => n4499, B1 => n3973, B2 => 
                           n4507, ZN => n2627);
   U2658 : OAI22_X1 port map( A1 => n4038, A2 => n4499, B1 => n3974, B2 => 
                           n4507, ZN => n2608);
   U2659 : OAI22_X1 port map( A1 => n4039, A2 => n4499, B1 => n3975, B2 => 
                           n4507, ZN => n2589);
   U2660 : OAI22_X1 port map( A1 => n4040, A2 => n4499, B1 => n3976, B2 => 
                           n4507, ZN => n2570);
   U2661 : OAI22_X1 port map( A1 => n4041, A2 => n4500, B1 => n3977, B2 => 
                           n4508, ZN => n2551);
   U2662 : OAI22_X1 port map( A1 => n4042, A2 => n4500, B1 => n3978, B2 => 
                           n4508, ZN => n2532);
   U2663 : OAI22_X1 port map( A1 => n4043, A2 => n4500, B1 => n3979, B2 => 
                           n4508, ZN => n2513);
   U2664 : OAI22_X1 port map( A1 => n4044, A2 => n4500, B1 => n3980, B2 => 
                           n4508, ZN => n2494);
   U2665 : OAI22_X1 port map( A1 => n4045, A2 => n4500, B1 => n3981, B2 => 
                           n4508, ZN => n2475);
   U2666 : OAI22_X1 port map( A1 => n4046, A2 => n4500, B1 => n3982, B2 => 
                           n4508, ZN => n2456);
   U2667 : OAI22_X1 port map( A1 => n4047, A2 => n4501, B1 => n3983, B2 => 
                           n4509, ZN => n2437);
   U2668 : OAI22_X1 port map( A1 => n4048, A2 => n4501, B1 => n3984, B2 => 
                           n4509, ZN => n2418);
   U2669 : OAI22_X1 port map( A1 => n4049, A2 => n4501, B1 => n3985, B2 => 
                           n4509, ZN => n2399);
   U2670 : OAI22_X1 port map( A1 => n4050, A2 => n4501, B1 => n3986, B2 => 
                           n4509, ZN => n2380);
   U2671 : OAI22_X1 port map( A1 => n4051, A2 => n4501, B1 => n3987, B2 => 
                           n4509, ZN => n2361);
   U2672 : OAI22_X1 port map( A1 => n4052, A2 => n4501, B1 => n3988, B2 => 
                           n4509, ZN => n2342);
   U2673 : OAI22_X1 port map( A1 => n4053, A2 => n4502, B1 => n3989, B2 => 
                           n4510, ZN => n1299);
   U2674 : OAI22_X1 port map( A1 => n4054, A2 => n4502, B1 => n3990, B2 => 
                           n4510, ZN => n1280);
   U2675 : OAI22_X1 port map( A1 => n4055, A2 => n4502, B1 => n3991, B2 => 
                           n4510, ZN => n1261);
   U2676 : OAI22_X1 port map( A1 => n4056, A2 => n4502, B1 => n3992, B2 => 
                           n4510, ZN => n1242);
   U2677 : OAI22_X1 port map( A1 => n4057, A2 => n4502, B1 => n3993, B2 => 
                           n4510, ZN => n1223);
   U2678 : OAI22_X1 port map( A1 => n4058, A2 => n4502, B1 => n3994, B2 => 
                           n4510, ZN => n1204);
   U2679 : OAI22_X1 port map( A1 => n4059, A2 => n4503, B1 => n3995, B2 => 
                           n4511, ZN => n1185);
   U2680 : OAI22_X1 port map( A1 => n4060, A2 => n4503, B1 => n3996, B2 => 
                           n4511, ZN => n1166);
   U2681 : OAI22_X1 port map( A1 => n4061, A2 => n4503, B1 => n3997, B2 => 
                           n4511, ZN => n1147);
   U2682 : OAI22_X1 port map( A1 => n4062, A2 => n4503, B1 => n3998, B2 => 
                           n4511, ZN => n1128);
   U2683 : OAI22_X1 port map( A1 => n4063, A2 => n4503, B1 => n3999, B2 => 
                           n4511, ZN => n1109);
   U2684 : OAI22_X1 port map( A1 => n4064, A2 => n4503, B1 => n4000, B2 => 
                           n4511, ZN => n1090);
   U2685 : OAI22_X1 port map( A1 => n4035, A2 => n4563, B1 => n3971, B2 => 
                           n4571, ZN => n1006);
   U2686 : OAI22_X1 port map( A1 => n4036, A2 => n4563, B1 => n3972, B2 => 
                           n4571, ZN => n984);
   U2687 : OAI22_X1 port map( A1 => n4037, A2 => n4563, B1 => n3973, B2 => 
                           n4571, ZN => n965);
   U2688 : OAI22_X1 port map( A1 => n4038, A2 => n4563, B1 => n3974, B2 => 
                           n4571, ZN => n946);
   U2689 : OAI22_X1 port map( A1 => n4039, A2 => n4563, B1 => n3975, B2 => 
                           n4571, ZN => n927);
   U2690 : OAI22_X1 port map( A1 => n4040, A2 => n4563, B1 => n3976, B2 => 
                           n4571, ZN => n908);
   U2691 : OAI22_X1 port map( A1 => n4041, A2 => n4564, B1 => n3977, B2 => 
                           n4572, ZN => n889);
   U2692 : OAI22_X1 port map( A1 => n4042, A2 => n4564, B1 => n3978, B2 => 
                           n4572, ZN => n870);
   U2693 : OAI22_X1 port map( A1 => n4043, A2 => n4564, B1 => n3979, B2 => 
                           n4572, ZN => n851);
   U2694 : OAI22_X1 port map( A1 => n4044, A2 => n4564, B1 => n3980, B2 => 
                           n4572, ZN => n832);
   U2695 : OAI22_X1 port map( A1 => n4045, A2 => n4564, B1 => n3981, B2 => 
                           n4572, ZN => n813);
   U2696 : OAI22_X1 port map( A1 => n4046, A2 => n4564, B1 => n3982, B2 => 
                           n4572, ZN => n794);
   U2697 : OAI22_X1 port map( A1 => n4047, A2 => n4565, B1 => n3983, B2 => 
                           n4573, ZN => n775);
   U2698 : OAI22_X1 port map( A1 => n4048, A2 => n4565, B1 => n3984, B2 => 
                           n4573, ZN => n756);
   U2699 : OAI22_X1 port map( A1 => n4049, A2 => n4565, B1 => n3985, B2 => 
                           n4573, ZN => n737);
   U2700 : OAI22_X1 port map( A1 => n4050, A2 => n4565, B1 => n3986, B2 => 
                           n4573, ZN => n718);
   U2701 : OAI22_X1 port map( A1 => n4051, A2 => n4565, B1 => n3987, B2 => 
                           n4573, ZN => n699);
   U2702 : OAI22_X1 port map( A1 => n4052, A2 => n4565, B1 => n3988, B2 => 
                           n4573, ZN => n680);
   U2703 : OAI22_X1 port map( A1 => n4053, A2 => n4566, B1 => n3989, B2 => 
                           n4574, ZN => n661);
   U2704 : OAI22_X1 port map( A1 => n4054, A2 => n4566, B1 => n3990, B2 => 
                           n4574, ZN => n642);
   U2705 : OAI22_X1 port map( A1 => n4055, A2 => n4566, B1 => n3991, B2 => 
                           n4574, ZN => n623);
   U2706 : OAI22_X1 port map( A1 => n4056, A2 => n4566, B1 => n3992, B2 => 
                           n4574, ZN => n604);
   U2707 : OAI22_X1 port map( A1 => n4057, A2 => n4566, B1 => n3993, B2 => 
                           n4574, ZN => n585);
   U2708 : OAI22_X1 port map( A1 => n4058, A2 => n4566, B1 => n3994, B2 => 
                           n4574, ZN => n566);
   U2709 : OAI22_X1 port map( A1 => n4059, A2 => n4567, B1 => n3995, B2 => 
                           n4575, ZN => n547);
   U2710 : OAI22_X1 port map( A1 => n4060, A2 => n4567, B1 => n3996, B2 => 
                           n4575, ZN => n528);
   U2711 : OAI22_X1 port map( A1 => n4061, A2 => n4567, B1 => n3997, B2 => 
                           n4575, ZN => n509);
   U2712 : OAI22_X1 port map( A1 => n4062, A2 => n4567, B1 => n3998, B2 => 
                           n4575, ZN => n490);
   U2713 : OAI22_X1 port map( A1 => n4063, A2 => n4567, B1 => n3999, B2 => 
                           n4575, ZN => n471);
   U2714 : OAI22_X1 port map( A1 => n4064, A2 => n4567, B1 => n4000, B2 => 
                           n4575, ZN => n452);
   U2715 : OAI22_X1 port map( A1 => n3073, A2 => n5042, B1 => n1061, B2 => 
                           n5038, ZN => n4129);
   U2716 : NOR4_X1 port map( A1 => n1062, A2 => n1063, A3 => n1064, A4 => n1065
                           , ZN => n1061);
   U2717 : OAI221_X1 port map( B1 => n3297, B2 => n4998, C1 => n3105, C2 => 
                           n4994, A => n1078, ZN => n1063);
   U2718 : OAI221_X1 port map( B1 => n3201, B2 => n4982, C1 => n3233, C2 => 
                           n4978, A => n1079, ZN => n1062);
   U2719 : OAI22_X1 port map( A1 => n3074, A2 => n5042, B1 => n1023, B2 => 
                           n5038, ZN => n4130);
   U2720 : NOR4_X1 port map( A1 => n1025, A2 => n1026, A3 => n1027, A4 => n1028
                           , ZN => n1023);
   U2721 : OAI221_X1 port map( B1 => n3298, B2 => n4998, C1 => n3106, C2 => 
                           n4994, A => n1052, ZN => n1026);
   U2722 : OAI221_X1 port map( B1 => n3202, B2 => n4982, C1 => n3234, C2 => 
                           n4978, A => n1057, ZN => n1025);
   U2723 : OAI22_X1 port map( A1 => n3681, A2 => n4488, B1 => n3617, B2 => 
                           n4496, ZN => n1076);
   U2724 : OAI22_X1 port map( A1 => n3682, A2 => n4488, B1 => n3618, B2 => 
                           n4496, ZN => n1043);
   U2725 : OAI22_X1 port map( A1 => n3041, A2 => n5122, B1 => n423, B2 => n5118
                           , ZN => n4161);
   U2726 : NOR4_X1 port map( A1 => n424, A2 => n425, A3 => n426, A4 => n427, ZN
                           => n423);
   U2727 : OAI221_X1 port map( B1 => n3201, B2 => n5062, C1 => n3233, C2 => 
                           n5058, A => n441, ZN => n424);
   U2728 : OAI221_X1 port map( B1 => n3297, B2 => n5078, C1 => n3105, C2 => 
                           n5074, A => n440, ZN => n425);
   U2729 : OAI22_X1 port map( A1 => n3042, A2 => n5122, B1 => n385, B2 => n5118
                           , ZN => n4162);
   U2730 : NOR4_X1 port map( A1 => n387, A2 => n388, A3 => n389, A4 => n390, ZN
                           => n385);
   U2731 : OAI221_X1 port map( B1 => n3202, B2 => n5062, C1 => n3234, C2 => 
                           n5058, A => n419, ZN => n387);
   U2732 : OAI221_X1 port map( B1 => n3298, B2 => n5078, C1 => n3106, C2 => 
                           n5074, A => n414, ZN => n388);
   U2733 : OAI22_X1 port map( A1 => n3681, A2 => n4552, B1 => n3617, B2 => 
                           n4560, ZN => n438);
   U2734 : OAI22_X1 port map( A1 => n3682, A2 => n4552, B1 => n3618, B2 => 
                           n4560, ZN => n405);
   U2735 : OAI22_X1 port map( A1 => n3809, A2 => n4504, B1 => n3745, B2 => 
                           n4512, ZN => n1075);
   U2736 : OAI22_X1 port map( A1 => n3810, A2 => n4504, B1 => n3746, B2 => 
                           n4512, ZN => n1042);
   U2737 : OAI22_X1 port map( A1 => n3809, A2 => n4568, B1 => n3745, B2 => 
                           n4576, ZN => n437);
   U2738 : OAI22_X1 port map( A1 => n3810, A2 => n4568, B1 => n3746, B2 => 
                           n4576, ZN => n404);
   U2739 : NOR3_X1 port map( A1 => n5136, A2 => ADD_RD2(0), A3 => n5137, ZN => 
                           n2676);
   U2740 : OAI22_X1 port map( A1 => n3683, A2 => n4515, B1 => n3619, B2 => 
                           n4523, ZN => n2671);
   U2741 : OAI22_X1 port map( A1 => n3684, A2 => n4515, B1 => n3620, B2 => 
                           n4523, ZN => n2649);
   U2742 : OAI22_X1 port map( A1 => n3685, A2 => n4515, B1 => n3621, B2 => 
                           n4523, ZN => n2630);
   U2743 : OAI22_X1 port map( A1 => n3686, A2 => n4515, B1 => n3622, B2 => 
                           n4523, ZN => n2611);
   U2744 : OAI22_X1 port map( A1 => n3687, A2 => n4515, B1 => n3623, B2 => 
                           n4523, ZN => n2592);
   U2745 : OAI22_X1 port map( A1 => n3688, A2 => n4515, B1 => n3624, B2 => 
                           n4523, ZN => n2573);
   U2746 : OAI22_X1 port map( A1 => n3689, A2 => n4516, B1 => n3625, B2 => 
                           n4524, ZN => n2554);
   U2747 : OAI22_X1 port map( A1 => n3690, A2 => n4516, B1 => n3626, B2 => 
                           n4524, ZN => n2535);
   U2748 : OAI22_X1 port map( A1 => n3691, A2 => n4516, B1 => n3627, B2 => 
                           n4524, ZN => n2516);
   U2749 : OAI22_X1 port map( A1 => n3692, A2 => n4516, B1 => n3628, B2 => 
                           n4524, ZN => n2497);
   U2750 : OAI22_X1 port map( A1 => n3693, A2 => n4516, B1 => n3629, B2 => 
                           n4524, ZN => n2478);
   U2751 : OAI22_X1 port map( A1 => n3694, A2 => n4516, B1 => n3630, B2 => 
                           n4524, ZN => n2459);
   U2752 : OAI22_X1 port map( A1 => n3695, A2 => n4517, B1 => n3631, B2 => 
                           n4525, ZN => n2440);
   U2753 : OAI22_X1 port map( A1 => n3696, A2 => n4517, B1 => n3632, B2 => 
                           n4525, ZN => n2421);
   U2754 : OAI22_X1 port map( A1 => n3697, A2 => n4517, B1 => n3633, B2 => 
                           n4525, ZN => n2402);
   U2755 : OAI22_X1 port map( A1 => n3698, A2 => n4517, B1 => n3634, B2 => 
                           n4525, ZN => n2383);
   U2756 : OAI22_X1 port map( A1 => n3699, A2 => n4517, B1 => n3635, B2 => 
                           n4525, ZN => n2364);
   U2757 : OAI22_X1 port map( A1 => n3700, A2 => n4517, B1 => n3636, B2 => 
                           n4525, ZN => n2345);
   U2758 : OAI22_X1 port map( A1 => n3701, A2 => n4518, B1 => n3637, B2 => 
                           n4526, ZN => n1302);
   U2759 : OAI22_X1 port map( A1 => n3702, A2 => n4518, B1 => n3638, B2 => 
                           n4526, ZN => n1283);
   U2760 : OAI22_X1 port map( A1 => n3703, A2 => n4518, B1 => n3639, B2 => 
                           n4526, ZN => n1264);
   U2761 : OAI22_X1 port map( A1 => n3704, A2 => n4518, B1 => n3640, B2 => 
                           n4526, ZN => n1245);
   U2762 : OAI22_X1 port map( A1 => n3705, A2 => n4518, B1 => n3641, B2 => 
                           n4526, ZN => n1226);
   U2763 : OAI22_X1 port map( A1 => n3706, A2 => n4518, B1 => n3642, B2 => 
                           n4526, ZN => n1207);
   U2764 : OAI22_X1 port map( A1 => n3707, A2 => n4519, B1 => n3643, B2 => 
                           n4527, ZN => n1188);
   U2765 : OAI22_X1 port map( A1 => n3708, A2 => n4519, B1 => n3644, B2 => 
                           n4527, ZN => n1169);
   U2766 : OAI22_X1 port map( A1 => n3709, A2 => n4519, B1 => n3645, B2 => 
                           n4527, ZN => n1150);
   U2767 : OAI22_X1 port map( A1 => n3710, A2 => n4519, B1 => n3646, B2 => 
                           n4527, ZN => n1131);
   U2768 : OAI22_X1 port map( A1 => n3711, A2 => n4519, B1 => n3647, B2 => 
                           n4527, ZN => n1112);
   U2769 : OAI22_X1 port map( A1 => n3712, A2 => n4519, B1 => n3648, B2 => 
                           n4527, ZN => n1093);
   U2770 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n5137, 
                           ZN => n2677);
   U2771 : OAI22_X1 port map( A1 => n3937, A2 => n4488, B1 => n3873, B2 => 
                           n4496, ZN => n1072);
   U2772 : OAI22_X1 port map( A1 => n3938, A2 => n4488, B1 => n3874, B2 => 
                           n4496, ZN => n1039);
   U2773 : OAI22_X1 port map( A1 => n3937, A2 => n4552, B1 => n3873, B2 => 
                           n4560, ZN => n434);
   U2774 : OAI22_X1 port map( A1 => n3938, A2 => n4552, B1 => n3874, B2 => 
                           n4560, ZN => n401);
   U2775 : OAI22_X1 port map( A1 => n4065, A2 => n4504, B1 => n4001, B2 => 
                           n4512, ZN => n1071);
   U2776 : OAI22_X1 port map( A1 => n4066, A2 => n4504, B1 => n4002, B2 => 
                           n4512, ZN => n1038);
   U2777 : OAI22_X1 port map( A1 => n4065, A2 => n4568, B1 => n4001, B2 => 
                           n4576, ZN => n433);
   U2778 : OAI22_X1 port map( A1 => n4066, A2 => n4568, B1 => n4002, B2 => 
                           n4576, ZN => n400);
   U2779 : NOR3_X1 port map( A1 => n5149, A2 => ADD_RD1(0), A3 => n5150, ZN => 
                           n1014);
   U2780 : OAI22_X1 port map( A1 => n3683, A2 => n4579, B1 => n3619, B2 => 
                           n4587, ZN => n1009);
   U2781 : OAI22_X1 port map( A1 => n3684, A2 => n4579, B1 => n3620, B2 => 
                           n4587, ZN => n987);
   U2782 : OAI22_X1 port map( A1 => n3685, A2 => n4579, B1 => n3621, B2 => 
                           n4587, ZN => n968);
   U2783 : OAI22_X1 port map( A1 => n3686, A2 => n4579, B1 => n3622, B2 => 
                           n4587, ZN => n949);
   U2784 : OAI22_X1 port map( A1 => n3687, A2 => n4579, B1 => n3623, B2 => 
                           n4587, ZN => n930);
   U2785 : OAI22_X1 port map( A1 => n3688, A2 => n4579, B1 => n3624, B2 => 
                           n4587, ZN => n911);
   U2786 : OAI22_X1 port map( A1 => n3689, A2 => n4580, B1 => n3625, B2 => 
                           n4588, ZN => n892);
   U2787 : OAI22_X1 port map( A1 => n3690, A2 => n4580, B1 => n3626, B2 => 
                           n4588, ZN => n873);
   U2788 : OAI22_X1 port map( A1 => n3691, A2 => n4580, B1 => n3627, B2 => 
                           n4588, ZN => n854);
   U2789 : OAI22_X1 port map( A1 => n3692, A2 => n4580, B1 => n3628, B2 => 
                           n4588, ZN => n835);
   U2790 : OAI22_X1 port map( A1 => n3693, A2 => n4580, B1 => n3629, B2 => 
                           n4588, ZN => n816);
   U2791 : OAI22_X1 port map( A1 => n3694, A2 => n4580, B1 => n3630, B2 => 
                           n4588, ZN => n797);
   U2792 : OAI22_X1 port map( A1 => n3695, A2 => n4581, B1 => n3631, B2 => 
                           n4589, ZN => n778);
   U2793 : OAI22_X1 port map( A1 => n3696, A2 => n4581, B1 => n3632, B2 => 
                           n4589, ZN => n759);
   U2794 : OAI22_X1 port map( A1 => n3697, A2 => n4581, B1 => n3633, B2 => 
                           n4589, ZN => n740);
   U2795 : OAI22_X1 port map( A1 => n3698, A2 => n4581, B1 => n3634, B2 => 
                           n4589, ZN => n721);
   U2796 : OAI22_X1 port map( A1 => n3699, A2 => n4581, B1 => n3635, B2 => 
                           n4589, ZN => n702);
   U2797 : OAI22_X1 port map( A1 => n3700, A2 => n4581, B1 => n3636, B2 => 
                           n4589, ZN => n683);
   U2798 : OAI22_X1 port map( A1 => n3701, A2 => n4582, B1 => n3637, B2 => 
                           n4590, ZN => n664);
   U2799 : OAI22_X1 port map( A1 => n3702, A2 => n4582, B1 => n3638, B2 => 
                           n4590, ZN => n645);
   U2800 : OAI22_X1 port map( A1 => n3703, A2 => n4582, B1 => n3639, B2 => 
                           n4590, ZN => n626);
   U2801 : OAI22_X1 port map( A1 => n3704, A2 => n4582, B1 => n3640, B2 => 
                           n4590, ZN => n607);
   U2802 : OAI22_X1 port map( A1 => n3705, A2 => n4582, B1 => n3641, B2 => 
                           n4590, ZN => n588);
   U2803 : OAI22_X1 port map( A1 => n3706, A2 => n4582, B1 => n3642, B2 => 
                           n4590, ZN => n569);
   U2804 : OAI22_X1 port map( A1 => n3707, A2 => n4583, B1 => n3643, B2 => 
                           n4591, ZN => n550);
   U2805 : OAI22_X1 port map( A1 => n3708, A2 => n4583, B1 => n3644, B2 => 
                           n4591, ZN => n531);
   U2806 : OAI22_X1 port map( A1 => n3709, A2 => n4583, B1 => n3645, B2 => 
                           n4591, ZN => n512);
   U2807 : OAI22_X1 port map( A1 => n3710, A2 => n4583, B1 => n3646, B2 => 
                           n4591, ZN => n493);
   U2808 : OAI22_X1 port map( A1 => n3711, A2 => n4583, B1 => n3647, B2 => 
                           n4591, ZN => n474);
   U2809 : OAI22_X1 port map( A1 => n3712, A2 => n4583, B1 => n3648, B2 => 
                           n4591, ZN => n455);
   U2810 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n5150, 
                           ZN => n1015);
   U2811 : OAI22_X1 port map( A1 => n3939, A2 => n4515, B1 => n3875, B2 => 
                           n4523, ZN => n2667);
   U2812 : OAI22_X1 port map( A1 => n3940, A2 => n4515, B1 => n3876, B2 => 
                           n4523, ZN => n2645);
   U2813 : OAI22_X1 port map( A1 => n3941, A2 => n4515, B1 => n3877, B2 => 
                           n4523, ZN => n2626);
   U2814 : OAI22_X1 port map( A1 => n3942, A2 => n4515, B1 => n3878, B2 => 
                           n4523, ZN => n2607);
   U2815 : OAI22_X1 port map( A1 => n3943, A2 => n4515, B1 => n3879, B2 => 
                           n4523, ZN => n2588);
   U2816 : OAI22_X1 port map( A1 => n3944, A2 => n4515, B1 => n3880, B2 => 
                           n4523, ZN => n2569);
   U2817 : OAI22_X1 port map( A1 => n3945, A2 => n4516, B1 => n3881, B2 => 
                           n4524, ZN => n2550);
   U2818 : OAI22_X1 port map( A1 => n3946, A2 => n4516, B1 => n3882, B2 => 
                           n4524, ZN => n2531);
   U2819 : OAI22_X1 port map( A1 => n3947, A2 => n4516, B1 => n3883, B2 => 
                           n4524, ZN => n2512);
   U2820 : OAI22_X1 port map( A1 => n3948, A2 => n4516, B1 => n3884, B2 => 
                           n4524, ZN => n2493);
   U2821 : OAI22_X1 port map( A1 => n3949, A2 => n4516, B1 => n3885, B2 => 
                           n4524, ZN => n2474);
   U2822 : OAI22_X1 port map( A1 => n3950, A2 => n4516, B1 => n3886, B2 => 
                           n4524, ZN => n2455);
   U2823 : OAI22_X1 port map( A1 => n3951, A2 => n4517, B1 => n3887, B2 => 
                           n4525, ZN => n2436);
   U2824 : OAI22_X1 port map( A1 => n3952, A2 => n4517, B1 => n3888, B2 => 
                           n4525, ZN => n2417);
   U2825 : OAI22_X1 port map( A1 => n3953, A2 => n4517, B1 => n3889, B2 => 
                           n4525, ZN => n2398);
   U2826 : OAI22_X1 port map( A1 => n3954, A2 => n4517, B1 => n3890, B2 => 
                           n4525, ZN => n2379);
   U2827 : OAI22_X1 port map( A1 => n3955, A2 => n4517, B1 => n3891, B2 => 
                           n4525, ZN => n2360);
   U2828 : OAI22_X1 port map( A1 => n3956, A2 => n4517, B1 => n3892, B2 => 
                           n4525, ZN => n2341);
   U2829 : OAI22_X1 port map( A1 => n3957, A2 => n4518, B1 => n3893, B2 => 
                           n4526, ZN => n1298);
   U2830 : OAI22_X1 port map( A1 => n3958, A2 => n4518, B1 => n3894, B2 => 
                           n4526, ZN => n1279);
   U2831 : OAI22_X1 port map( A1 => n3959, A2 => n4518, B1 => n3895, B2 => 
                           n4526, ZN => n1260);
   U2832 : OAI22_X1 port map( A1 => n3960, A2 => n4518, B1 => n3896, B2 => 
                           n4526, ZN => n1241);
   U2833 : OAI22_X1 port map( A1 => n3961, A2 => n4518, B1 => n3897, B2 => 
                           n4526, ZN => n1222);
   U2834 : OAI22_X1 port map( A1 => n3962, A2 => n4518, B1 => n3898, B2 => 
                           n4526, ZN => n1203);
   U2835 : OAI22_X1 port map( A1 => n3963, A2 => n4519, B1 => n3899, B2 => 
                           n4527, ZN => n1184);
   U2836 : OAI22_X1 port map( A1 => n3964, A2 => n4519, B1 => n3900, B2 => 
                           n4527, ZN => n1165);
   U2837 : OAI22_X1 port map( A1 => n3965, A2 => n4519, B1 => n3901, B2 => 
                           n4527, ZN => n1146);
   U2838 : OAI22_X1 port map( A1 => n3966, A2 => n4519, B1 => n3902, B2 => 
                           n4527, ZN => n1127);
   U2839 : OAI22_X1 port map( A1 => n3967, A2 => n4519, B1 => n3903, B2 => 
                           n4527, ZN => n1108);
   U2840 : OAI22_X1 port map( A1 => n3968, A2 => n4519, B1 => n3904, B2 => 
                           n4527, ZN => n1089);
   U2841 : OAI22_X1 port map( A1 => n3713, A2 => n4520, B1 => n3649, B2 => 
                           n4528, ZN => n1074);
   U2842 : OAI22_X1 port map( A1 => n3714, A2 => n4520, B1 => n3650, B2 => 
                           n4528, ZN => n1041);
   U2843 : OAI22_X1 port map( A1 => n3939, A2 => n4579, B1 => n3875, B2 => 
                           n4587, ZN => n1005);
   U2844 : OAI22_X1 port map( A1 => n3940, A2 => n4579, B1 => n3876, B2 => 
                           n4587, ZN => n983);
   U2845 : OAI22_X1 port map( A1 => n3941, A2 => n4579, B1 => n3877, B2 => 
                           n4587, ZN => n964);
   U2846 : OAI22_X1 port map( A1 => n3942, A2 => n4579, B1 => n3878, B2 => 
                           n4587, ZN => n945);
   U2847 : OAI22_X1 port map( A1 => n3943, A2 => n4579, B1 => n3879, B2 => 
                           n4587, ZN => n926);
   U2848 : OAI22_X1 port map( A1 => n3944, A2 => n4579, B1 => n3880, B2 => 
                           n4587, ZN => n907);
   U2849 : OAI22_X1 port map( A1 => n3945, A2 => n4580, B1 => n3881, B2 => 
                           n4588, ZN => n888);
   U2850 : OAI22_X1 port map( A1 => n3946, A2 => n4580, B1 => n3882, B2 => 
                           n4588, ZN => n869);
   U2851 : OAI22_X1 port map( A1 => n3947, A2 => n4580, B1 => n3883, B2 => 
                           n4588, ZN => n850);
   U2852 : OAI22_X1 port map( A1 => n3948, A2 => n4580, B1 => n3884, B2 => 
                           n4588, ZN => n831);
   U2853 : OAI22_X1 port map( A1 => n3949, A2 => n4580, B1 => n3885, B2 => 
                           n4588, ZN => n812);
   U2854 : OAI22_X1 port map( A1 => n3950, A2 => n4580, B1 => n3886, B2 => 
                           n4588, ZN => n793);
   U2855 : OAI22_X1 port map( A1 => n3951, A2 => n4581, B1 => n3887, B2 => 
                           n4589, ZN => n774);
   U2856 : OAI22_X1 port map( A1 => n3952, A2 => n4581, B1 => n3888, B2 => 
                           n4589, ZN => n755);
   U2857 : OAI22_X1 port map( A1 => n3953, A2 => n4581, B1 => n3889, B2 => 
                           n4589, ZN => n736);
   U2858 : OAI22_X1 port map( A1 => n3954, A2 => n4581, B1 => n3890, B2 => 
                           n4589, ZN => n717);
   U2859 : OAI22_X1 port map( A1 => n3955, A2 => n4581, B1 => n3891, B2 => 
                           n4589, ZN => n698);
   U2860 : OAI22_X1 port map( A1 => n3956, A2 => n4581, B1 => n3892, B2 => 
                           n4589, ZN => n679);
   U2861 : OAI22_X1 port map( A1 => n3957, A2 => n4582, B1 => n3893, B2 => 
                           n4590, ZN => n660);
   U2862 : OAI22_X1 port map( A1 => n3958, A2 => n4582, B1 => n3894, B2 => 
                           n4590, ZN => n641);
   U2863 : OAI22_X1 port map( A1 => n3959, A2 => n4582, B1 => n3895, B2 => 
                           n4590, ZN => n622);
   U2864 : OAI22_X1 port map( A1 => n3960, A2 => n4582, B1 => n3896, B2 => 
                           n4590, ZN => n603);
   U2865 : OAI22_X1 port map( A1 => n3961, A2 => n4582, B1 => n3897, B2 => 
                           n4590, ZN => n584);
   U2866 : OAI22_X1 port map( A1 => n3962, A2 => n4582, B1 => n3898, B2 => 
                           n4590, ZN => n565);
   U2867 : OAI22_X1 port map( A1 => n3963, A2 => n4583, B1 => n3899, B2 => 
                           n4591, ZN => n546);
   U2868 : OAI22_X1 port map( A1 => n3964, A2 => n4583, B1 => n3900, B2 => 
                           n4591, ZN => n527);
   U2869 : OAI22_X1 port map( A1 => n3965, A2 => n4583, B1 => n3901, B2 => 
                           n4591, ZN => n508);
   U2870 : OAI22_X1 port map( A1 => n3966, A2 => n4583, B1 => n3902, B2 => 
                           n4591, ZN => n489);
   U2871 : OAI22_X1 port map( A1 => n3967, A2 => n4583, B1 => n3903, B2 => 
                           n4591, ZN => n470);
   U2872 : OAI22_X1 port map( A1 => n3968, A2 => n4583, B1 => n3904, B2 => 
                           n4591, ZN => n451);
   U2873 : OAI22_X1 port map( A1 => n3713, A2 => n4584, B1 => n3649, B2 => 
                           n4592, ZN => n436);
   U2874 : OAI22_X1 port map( A1 => n3714, A2 => n4584, B1 => n3650, B2 => 
                           n4592, ZN => n403);
   U2875 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n2709);
   U2876 : OAI22_X1 port map( A1 => n3969, A2 => n4520, B1 => n3905, B2 => 
                           n4528, ZN => n1070);
   U2877 : OAI22_X1 port map( A1 => n3970, A2 => n4520, B1 => n3906, B2 => 
                           n4528, ZN => n1037);
   U2878 : OAI22_X1 port map( A1 => n3969, A2 => n4584, B1 => n3905, B2 => 
                           n4592, ZN => n432);
   U2879 : OAI22_X1 port map( A1 => n3970, A2 => n4584, B1 => n3906, B2 => 
                           n4592, ZN => n399);
   U2880 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n5136, 
                           ZN => n2678);
   U2881 : OAI22_X1 port map( A1 => n3811, A2 => n4539, B1 => n3747, B2 => 
                           n4531, ZN => n2670);
   U2882 : OAI22_X1 port map( A1 => n3812, A2 => n4539, B1 => n3748, B2 => 
                           n4531, ZN => n2648);
   U2883 : OAI22_X1 port map( A1 => n3813, A2 => n4539, B1 => n3749, B2 => 
                           n4531, ZN => n2629);
   U2884 : OAI22_X1 port map( A1 => n3814, A2 => n4539, B1 => n3750, B2 => 
                           n4531, ZN => n2610);
   U2885 : OAI22_X1 port map( A1 => n3815, A2 => n4539, B1 => n3751, B2 => 
                           n4531, ZN => n2591);
   U2886 : OAI22_X1 port map( A1 => n3816, A2 => n4539, B1 => n3752, B2 => 
                           n4531, ZN => n2572);
   U2887 : OAI22_X1 port map( A1 => n3817, A2 => n4540, B1 => n3753, B2 => 
                           n4532, ZN => n2553);
   U2888 : OAI22_X1 port map( A1 => n3818, A2 => n4540, B1 => n3754, B2 => 
                           n4532, ZN => n2534);
   U2889 : OAI22_X1 port map( A1 => n3819, A2 => n4540, B1 => n3755, B2 => 
                           n4532, ZN => n2515);
   U2890 : OAI22_X1 port map( A1 => n3820, A2 => n4540, B1 => n3756, B2 => 
                           n4532, ZN => n2496);
   U2891 : OAI22_X1 port map( A1 => n3821, A2 => n4540, B1 => n3757, B2 => 
                           n4532, ZN => n2477);
   U2892 : OAI22_X1 port map( A1 => n3822, A2 => n4540, B1 => n3758, B2 => 
                           n4532, ZN => n2458);
   U2893 : OAI22_X1 port map( A1 => n3823, A2 => n4541, B1 => n3759, B2 => 
                           n4533, ZN => n2439);
   U2894 : OAI22_X1 port map( A1 => n3824, A2 => n4541, B1 => n3760, B2 => 
                           n4533, ZN => n2420);
   U2895 : OAI22_X1 port map( A1 => n3825, A2 => n4541, B1 => n3761, B2 => 
                           n4533, ZN => n2401);
   U2896 : OAI22_X1 port map( A1 => n3826, A2 => n4541, B1 => n3762, B2 => 
                           n4533, ZN => n2382);
   U2897 : OAI22_X1 port map( A1 => n3827, A2 => n4541, B1 => n3763, B2 => 
                           n4533, ZN => n2363);
   U2898 : OAI22_X1 port map( A1 => n3828, A2 => n4541, B1 => n3764, B2 => 
                           n4533, ZN => n2344);
   U2899 : OAI22_X1 port map( A1 => n3829, A2 => n4542, B1 => n3765, B2 => 
                           n4534, ZN => n1301);
   U2900 : OAI22_X1 port map( A1 => n3830, A2 => n4542, B1 => n3766, B2 => 
                           n4534, ZN => n1282);
   U2901 : OAI22_X1 port map( A1 => n3831, A2 => n4542, B1 => n3767, B2 => 
                           n4534, ZN => n1263);
   U2902 : OAI22_X1 port map( A1 => n3832, A2 => n4542, B1 => n3768, B2 => 
                           n4534, ZN => n1244);
   U2903 : OAI22_X1 port map( A1 => n3833, A2 => n4542, B1 => n3769, B2 => 
                           n4534, ZN => n1225);
   U2904 : OAI22_X1 port map( A1 => n3834, A2 => n4542, B1 => n3770, B2 => 
                           n4534, ZN => n1206);
   U2905 : OAI22_X1 port map( A1 => n3835, A2 => n4543, B1 => n3771, B2 => 
                           n4535, ZN => n1187);
   U2906 : OAI22_X1 port map( A1 => n3836, A2 => n4543, B1 => n3772, B2 => 
                           n4535, ZN => n1168);
   U2907 : OAI22_X1 port map( A1 => n3837, A2 => n4543, B1 => n3773, B2 => 
                           n4535, ZN => n1149);
   U2908 : OAI22_X1 port map( A1 => n3838, A2 => n4543, B1 => n3774, B2 => 
                           n4535, ZN => n1130);
   U2909 : OAI22_X1 port map( A1 => n3839, A2 => n4543, B1 => n3775, B2 => 
                           n4535, ZN => n1111);
   U2910 : OAI22_X1 port map( A1 => n3840, A2 => n4543, B1 => n3776, B2 => 
                           n4535, ZN => n1092);
   U2911 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n5149, 
                           ZN => n1016);
   U2912 : OAI22_X1 port map( A1 => n3811, A2 => n4603, B1 => n3747, B2 => 
                           n4595, ZN => n1008);
   U2913 : OAI22_X1 port map( A1 => n3812, A2 => n4603, B1 => n3748, B2 => 
                           n4595, ZN => n986);
   U2914 : OAI22_X1 port map( A1 => n3813, A2 => n4603, B1 => n3749, B2 => 
                           n4595, ZN => n967);
   U2915 : OAI22_X1 port map( A1 => n3814, A2 => n4603, B1 => n3750, B2 => 
                           n4595, ZN => n948);
   U2916 : OAI22_X1 port map( A1 => n3815, A2 => n4603, B1 => n3751, B2 => 
                           n4595, ZN => n929);
   U2917 : OAI22_X1 port map( A1 => n3816, A2 => n4603, B1 => n3752, B2 => 
                           n4595, ZN => n910);
   U2918 : OAI22_X1 port map( A1 => n3817, A2 => n4604, B1 => n3753, B2 => 
                           n4596, ZN => n891);
   U2919 : OAI22_X1 port map( A1 => n3818, A2 => n4604, B1 => n3754, B2 => 
                           n4596, ZN => n872);
   U2920 : OAI22_X1 port map( A1 => n3819, A2 => n4604, B1 => n3755, B2 => 
                           n4596, ZN => n853);
   U2921 : OAI22_X1 port map( A1 => n3820, A2 => n4604, B1 => n3756, B2 => 
                           n4596, ZN => n834);
   U2922 : OAI22_X1 port map( A1 => n3821, A2 => n4604, B1 => n3757, B2 => 
                           n4596, ZN => n815);
   U2923 : OAI22_X1 port map( A1 => n3822, A2 => n4604, B1 => n3758, B2 => 
                           n4596, ZN => n796);
   U2924 : OAI22_X1 port map( A1 => n3823, A2 => n4605, B1 => n3759, B2 => 
                           n4597, ZN => n777);
   U2925 : OAI22_X1 port map( A1 => n3824, A2 => n4605, B1 => n3760, B2 => 
                           n4597, ZN => n758);
   U2926 : OAI22_X1 port map( A1 => n3825, A2 => n4605, B1 => n3761, B2 => 
                           n4597, ZN => n739);
   U2927 : OAI22_X1 port map( A1 => n3826, A2 => n4605, B1 => n3762, B2 => 
                           n4597, ZN => n720);
   U2928 : OAI22_X1 port map( A1 => n3827, A2 => n4605, B1 => n3763, B2 => 
                           n4597, ZN => n701);
   U2929 : OAI22_X1 port map( A1 => n3828, A2 => n4605, B1 => n3764, B2 => 
                           n4597, ZN => n682);
   U2930 : OAI22_X1 port map( A1 => n3829, A2 => n4606, B1 => n3765, B2 => 
                           n4598, ZN => n663);
   U2931 : OAI22_X1 port map( A1 => n3830, A2 => n4606, B1 => n3766, B2 => 
                           n4598, ZN => n644);
   U2932 : OAI22_X1 port map( A1 => n3831, A2 => n4606, B1 => n3767, B2 => 
                           n4598, ZN => n625);
   U2933 : OAI22_X1 port map( A1 => n3832, A2 => n4606, B1 => n3768, B2 => 
                           n4598, ZN => n606);
   U2934 : OAI22_X1 port map( A1 => n3833, A2 => n4606, B1 => n3769, B2 => 
                           n4598, ZN => n587);
   U2935 : OAI22_X1 port map( A1 => n3834, A2 => n4606, B1 => n3770, B2 => 
                           n4598, ZN => n568);
   U2936 : OAI22_X1 port map( A1 => n3835, A2 => n4607, B1 => n3771, B2 => 
                           n4599, ZN => n549);
   U2937 : OAI22_X1 port map( A1 => n3836, A2 => n4607, B1 => n3772, B2 => 
                           n4599, ZN => n530);
   U2938 : OAI22_X1 port map( A1 => n3837, A2 => n4607, B1 => n3773, B2 => 
                           n4599, ZN => n511);
   U2939 : OAI22_X1 port map( A1 => n3838, A2 => n4607, B1 => n3774, B2 => 
                           n4599, ZN => n492);
   U2940 : OAI22_X1 port map( A1 => n3839, A2 => n4607, B1 => n3775, B2 => 
                           n4599, ZN => n473);
   U2941 : OAI22_X1 port map( A1 => n3840, A2 => n4607, B1 => n3776, B2 => 
                           n4599, ZN => n454);
   U2942 : OAI22_X1 port map( A1 => n4067, A2 => n4539, B1 => n4003, B2 => 
                           n4531, ZN => n2666);
   U2943 : OAI22_X1 port map( A1 => n4068, A2 => n4539, B1 => n4004, B2 => 
                           n4531, ZN => n2644);
   U2944 : OAI22_X1 port map( A1 => n4069, A2 => n4539, B1 => n4005, B2 => 
                           n4531, ZN => n2625);
   U2945 : OAI22_X1 port map( A1 => n4070, A2 => n4539, B1 => n4006, B2 => 
                           n4531, ZN => n2606);
   U2946 : OAI22_X1 port map( A1 => n4071, A2 => n4539, B1 => n4007, B2 => 
                           n4531, ZN => n2587);
   U2947 : OAI22_X1 port map( A1 => n4072, A2 => n4539, B1 => n4008, B2 => 
                           n4531, ZN => n2568);
   U2948 : OAI22_X1 port map( A1 => n4073, A2 => n4540, B1 => n4009, B2 => 
                           n4532, ZN => n2549);
   U2949 : OAI22_X1 port map( A1 => n4074, A2 => n4540, B1 => n4010, B2 => 
                           n4532, ZN => n2530);
   U2950 : OAI22_X1 port map( A1 => n4075, A2 => n4540, B1 => n4011, B2 => 
                           n4532, ZN => n2511);
   U2951 : OAI22_X1 port map( A1 => n4076, A2 => n4540, B1 => n4012, B2 => 
                           n4532, ZN => n2492);
   U2952 : OAI22_X1 port map( A1 => n4077, A2 => n4540, B1 => n4013, B2 => 
                           n4532, ZN => n2473);
   U2953 : OAI22_X1 port map( A1 => n4078, A2 => n4540, B1 => n4014, B2 => 
                           n4532, ZN => n2454);
   U2954 : OAI22_X1 port map( A1 => n4079, A2 => n4541, B1 => n4015, B2 => 
                           n4533, ZN => n2435);
   U2955 : OAI22_X1 port map( A1 => n4080, A2 => n4541, B1 => n4016, B2 => 
                           n4533, ZN => n2416);
   U2956 : OAI22_X1 port map( A1 => n4081, A2 => n4541, B1 => n4017, B2 => 
                           n4533, ZN => n2397);
   U2957 : OAI22_X1 port map( A1 => n4082, A2 => n4541, B1 => n4018, B2 => 
                           n4533, ZN => n2378);
   U2958 : OAI22_X1 port map( A1 => n4083, A2 => n4541, B1 => n4019, B2 => 
                           n4533, ZN => n2359);
   U2959 : OAI22_X1 port map( A1 => n4084, A2 => n4541, B1 => n4020, B2 => 
                           n4533, ZN => n2340);
   U2960 : OAI22_X1 port map( A1 => n4085, A2 => n4542, B1 => n4021, B2 => 
                           n4534, ZN => n1297);
   U2961 : OAI22_X1 port map( A1 => n4086, A2 => n4542, B1 => n4022, B2 => 
                           n4534, ZN => n1278);
   U2962 : OAI22_X1 port map( A1 => n4087, A2 => n4542, B1 => n4023, B2 => 
                           n4534, ZN => n1259);
   U2963 : OAI22_X1 port map( A1 => n4088, A2 => n4542, B1 => n4024, B2 => 
                           n4534, ZN => n1240);
   U2964 : OAI22_X1 port map( A1 => n4089, A2 => n4542, B1 => n4025, B2 => 
                           n4534, ZN => n1221);
   U2965 : OAI22_X1 port map( A1 => n4090, A2 => n4542, B1 => n4026, B2 => 
                           n4534, ZN => n1202);
   U2966 : OAI22_X1 port map( A1 => n4091, A2 => n4543, B1 => n4027, B2 => 
                           n4535, ZN => n1183);
   U2967 : OAI22_X1 port map( A1 => n4092, A2 => n4543, B1 => n4028, B2 => 
                           n4535, ZN => n1164);
   U2968 : OAI22_X1 port map( A1 => n4093, A2 => n4543, B1 => n4029, B2 => 
                           n4535, ZN => n1145);
   U2969 : OAI22_X1 port map( A1 => n4094, A2 => n4543, B1 => n4030, B2 => 
                           n4535, ZN => n1126);
   U2970 : OAI22_X1 port map( A1 => n4095, A2 => n4543, B1 => n4031, B2 => 
                           n4535, ZN => n1107);
   U2971 : OAI22_X1 port map( A1 => n4096, A2 => n4543, B1 => n4032, B2 => 
                           n4535, ZN => n1088);
   U2972 : OAI22_X1 port map( A1 => n4067, A2 => n4603, B1 => n4003, B2 => 
                           n4595, ZN => n1004);
   U2973 : OAI22_X1 port map( A1 => n4068, A2 => n4603, B1 => n4004, B2 => 
                           n4595, ZN => n982);
   U2974 : OAI22_X1 port map( A1 => n4069, A2 => n4603, B1 => n4005, B2 => 
                           n4595, ZN => n963);
   U2975 : OAI22_X1 port map( A1 => n4070, A2 => n4603, B1 => n4006, B2 => 
                           n4595, ZN => n944);
   U2976 : OAI22_X1 port map( A1 => n4071, A2 => n4603, B1 => n4007, B2 => 
                           n4595, ZN => n925);
   U2977 : OAI22_X1 port map( A1 => n4072, A2 => n4603, B1 => n4008, B2 => 
                           n4595, ZN => n906);
   U2978 : OAI22_X1 port map( A1 => n4073, A2 => n4604, B1 => n4009, B2 => 
                           n4596, ZN => n887);
   U2979 : OAI22_X1 port map( A1 => n4074, A2 => n4604, B1 => n4010, B2 => 
                           n4596, ZN => n868);
   U2980 : OAI22_X1 port map( A1 => n4075, A2 => n4604, B1 => n4011, B2 => 
                           n4596, ZN => n849);
   U2981 : OAI22_X1 port map( A1 => n4076, A2 => n4604, B1 => n4012, B2 => 
                           n4596, ZN => n830);
   U2982 : OAI22_X1 port map( A1 => n4077, A2 => n4604, B1 => n4013, B2 => 
                           n4596, ZN => n811);
   U2983 : OAI22_X1 port map( A1 => n4078, A2 => n4604, B1 => n4014, B2 => 
                           n4596, ZN => n792);
   U2984 : OAI22_X1 port map( A1 => n4079, A2 => n4605, B1 => n4015, B2 => 
                           n4597, ZN => n773);
   U2985 : OAI22_X1 port map( A1 => n4080, A2 => n4605, B1 => n4016, B2 => 
                           n4597, ZN => n754);
   U2986 : OAI22_X1 port map( A1 => n4081, A2 => n4605, B1 => n4017, B2 => 
                           n4597, ZN => n735);
   U2987 : OAI22_X1 port map( A1 => n4082, A2 => n4605, B1 => n4018, B2 => 
                           n4597, ZN => n716);
   U2988 : OAI22_X1 port map( A1 => n4083, A2 => n4605, B1 => n4019, B2 => 
                           n4597, ZN => n697);
   U2989 : OAI22_X1 port map( A1 => n4084, A2 => n4605, B1 => n4020, B2 => 
                           n4597, ZN => n678);
   U2990 : OAI22_X1 port map( A1 => n4085, A2 => n4606, B1 => n4021, B2 => 
                           n4598, ZN => n659);
   U2991 : OAI22_X1 port map( A1 => n4086, A2 => n4606, B1 => n4022, B2 => 
                           n4598, ZN => n640);
   U2992 : OAI22_X1 port map( A1 => n4087, A2 => n4606, B1 => n4023, B2 => 
                           n4598, ZN => n621);
   U2993 : OAI22_X1 port map( A1 => n4088, A2 => n4606, B1 => n4024, B2 => 
                           n4598, ZN => n602);
   U2994 : OAI22_X1 port map( A1 => n4089, A2 => n4606, B1 => n4025, B2 => 
                           n4598, ZN => n583);
   U2995 : OAI22_X1 port map( A1 => n4090, A2 => n4606, B1 => n4026, B2 => 
                           n4598, ZN => n564);
   U2996 : OAI22_X1 port map( A1 => n4091, A2 => n4607, B1 => n4027, B2 => 
                           n4599, ZN => n545);
   U2997 : OAI22_X1 port map( A1 => n4092, A2 => n4607, B1 => n4028, B2 => 
                           n4599, ZN => n526);
   U2998 : OAI22_X1 port map( A1 => n4093, A2 => n4607, B1 => n4029, B2 => 
                           n4599, ZN => n507);
   U2999 : OAI22_X1 port map( A1 => n4094, A2 => n4607, B1 => n4030, B2 => 
                           n4599, ZN => n488);
   U3000 : OAI22_X1 port map( A1 => n4095, A2 => n4607, B1 => n4031, B2 => 
                           n4599, ZN => n469);
   U3001 : OAI22_X1 port map( A1 => n4096, A2 => n4607, B1 => n4032, B2 => 
                           n4599, ZN => n450);
   U3002 : OAI22_X1 port map( A1 => n3841, A2 => n4544, B1 => n3777, B2 => 
                           n4536, ZN => n1073);
   U3003 : OAI22_X1 port map( A1 => n3842, A2 => n4544, B1 => n3778, B2 => 
                           n4536, ZN => n1040);
   U3004 : OAI22_X1 port map( A1 => n3841, A2 => n4608, B1 => n3777, B2 => 
                           n4600, ZN => n435);
   U3005 : OAI22_X1 port map( A1 => n3842, A2 => n4608, B1 => n3778, B2 => 
                           n4600, ZN => n402);
   U3006 : OAI22_X1 port map( A1 => n4097, A2 => n4544, B1 => n4033, B2 => 
                           n4536, ZN => n1069);
   U3007 : OAI22_X1 port map( A1 => n4098, A2 => n4544, B1 => n4034, B2 => 
                           n4536, ZN => n1036);
   U3008 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(0), ZN => n1017);
   U3009 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n2679);
   U3010 : OAI22_X1 port map( A1 => n4097, A2 => n4608, B1 => n4033, B2 => 
                           n4600, ZN => n431);
   U3011 : OAI22_X1 port map( A1 => n4098, A2 => n4608, B1 => n4034, B2 => 
                           n4600, ZN => n398);
   U3012 : OAI221_X1 port map( B1 => n3483, B2 => n5018, C1 => n3547, C2 => 
                           n5014, A => n1191, ZN => n1178);
   U3013 : AOI222_X1 port map( A1 => n5010, A2 => n4379, B1 => n5003, B2 => 
                           n4251, C1 => n4999, C2 => n4187, ZN => n1191);
   U3014 : OAI221_X1 port map( B1 => n3484, B2 => n5018, C1 => n3548, C2 => 
                           n5014, A => n1172, ZN => n1159);
   U3015 : AOI222_X1 port map( A1 => n5010, A2 => n4380, B1 => n5003, B2 => 
                           n4252, C1 => n4999, C2 => n4188, ZN => n1172);
   U3016 : OAI221_X1 port map( B1 => n3485, B2 => n5018, C1 => n3549, C2 => 
                           n5014, A => n1153, ZN => n1140);
   U3017 : AOI222_X1 port map( A1 => n5010, A2 => n4381, B1 => n5003, B2 => 
                           n4253, C1 => n4999, C2 => n4189, ZN => n1153);
   U3018 : OAI221_X1 port map( B1 => n3486, B2 => n5018, C1 => n3550, C2 => 
                           n5014, A => n1134, ZN => n1121);
   U3019 : AOI222_X1 port map( A1 => n5010, A2 => n4382, B1 => n5003, B2 => 
                           n4254, C1 => n4999, C2 => n4190, ZN => n1134);
   U3020 : OAI221_X1 port map( B1 => n3487, B2 => n5018, C1 => n3551, C2 => 
                           n5014, A => n1115, ZN => n1102);
   U3021 : AOI222_X1 port map( A1 => n5010, A2 => n4383, B1 => n5003, B2 => 
                           n4255, C1 => n4999, C2 => n4191, ZN => n1115);
   U3022 : OAI221_X1 port map( B1 => n3488, B2 => n5018, C1 => n3552, C2 => 
                           n5014, A => n1096, ZN => n1083);
   U3023 : AOI222_X1 port map( A1 => n5010, A2 => n4384, B1 => n5003, B2 => 
                           n4256, C1 => n4999, C2 => n4192, ZN => n1096);
   U3024 : OAI221_X1 port map( B1 => n3489, B2 => n5018, C1 => n3553, C2 => 
                           n5014, A => n1077, ZN => n1064);
   U3025 : AOI222_X1 port map( A1 => n5010, A2 => n4385, B1 => n5003, B2 => 
                           n4257, C1 => n4999, C2 => n4193, ZN => n1077);
   U3026 : OAI221_X1 port map( B1 => n3490, B2 => n5018, C1 => n3554, C2 => 
                           n5014, A => n1046, ZN => n1027);
   U3027 : AOI222_X1 port map( A1 => n5010, A2 => n4386, B1 => n5003, B2 => 
                           n4258, C1 => n4999, C2 => n4194, ZN => n1046);
   U3028 : OAI221_X1 port map( B1 => n3459, B2 => n5016, C1 => n3523, C2 => 
                           n5012, A => n2680, ZN => n2658);
   U3029 : AOI222_X1 port map( A1 => n5008, A2 => n4355, B1 => n5005, B2 => 
                           n4227, C1 => n5001, C2 => n4163, ZN => n2680);
   U3030 : OAI221_X1 port map( B1 => n3460, B2 => n5016, C1 => n3524, C2 => 
                           n5012, A => n2652, ZN => n2639);
   U3031 : AOI222_X1 port map( A1 => n5008, A2 => n4356, B1 => n5005, B2 => 
                           n4228, C1 => n5001, C2 => n4164, ZN => n2652);
   U3032 : OAI221_X1 port map( B1 => n3461, B2 => n5016, C1 => n3525, C2 => 
                           n5012, A => n2633, ZN => n2620);
   U3033 : AOI222_X1 port map( A1 => n5008, A2 => n4357, B1 => n5005, B2 => 
                           n4229, C1 => n5001, C2 => n4165, ZN => n2633);
   U3034 : OAI221_X1 port map( B1 => n3462, B2 => n5016, C1 => n3526, C2 => 
                           n5012, A => n2614, ZN => n2601);
   U3035 : AOI222_X1 port map( A1 => n5008, A2 => n4358, B1 => n5005, B2 => 
                           n4230, C1 => n5001, C2 => n4166, ZN => n2614);
   U3036 : OAI221_X1 port map( B1 => n3463, B2 => n5016, C1 => n3527, C2 => 
                           n5012, A => n2595, ZN => n2582);
   U3037 : AOI222_X1 port map( A1 => n5008, A2 => n4359, B1 => n5005, B2 => 
                           n4231, C1 => n5001, C2 => n4167, ZN => n2595);
   U3038 : OAI221_X1 port map( B1 => n3464, B2 => n5016, C1 => n3528, C2 => 
                           n5012, A => n2576, ZN => n2563);
   U3039 : AOI222_X1 port map( A1 => n5008, A2 => n4360, B1 => n5005, B2 => 
                           n4232, C1 => n5001, C2 => n4168, ZN => n2576);
   U3040 : OAI221_X1 port map( B1 => n3465, B2 => n5016, C1 => n3529, C2 => 
                           n5012, A => n2557, ZN => n2544);
   U3041 : AOI222_X1 port map( A1 => n5008, A2 => n4361, B1 => n5005, B2 => 
                           n4233, C1 => n5001, C2 => n4169, ZN => n2557);
   U3042 : OAI221_X1 port map( B1 => n3466, B2 => n5016, C1 => n3530, C2 => 
                           n5012, A => n2538, ZN => n2525);
   U3043 : AOI222_X1 port map( A1 => n5008, A2 => n4362, B1 => n5005, B2 => 
                           n4234, C1 => n5001, C2 => n4170, ZN => n2538);
   U3044 : OAI221_X1 port map( B1 => n3467, B2 => n5016, C1 => n3531, C2 => 
                           n5012, A => n2519, ZN => n2506);
   U3045 : AOI222_X1 port map( A1 => n5008, A2 => n4363, B1 => n5004, B2 => 
                           n4235, C1 => n5000, C2 => n4171, ZN => n2519);
   U3046 : OAI221_X1 port map( B1 => n3468, B2 => n5016, C1 => n3532, C2 => 
                           n5012, A => n2500, ZN => n2487);
   U3047 : AOI222_X1 port map( A1 => n5008, A2 => n4364, B1 => n5004, B2 => 
                           n4236, C1 => n5000, C2 => n4172, ZN => n2500);
   U3048 : OAI221_X1 port map( B1 => n3469, B2 => n5016, C1 => n3533, C2 => 
                           n5012, A => n2481, ZN => n2468);
   U3049 : AOI222_X1 port map( A1 => n5008, A2 => n4365, B1 => n5004, B2 => 
                           n4237, C1 => n5000, C2 => n4173, ZN => n2481);
   U3050 : OAI221_X1 port map( B1 => n3470, B2 => n5016, C1 => n3534, C2 => 
                           n5012, A => n2462, ZN => n2449);
   U3051 : AOI222_X1 port map( A1 => n5008, A2 => n4366, B1 => n5004, B2 => 
                           n4238, C1 => n5000, C2 => n4174, ZN => n2462);
   U3052 : OAI221_X1 port map( B1 => n3471, B2 => n5017, C1 => n3535, C2 => 
                           n5013, A => n2443, ZN => n2430);
   U3053 : AOI222_X1 port map( A1 => n5009, A2 => n4367, B1 => n5004, B2 => 
                           n4239, C1 => n5000, C2 => n4175, ZN => n2443);
   U3054 : OAI221_X1 port map( B1 => n3472, B2 => n5017, C1 => n3536, C2 => 
                           n5013, A => n2424, ZN => n2411);
   U3055 : AOI222_X1 port map( A1 => n5009, A2 => n4368, B1 => n5004, B2 => 
                           n4240, C1 => n5000, C2 => n4176, ZN => n2424);
   U3056 : OAI221_X1 port map( B1 => n3473, B2 => n5017, C1 => n3537, C2 => 
                           n5013, A => n2405, ZN => n2392);
   U3057 : AOI222_X1 port map( A1 => n5009, A2 => n4369, B1 => n5004, B2 => 
                           n4241, C1 => n5000, C2 => n4177, ZN => n2405);
   U3058 : OAI221_X1 port map( B1 => n3474, B2 => n5017, C1 => n3538, C2 => 
                           n5013, A => n2386, ZN => n2373);
   U3059 : AOI222_X1 port map( A1 => n5009, A2 => n4370, B1 => n5004, B2 => 
                           n4242, C1 => n5000, C2 => n4178, ZN => n2386);
   U3060 : OAI221_X1 port map( B1 => n3475, B2 => n5017, C1 => n3539, C2 => 
                           n5013, A => n2367, ZN => n2354);
   U3061 : AOI222_X1 port map( A1 => n5009, A2 => n4371, B1 => n5004, B2 => 
                           n4243, C1 => n5000, C2 => n4179, ZN => n2367);
   U3062 : OAI221_X1 port map( B1 => n3476, B2 => n5017, C1 => n3540, C2 => 
                           n5013, A => n2348, ZN => n2335);
   U3063 : AOI222_X1 port map( A1 => n5009, A2 => n4372, B1 => n5004, B2 => 
                           n4244, C1 => n5000, C2 => n4180, ZN => n2348);
   U3064 : OAI221_X1 port map( B1 => n3477, B2 => n5017, C1 => n3541, C2 => 
                           n5013, A => n2329, ZN => n1292);
   U3065 : AOI222_X1 port map( A1 => n5009, A2 => n4373, B1 => n5004, B2 => 
                           n4245, C1 => n5000, C2 => n4181, ZN => n2329);
   U3066 : OAI221_X1 port map( B1 => n3478, B2 => n5017, C1 => n3542, C2 => 
                           n5013, A => n1286, ZN => n1273);
   U3067 : AOI222_X1 port map( A1 => n5009, A2 => n4374, B1 => n5004, B2 => 
                           n4246, C1 => n5000, C2 => n4182, ZN => n1286);
   U3068 : OAI221_X1 port map( B1 => n3479, B2 => n5017, C1 => n3543, C2 => 
                           n5013, A => n1267, ZN => n1254);
   U3069 : AOI222_X1 port map( A1 => n5009, A2 => n4375, B1 => n5003, B2 => 
                           n4247, C1 => n4999, C2 => n4183, ZN => n1267);
   U3070 : OAI221_X1 port map( B1 => n3480, B2 => n5017, C1 => n3544, C2 => 
                           n5013, A => n1248, ZN => n1235);
   U3071 : AOI222_X1 port map( A1 => n5009, A2 => n4376, B1 => n5003, B2 => 
                           n4248, C1 => n4999, C2 => n4184, ZN => n1248);
   U3072 : OAI221_X1 port map( B1 => n3481, B2 => n5017, C1 => n3545, C2 => 
                           n5013, A => n1229, ZN => n1216);
   U3073 : AOI222_X1 port map( A1 => n5009, A2 => n4377, B1 => n5003, B2 => 
                           n4249, C1 => n4999, C2 => n4185, ZN => n1229);
   U3074 : OAI221_X1 port map( B1 => n3482, B2 => n5017, C1 => n3546, C2 => 
                           n5013, A => n1210, ZN => n1197);
   U3075 : AOI222_X1 port map( A1 => n5009, A2 => n4378, B1 => n5003, B2 => 
                           n4250, C1 => n4999, C2 => n4186, ZN => n1210);
   U3076 : OAI221_X1 port map( B1 => n3483, B2 => n5098, C1 => n3547, C2 => 
                           n5094, A => n553, ZN => n540);
   U3077 : AOI222_X1 port map( A1 => n5090, A2 => n4379, B1 => n5083, B2 => 
                           n4251, C1 => n5079, C2 => n4187, ZN => n553);
   U3078 : OAI221_X1 port map( B1 => n3484, B2 => n5098, C1 => n3548, C2 => 
                           n5094, A => n534, ZN => n521);
   U3079 : AOI222_X1 port map( A1 => n5090, A2 => n4380, B1 => n5083, B2 => 
                           n4252, C1 => n5079, C2 => n4188, ZN => n534);
   U3080 : OAI221_X1 port map( B1 => n3485, B2 => n5098, C1 => n3549, C2 => 
                           n5094, A => n515, ZN => n502);
   U3081 : AOI222_X1 port map( A1 => n5090, A2 => n4381, B1 => n5083, B2 => 
                           n4253, C1 => n5079, C2 => n4189, ZN => n515);
   U3082 : OAI221_X1 port map( B1 => n3486, B2 => n5098, C1 => n3550, C2 => 
                           n5094, A => n496, ZN => n483);
   U3083 : AOI222_X1 port map( A1 => n5090, A2 => n4382, B1 => n5083, B2 => 
                           n4254, C1 => n5079, C2 => n4190, ZN => n496);
   U3084 : OAI221_X1 port map( B1 => n3487, B2 => n5098, C1 => n3551, C2 => 
                           n5094, A => n477, ZN => n464);
   U3085 : AOI222_X1 port map( A1 => n5090, A2 => n4383, B1 => n5083, B2 => 
                           n4255, C1 => n5079, C2 => n4191, ZN => n477);
   U3086 : OAI221_X1 port map( B1 => n3488, B2 => n5098, C1 => n3552, C2 => 
                           n5094, A => n458, ZN => n445);
   U3087 : AOI222_X1 port map( A1 => n5090, A2 => n4384, B1 => n5083, B2 => 
                           n4256, C1 => n5079, C2 => n4192, ZN => n458);
   U3088 : OAI221_X1 port map( B1 => n3489, B2 => n5098, C1 => n3553, C2 => 
                           n5094, A => n439, ZN => n426);
   U3089 : AOI222_X1 port map( A1 => n5090, A2 => n4385, B1 => n5083, B2 => 
                           n4257, C1 => n5079, C2 => n4193, ZN => n439);
   U3090 : OAI221_X1 port map( B1 => n3490, B2 => n5098, C1 => n3554, C2 => 
                           n5094, A => n408, ZN => n389);
   U3091 : AOI222_X1 port map( A1 => n5090, A2 => n4386, B1 => n5083, B2 => 
                           n4258, C1 => n5079, C2 => n4194, ZN => n408);
   U3092 : OAI221_X1 port map( B1 => n3459, B2 => n5096, C1 => n3523, C2 => 
                           n5092, A => n1018, ZN => n996);
   U3093 : AOI222_X1 port map( A1 => n5088, A2 => n4355, B1 => n5085, B2 => 
                           n4227, C1 => n5081, C2 => n4163, ZN => n1018);
   U3094 : OAI221_X1 port map( B1 => n3460, B2 => n5096, C1 => n3524, C2 => 
                           n5092, A => n990, ZN => n977);
   U3095 : AOI222_X1 port map( A1 => n5088, A2 => n4356, B1 => n5085, B2 => 
                           n4228, C1 => n5081, C2 => n4164, ZN => n990);
   U3096 : OAI221_X1 port map( B1 => n3461, B2 => n5096, C1 => n3525, C2 => 
                           n5092, A => n971, ZN => n958);
   U3097 : AOI222_X1 port map( A1 => n5088, A2 => n4357, B1 => n5085, B2 => 
                           n4229, C1 => n5081, C2 => n4165, ZN => n971);
   U3098 : OAI221_X1 port map( B1 => n3462, B2 => n5096, C1 => n3526, C2 => 
                           n5092, A => n952, ZN => n939);
   U3099 : AOI222_X1 port map( A1 => n5088, A2 => n4358, B1 => n5085, B2 => 
                           n4230, C1 => n5081, C2 => n4166, ZN => n952);
   U3100 : OAI221_X1 port map( B1 => n3463, B2 => n5096, C1 => n3527, C2 => 
                           n5092, A => n933, ZN => n920);
   U3101 : AOI222_X1 port map( A1 => n5088, A2 => n4359, B1 => n5085, B2 => 
                           n4231, C1 => n5081, C2 => n4167, ZN => n933);
   U3102 : OAI221_X1 port map( B1 => n3464, B2 => n5096, C1 => n3528, C2 => 
                           n5092, A => n914, ZN => n901);
   U3103 : AOI222_X1 port map( A1 => n5088, A2 => n4360, B1 => n5085, B2 => 
                           n4232, C1 => n5081, C2 => n4168, ZN => n914);
   U3104 : OAI221_X1 port map( B1 => n3465, B2 => n5096, C1 => n3529, C2 => 
                           n5092, A => n895, ZN => n882);
   U3105 : AOI222_X1 port map( A1 => n5088, A2 => n4361, B1 => n5085, B2 => 
                           n4233, C1 => n5081, C2 => n4169, ZN => n895);
   U3106 : OAI221_X1 port map( B1 => n3466, B2 => n5096, C1 => n3530, C2 => 
                           n5092, A => n876, ZN => n863);
   U3107 : AOI222_X1 port map( A1 => n5088, A2 => n4362, B1 => n5085, B2 => 
                           n4234, C1 => n5081, C2 => n4170, ZN => n876);
   U3108 : OAI221_X1 port map( B1 => n3467, B2 => n5096, C1 => n3531, C2 => 
                           n5092, A => n857, ZN => n844);
   U3109 : AOI222_X1 port map( A1 => n5088, A2 => n4363, B1 => n5084, B2 => 
                           n4235, C1 => n5080, C2 => n4171, ZN => n857);
   U3110 : OAI221_X1 port map( B1 => n3468, B2 => n5096, C1 => n3532, C2 => 
                           n5092, A => n838, ZN => n825);
   U3111 : AOI222_X1 port map( A1 => n5088, A2 => n4364, B1 => n5084, B2 => 
                           n4236, C1 => n5080, C2 => n4172, ZN => n838);
   U3112 : OAI221_X1 port map( B1 => n3469, B2 => n5096, C1 => n3533, C2 => 
                           n5092, A => n819, ZN => n806);
   U3113 : AOI222_X1 port map( A1 => n5088, A2 => n4365, B1 => n5084, B2 => 
                           n4237, C1 => n5080, C2 => n4173, ZN => n819);
   U3114 : OAI221_X1 port map( B1 => n3470, B2 => n5096, C1 => n3534, C2 => 
                           n5092, A => n800, ZN => n787);
   U3115 : AOI222_X1 port map( A1 => n5088, A2 => n4366, B1 => n5084, B2 => 
                           n4238, C1 => n5080, C2 => n4174, ZN => n800);
   U3116 : OAI221_X1 port map( B1 => n3471, B2 => n5097, C1 => n3535, C2 => 
                           n5093, A => n781, ZN => n768);
   U3117 : AOI222_X1 port map( A1 => n5089, A2 => n4367, B1 => n5084, B2 => 
                           n4239, C1 => n5080, C2 => n4175, ZN => n781);
   U3118 : OAI221_X1 port map( B1 => n3472, B2 => n5097, C1 => n3536, C2 => 
                           n5093, A => n762, ZN => n749);
   U3119 : AOI222_X1 port map( A1 => n5089, A2 => n4368, B1 => n5084, B2 => 
                           n4240, C1 => n5080, C2 => n4176, ZN => n762);
   U3120 : OAI221_X1 port map( B1 => n3473, B2 => n5097, C1 => n3537, C2 => 
                           n5093, A => n743, ZN => n730);
   U3121 : AOI222_X1 port map( A1 => n5089, A2 => n4369, B1 => n5084, B2 => 
                           n4241, C1 => n5080, C2 => n4177, ZN => n743);
   U3122 : OAI221_X1 port map( B1 => n3474, B2 => n5097, C1 => n3538, C2 => 
                           n5093, A => n724, ZN => n711);
   U3123 : AOI222_X1 port map( A1 => n5089, A2 => n4370, B1 => n5084, B2 => 
                           n4242, C1 => n5080, C2 => n4178, ZN => n724);
   U3124 : OAI221_X1 port map( B1 => n3475, B2 => n5097, C1 => n3539, C2 => 
                           n5093, A => n705, ZN => n692);
   U3125 : AOI222_X1 port map( A1 => n5089, A2 => n4371, B1 => n5084, B2 => 
                           n4243, C1 => n5080, C2 => n4179, ZN => n705);
   U3126 : OAI221_X1 port map( B1 => n3476, B2 => n5097, C1 => n3540, C2 => 
                           n5093, A => n686, ZN => n673);
   U3127 : AOI222_X1 port map( A1 => n5089, A2 => n4372, B1 => n5084, B2 => 
                           n4244, C1 => n5080, C2 => n4180, ZN => n686);
   U3128 : OAI221_X1 port map( B1 => n3477, B2 => n5097, C1 => n3541, C2 => 
                           n5093, A => n667, ZN => n654);
   U3129 : AOI222_X1 port map( A1 => n5089, A2 => n4373, B1 => n5084, B2 => 
                           n4245, C1 => n5080, C2 => n4181, ZN => n667);
   U3130 : OAI221_X1 port map( B1 => n3478, B2 => n5097, C1 => n3542, C2 => 
                           n5093, A => n648, ZN => n635);
   U3131 : AOI222_X1 port map( A1 => n5089, A2 => n4374, B1 => n5084, B2 => 
                           n4246, C1 => n5080, C2 => n4182, ZN => n648);
   U3132 : OAI221_X1 port map( B1 => n3479, B2 => n5097, C1 => n3543, C2 => 
                           n5093, A => n629, ZN => n616);
   U3133 : AOI222_X1 port map( A1 => n5089, A2 => n4375, B1 => n5083, B2 => 
                           n4247, C1 => n5079, C2 => n4183, ZN => n629);
   U3134 : OAI221_X1 port map( B1 => n3480, B2 => n5097, C1 => n3544, C2 => 
                           n5093, A => n610, ZN => n597);
   U3135 : AOI222_X1 port map( A1 => n5089, A2 => n4376, B1 => n5083, B2 => 
                           n4248, C1 => n5079, C2 => n4184, ZN => n610);
   U3136 : OAI221_X1 port map( B1 => n3481, B2 => n5097, C1 => n3545, C2 => 
                           n5093, A => n591, ZN => n578);
   U3137 : AOI222_X1 port map( A1 => n5089, A2 => n4377, B1 => n5083, B2 => 
                           n4249, C1 => n5079, C2 => n4185, ZN => n591);
   U3138 : OAI221_X1 port map( B1 => n3482, B2 => n5097, C1 => n3546, C2 => 
                           n5093, A => n572, ZN => n559);
   U3139 : AOI222_X1 port map( A1 => n5089, A2 => n4378, B1 => n5083, B2 => 
                           n4250, C1 => n5079, C2 => n4186, ZN => n572);
   U3140 : INV_X1 port map( A => ADD_RD1(3), ZN => n5151);
   U3141 : INV_X1 port map( A => ADD_RD2(3), ZN => n5138);
   U3142 : NOR2_X1 port map( A1 => n5152, A2 => ADD_RD1(3), ZN => n1001);
   U3143 : INV_X1 port map( A => ADD_RD1(4), ZN => n5152);
   U3144 : NOR2_X1 port map( A1 => n5139, A2 => ADD_RD2(3), ZN => n2663);
   U3145 : INV_X1 port map( A => ADD_RD2(4), ZN => n5139);
   U3146 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => n5152, ZN => n392);
   U3147 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => n5139, ZN => n1030);
   U3148 : NAND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => n386);
   U3149 : NAND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => n1024);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity SIGN_EXT_bits16 is

   port( inputt : in std_logic_vector (15 downto 0);  outputt : out 
         std_logic_vector (31 downto 0));

end SIGN_EXT_bits16;

architecture SYN_BEHAVIORAL of SIGN_EXT_bits16 is

begin
   outputt <= ( inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), 
      inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), 
      inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), 
      inputt(14), inputt(13), inputt(12), inputt(11), inputt(10), inputt(9), 
      inputt(8), inputt(7), inputt(6), inputt(5), inputt(4), inputt(3), 
      inputt(2), inputt(1), inputt(0) );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_8 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_8;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_8 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_225
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_226
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_227
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_228
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_229
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_230
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_231
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_232
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_233
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_234
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_235
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_236
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_237
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_238
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_239
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_240
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_241
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_242
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_243
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_244
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_245
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_246
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_247
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_248
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_249
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_250
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_251
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_252
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_253
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_254
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_255
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_256
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12 : std_logic;

begin
   
   FF_0 : FD_256 port map( D => data_in(0), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_255 port map( D => data_in(1), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_254 port map( D => data_in(2), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_253 port map( D => data_in(3), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_252 port map( D => data_in(4), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_251 port map( D => data_in(5), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_250 port map( D => data_in(6), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_249 port map( D => data_in(7), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_248 port map( D => data_in(8), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_247 port map( D => data_in(9), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_246 port map( D => data_in(10), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_245 port map( D => data_in(11), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_244 port map( D => data_in(12), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(12));
   FF_13 : FD_243 port map( D => data_in(13), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(13));
   FF_14 : FD_242 port map( D => data_in(14), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(14));
   FF_15 : FD_241 port map( D => data_in(15), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(15));
   FF_16 : FD_240 port map( D => data_in(16), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(16));
   FF_17 : FD_239 port map( D => data_in(17), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(17));
   FF_18 : FD_238 port map( D => data_in(18), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(18));
   FF_19 : FD_237 port map( D => data_in(19), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(19));
   FF_20 : FD_236 port map( D => data_in(20), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(20));
   FF_21 : FD_235 port map( D => data_in(21), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(21));
   FF_22 : FD_234 port map( D => data_in(22), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(22));
   FF_23 : FD_233 port map( D => data_in(23), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(23));
   FF_24 : FD_232 port map( D => data_in(24), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(24));
   FF_25 : FD_231 port map( D => data_in(25), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(25));
   FF_26 : FD_230 port map( D => data_in(26), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(26));
   FF_27 : FD_229 port map( D => data_in(27), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(27));
   FF_28 : FD_228 port map( D => data_in(28), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(28));
   FF_29 : FD_227 port map( D => data_in(29), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(29));
   FF_30 : FD_226 port map( D => data_in(30), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(30));
   FF_31 : FD_225 port map( D => data_in(31), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => n12, Z => n9);
   U3 : BUF_X1 port map( A => n12, Z => n10);
   U4 : BUF_X1 port map( A => n12, Z => n11);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_0 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_0;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_321
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_322
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_323
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_324
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_325
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_326
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_327
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_328
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_329
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_330
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_331
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_332
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_333
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_334
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_335
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_336
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_337
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_338
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_339
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_340
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_341
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_342
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_343
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_344
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_345
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_346
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_347
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_348
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_349
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_350
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_351
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_352
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12 : std_logic;

begin
   
   FF_0 : FD_352 port map( D => data_in(0), CK => CK, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_351 port map( D => data_in(1), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_350 port map( D => data_in(2), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_349 port map( D => data_in(3), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_348 port map( D => data_in(4), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_347 port map( D => data_in(5), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_346 port map( D => data_in(6), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_345 port map( D => data_in(7), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_344 port map( D => data_in(8), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_343 port map( D => data_in(9), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_342 port map( D => data_in(10), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_341 port map( D => data_in(11), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_340 port map( D => data_in(12), CK => CK, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_339 port map( D => data_in(13), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(13));
   FF_14 : FD_338 port map( D => data_in(14), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(14));
   FF_15 : FD_337 port map( D => data_in(15), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(15));
   FF_16 : FD_336 port map( D => data_in(16), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(16));
   FF_17 : FD_335 port map( D => data_in(17), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(17));
   FF_18 : FD_334 port map( D => data_in(18), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(18));
   FF_19 : FD_333 port map( D => data_in(19), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(19));
   FF_20 : FD_332 port map( D => data_in(20), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(20));
   FF_21 : FD_331 port map( D => data_in(21), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(21));
   FF_22 : FD_330 port map( D => data_in(22), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(22));
   FF_23 : FD_329 port map( D => data_in(23), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(23));
   FF_24 : FD_328 port map( D => data_in(24), CK => CK, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(24));
   FF_25 : FD_327 port map( D => data_in(25), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(25));
   FF_26 : FD_326 port map( D => data_in(26), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(26));
   FF_27 : FD_325 port map( D => data_in(27), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(27));
   FF_28 : FD_324 port map( D => data_in(28), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(28));
   FF_29 : FD_323 port map( D => data_in(29), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(29));
   FF_30 : FD_322 port map( D => data_in(30), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(30));
   FF_31 : FD_321 port map( D => data_in(31), CK => CK, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => n12, Z => n9);
   U3 : BUF_X1 port map( A => n12, Z => n10);
   U4 : BUF_X1 port map( A => n12, Z => n11);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end RCA_NBITS32;

architecture SYN_BEHAVIORAL of RCA_NBITS32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n54, n55, n56, n57, n59, n60, n63, n64, n65, n70, n71, n73, n74, n75,
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n109, n110, n111, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n180, n179, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n258, n259, n260, n261, n262, n263, n264, n265, 
      n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
      n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
      n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300 : 
      std_logic;

begin
   
   U126 : XOR2_X1 port map( A => n54, B => n55, Z => S(9));
   U127 : XOR2_X1 port map( A => Ci, B => B(9), Z => n55);
   U128 : XOR2_X1 port map( A => n274, B => A(9), Z => n54);
   U129 : XOR2_X1 port map( A => n56, B => n57, Z => S(8));
   U130 : XOR2_X1 port map( A => A(8), B => n204, Z => n57);
   U131 : XOR2_X1 port map( A => Ci, B => B(8), Z => n56);
   U132 : XOR2_X1 port map( A => n59, B => n60, Z => S(7));
   U133 : XOR2_X1 port map( A => Ci, B => B(7), Z => n60);
   U137 : XOR2_X1 port map( A => n64, B => n65, Z => S(5));
   U138 : XOR2_X1 port map( A => Ci, B => B(5), Z => n65);
   U139 : XOR2_X1 port map( A => n221, B => A(5), Z => n64);
   U146 : XOR2_X1 port map( A => Ci, B => B(31), Z => n71);
   U147 : XOR2_X1 port map( A => n74, B => n75, Z => S(30));
   U149 : XOR2_X1 port map( A => Ci, B => B(30), Z => n74);
   U150 : XOR2_X1 port map( A => n76, B => n77, Z => S(2));
   U151 : XOR2_X1 port map( A => Ci, B => B(2), Z => n77);
   U152 : XOR2_X1 port map( A => A(2), B => n234, Z => n76);
   U153 : XOR2_X1 port map( A => n78, B => n79, Z => S(29));
   U154 : XOR2_X1 port map( A => Ci, B => B(29), Z => n79);
   U155 : XOR2_X1 port map( A => n206, B => A(29), Z => n78);
   U156 : XOR2_X1 port map( A => n81, B => n82, Z => S(28));
   U157 : XOR2_X1 port map( A => Ci, B => B(28), Z => n82);
   U158 : XOR2_X1 port map( A => n211, B => A(28), Z => n81);
   U159 : XOR2_X1 port map( A => n84, B => n85, Z => S(27));
   U160 : XOR2_X1 port map( A => Ci, B => B(27), Z => n85);
   U161 : XOR2_X1 port map( A => n209, B => A(27), Z => n84);
   U162 : XOR2_X1 port map( A => n87, B => n88, Z => S(26));
   U163 : XOR2_X1 port map( A => Ci, B => B(26), Z => n88);
   U164 : XOR2_X1 port map( A => n208, B => A(26), Z => n87);
   U165 : XOR2_X1 port map( A => n90, B => n91, Z => S(25));
   U166 : XOR2_X1 port map( A => Ci, B => B(25), Z => n91);
   U167 : XOR2_X1 port map( A => n207, B => A(25), Z => n90);
   U168 : XOR2_X1 port map( A => n93, B => n94, Z => S(24));
   U169 : XOR2_X1 port map( A => Ci, B => B(24), Z => n94);
   U170 : XOR2_X1 port map( A => n243, B => A(24), Z => n93);
   U171 : XOR2_X1 port map( A => n96, B => n97, Z => S(23));
   U172 : XOR2_X1 port map( A => Ci, B => B(23), Z => n97);
   U173 : XOR2_X1 port map( A => n242, B => A(23), Z => n96);
   U174 : XOR2_X1 port map( A => n99, B => n100, Z => S(22));
   U175 : XOR2_X1 port map( A => Ci, B => B(22), Z => n100);
   U176 : XOR2_X1 port map( A => n239, B => A(22), Z => n99);
   U177 : XOR2_X1 port map( A => n102, B => n103, Z => S(21));
   U178 : XOR2_X1 port map( A => Ci, B => B(21), Z => n103);
   U179 : XOR2_X1 port map( A => n267, B => A(21), Z => n102);
   U180 : XOR2_X1 port map( A => n104, B => n105, Z => S(20));
   U181 : XOR2_X1 port map( A => Ci, B => B(20), Z => n105);
   U182 : XOR2_X1 port map( A => n106, B => A(20), Z => n104);
   U185 : XOR2_X1 port map( A => n110, B => n111, Z => S(19));
   U186 : XOR2_X1 port map( A => n288, B => n226, Z => n111);
   U187 : XOR2_X1 port map( A => B(19), B => n300, Z => n110);
   U190 : XOR2_X1 port map( A => n115, B => n116, Z => S(17));
   U191 : XOR2_X1 port map( A => Ci, B => B(17), Z => n116);
   U192 : XOR2_X1 port map( A => n287, B => n270, Z => n115);
   U193 : XOR2_X1 port map( A => n117, B => n118, Z => S(16));
   U194 : XOR2_X1 port map( A => n233, B => A(16), Z => n118);
   U195 : XOR2_X1 port map( A => B(16), B => n300, Z => n117);
   U196 : XOR2_X1 port map( A => n120, B => n121, Z => S(15));
   U198 : XOR2_X1 port map( A => B(15), B => n300, Z => n120);
   U199 : XOR2_X1 port map( A => n123, B => n124, Z => S(14));
   U200 : XOR2_X1 port map( A => B(14), B => n300, Z => n123);
   U201 : XOR2_X1 port map( A => n126, B => n127, Z => S(13));
   U202 : XOR2_X1 port map( A => n222, B => A(13), Z => n127);
   U203 : XOR2_X1 port map( A => B(13), B => n300, Z => n126);
   U204 : XOR2_X1 port map( A => n129, B => n130, Z => S(12));
   U205 : XOR2_X1 port map( A => A(12), B => n216, Z => n130);
   U206 : XOR2_X1 port map( A => Ci, B => B(12), Z => n129);
   U207 : XOR2_X1 port map( A => n132, B => n133, Z => S(11));
   U208 : XOR2_X1 port map( A => Ci, B => B(11), Z => n133);
   U209 : XOR2_X1 port map( A => n235, B => A(11), Z => n132);
   U210 : XOR2_X1 port map( A => n134, B => n135, Z => S(10));
   U211 : XOR2_X1 port map( A => A(10), B => n237, Z => n135);
   U212 : XOR2_X1 port map( A => Ci, B => B(10), Z => n134);
   U213 : XOR2_X1 port map( A => n298, B => B(0), Z => n138);
   U2 : OAI21_X2 port map( B1 => n154, B2 => n288, A => n155, ZN => n106);
   U3 : NAND2_X1 port map( A1 => n179, A2 => n172, ZN => n220);
   U4 : NAND2_X1 port map( A1 => n227, A2 => A(6), ZN => n179);
   U5 : AOI21_X1 port map( B1 => n281, B2 => n173, A => n174, ZN => n181);
   U6 : CLKBUF_X1 port map( A => n174, Z => n182);
   U7 : CLKBUF_X1 port map( A => n168, Z => n183);
   U8 : BUF_X1 port map( A => n171, Z => n188);
   U9 : AOI21_X1 port map( B1 => n281, B2 => n173, A => n174, ZN => n227);
   U10 : AOI21_X1 port map( B1 => n185, B2 => A(5), A => B(5), ZN => n174);
   U11 : OAI21_X1 port map( B1 => n176, B2 => n184, A => n175, ZN => n185);
   U12 : INV_X1 port map( A => A(4), ZN => n184);
   U13 : INV_X1 port map( A => n185, ZN => n173);
   U14 : CLKBUF_X1 port map( A => n187, Z => n186);
   U15 : AND2_X1 port map( A1 => n181, A2 => A(6), ZN => n187);
   U16 : OR2_X1 port map( A1 => n187, A2 => n189, ZN => n192);
   U17 : NAND2_X1 port map( A1 => n172, A2 => n282, ZN => n189);
   U18 : NOR2_X1 port map( A1 => n188, A2 => n191, ZN => n190);
   U19 : NOR2_X1 port map( A1 => n191, A2 => n171, ZN => n238);
   U20 : NAND2_X1 port map( A1 => n192, A2 => A(8), ZN => n191);
   U21 : AND2_X1 port map( A1 => n282, A2 => n170, ZN => n193);
   U22 : CLKBUF_X1 port map( A => n141, Z => n218);
   U23 : CLKBUF_X1 port map( A => n165, Z => n194);
   U24 : BUF_X1 port map( A => n232, Z => n202);
   U25 : NAND2_X1 port map( A1 => n180, A2 => n197, ZN => n195);
   U26 : AND2_X1 port map( A1 => n195, A2 => n196, ZN => n201);
   U27 : OR2_X1 port map( A1 => n280, A2 => A(2), ZN => n196);
   U28 : AND2_X1 port map( A1 => n202, A2 => n178, ZN => n197);
   U29 : NOR2_X1 port map( A1 => n198, A2 => n199, ZN => n219);
   U30 : NOR2_X1 port map( A1 => n200, A2 => n280, ZN => n198);
   U31 : NOR2_X1 port map( A1 => n280, A2 => A(2), ZN => n199);
   U32 : XNOR2_X1 port map( A => n218, B => A(30), ZN => n75);
   U33 : NAND2_X1 port map( A1 => n232, A2 => n180, ZN => n200);
   U34 : CLKBUF_X1 port map( A => n240, Z => n203);
   U35 : NOR2_X1 port map( A1 => n188, A2 => n193, ZN => n204);
   U36 : AOI21_X1 port map( B1 => n283, B2 => n167, A => n183, ZN => n205);
   U37 : CLKBUF_X1 port map( A => n80, Z => n206);
   U38 : OAI21_X1 port map( B1 => n260, B2 => n296, A => n144, ZN => n80);
   U39 : CLKBUF_X1 port map( A => n92, Z => n207);
   U40 : OAI21_X1 port map( B1 => n264, B2 => n292, A => n148, ZN => n92);
   U41 : CLKBUF_X1 port map( A => n89, Z => n208);
   U42 : OAI21_X1 port map( B1 => n263, B2 => n293, A => n147, ZN => n89);
   U43 : CLKBUF_X1 port map( A => n86, Z => n209);
   U44 : OAI21_X1 port map( B1 => n262, B2 => n294, A => n146, ZN => n86);
   U45 : CLKBUF_X1 port map( A => n114, Z => n210);
   U46 : OAI21_X1 port map( B1 => n270, B2 => n287, A => n157, ZN => n114);
   U47 : CLKBUF_X1 port map( A => n83, Z => n211);
   U48 : OAI21_X1 port map( B1 => n261, B2 => n295, A => n145, ZN => n83);
   U49 : AOI21_X1 port map( B1 => n297, B2 => n218, A => n142, ZN => n212);
   U50 : AOI21_X1 port map( B1 => n297, B2 => n218, A => n142, ZN => n73);
   U51 : AOI21_X1 port map( B1 => n285, B2 => n222, A => n162, ZN => n213);
   U52 : AOI21_X1 port map( B1 => n285, B2 => n222, A => n162, ZN => n125);
   U53 : INV_X1 port map( A => n270, ZN => n214);
   U54 : CLKBUF_X1 port map( A => n173, Z => n255);
   U55 : AOI21_X1 port map( B1 => n284, B2 => n164, A => n165, ZN => n215);
   U56 : AOI21_X1 port map( B1 => n284, B2 => n164, A => n194, ZN => n216);
   U57 : AOI21_X1 port map( B1 => n284, B2 => n164, A => n165, ZN => n131);
   U58 : OR2_X1 port map( A1 => n163, A2 => n223, ZN => n222);
   U59 : OR2_X1 port map( A1 => n238, A2 => n275, ZN => n217);
   U60 : INV_X1 port map( A => n255, ZN => n221);
   U61 : NOR2_X1 port map( A1 => n163, A2 => n223, ZN => n225);
   U62 : NOR2_X1 port map( A1 => n215, A2 => A(12), ZN => n223);
   U63 : AND2_X1 port map( A1 => n210, A2 => A(18), ZN => n224);
   U64 : OR2_X1 port map( A1 => n224, A2 => n269, ZN => n226);
   U65 : AOI21_X1 port map( B1 => n281, B2 => n255, A => n182, ZN => n63);
   U66 : CLKBUF_X1 port map( A => A(1), Z => n228);
   U67 : NAND2_X1 port map( A1 => n180, A2 => n202, ZN => n229);
   U68 : CLKBUF_X1 port map( A => A(0), Z => n230);
   U69 : AND2_X1 port map( A1 => n114, A2 => A(18), ZN => n231);
   U70 : NOR2_X1 port map( A1 => n231, A2 => n269, ZN => n154);
   U71 : NAND2_X1 port map( A1 => n109, A2 => A(1), ZN => n232);
   U72 : BUF_X1 port map( A => n119, Z => n233);
   U73 : CLKBUF_X1 port map( A => n229, Z => n234);
   U74 : OR2_X1 port map( A1 => n240, A2 => n273, ZN => n235);
   U75 : AND2_X1 port map( A1 => n229, A2 => A(2), ZN => n236);
   U76 : NOR2_X1 port map( A1 => n236, A2 => n280, ZN => n70);
   U77 : NOR2_X1 port map( A1 => n186, A2 => n277, ZN => n170);
   U78 : CLKBUF_X1 port map( A => n205, Z => n237);
   U79 : NOR2_X1 port map( A1 => n190, A2 => n275, ZN => n167);
   U80 : AOI21_X1 port map( B1 => n283, B2 => n167, A => n168, ZN => n136);
   U81 : CLKBUF_X1 port map( A => n101, Z => n239);
   U82 : AND2_X1 port map( A1 => n136, A2 => A(10), ZN => n240);
   U83 : NOR2_X1 port map( A1 => n203, A2 => n273, ZN => n164);
   U84 : AND2_X1 port map( A1 => B(0), A2 => n230, ZN => n241);
   U85 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n109);
   U86 : CLKBUF_X1 port map( A => n98, Z => n242);
   U87 : CLKBUF_X1 port map( A => n95, Z => n243);
   U88 : XOR2_X1 port map( A => n276, B => A(7), Z => n59);
   U89 : INV_X1 port map( A => n139, ZN => Co);
   U90 : INV_X1 port map( A => A(15), ZN => n256);
   U91 : INV_X1 port map( A => A(21), ZN => n289);
   U92 : INV_X1 port map( A => n169, ZN => n275);
   U93 : INV_X1 port map( A => n166, ZN => n273);
   U94 : INV_X1 port map( A => A(16), ZN => n286);
   U95 : OAI21_X1 port map( B1 => n266, B2 => n290, A => n150, ZN => n98);
   U96 : INV_X1 port map( A => A(22), ZN => n290);
   U97 : INV_X1 port map( A => A(27), ZN => n295);
   U98 : INV_X1 port map( A => A(11), ZN => n284);
   U99 : INV_X1 port map( A => A(13), ZN => n285);
   U100 : INV_X1 port map( A => A(7), ZN => n282);
   U101 : INV_X1 port map( A => A(9), ZN => n283);
   U102 : INV_X1 port map( A => A(5), ZN => n281);
   U103 : XNOR2_X1 port map( A => n244, B => n71, ZN => S(31));
   U104 : XNOR2_X1 port map( A => n73, B => A(31), ZN => n244);
   U105 : INV_X1 port map( A => A(30), ZN => n297);
   U106 : OAI21_X1 port map( B1 => n265, B2 => n291, A => n149, ZN => n95);
   U107 : OAI21_X1 port map( B1 => A(23), B2 => n242, A => B(23), ZN => n149);
   U108 : INV_X1 port map( A => A(23), ZN => n291);
   U109 : INV_X1 port map( A => A(24), ZN => n292);
   U110 : INV_X1 port map( A => A(25), ZN => n293);
   U111 : INV_X1 port map( A => A(26), ZN => n294);
   U112 : OAI21_X1 port map( B1 => A(19), B2 => n226, A => B(19), ZN => n155);
   U113 : OAI21_X1 port map( B1 => A(28), B2 => n211, A => B(28), ZN => n144);
   U114 : INV_X1 port map( A => A(28), ZN => n296);
   U115 : XOR2_X1 port map( A => n245, B => n246, Z => S(18));
   U116 : XNOR2_X1 port map( A => B(18), B => n300, ZN => n245);
   U117 : XOR2_X1 port map( A => A(18), B => n210, Z => n246);
   U118 : XNOR2_X1 port map( A => n272, B => A(15), ZN => n121);
   U119 : INV_X1 port map( A => A(17), ZN => n287);
   U120 : INV_X1 port map( A => A(19), ZN => n288);
   U121 : XOR2_X1 port map( A => n247, B => n248, Z => S(6));
   U122 : XNOR2_X1 port map( A => B(6), B => n300, ZN => n247);
   U123 : XOR2_X1 port map( A => n63, B => A(6), Z => n248);
   U124 : XOR2_X1 port map( A => n249, B => n250, Z => S(4));
   U125 : XNOR2_X1 port map( A => B(4), B => n300, ZN => n249);
   U134 : XOR2_X1 port map( A => n278, B => A(4), Z => n250);
   U135 : XOR2_X1 port map( A => n251, B => n252, Z => S(3));
   U136 : XOR2_X1 port map( A => n70, B => A(3), Z => n251);
   U140 : XNOR2_X1 port map( A => Ci, B => B(3), ZN => n252);
   U141 : OAI22_X1 port map( A1 => n137, A2 => n300, B1 => Ci, B2 => n138, ZN 
                           => S(0));
   U142 : XOR2_X1 port map( A => n253, B => n254, Z => S(1));
   U143 : XNOR2_X1 port map( A => B(1), B => n300, ZN => n253);
   U144 : XOR2_X1 port map( A => n241, B => n228, Z => n254);
   U145 : INV_X1 port map( A => Ci, ZN => n300);
   U148 : INV_X1 port map( A => B(0), ZN => n299);
   U183 : OAI21_X1 port map( B1 => A(27), B2 => n209, A => B(27), ZN => n145);
   U184 : INV_X1 port map( A => n176, ZN => n278);
   U188 : OAI21_X1 port map( B1 => A(17), B2 => n214, A => B(17), ZN => n157);
   U189 : OAI21_X1 port map( B1 => n271, B2 => A(16), A => B(16), ZN => n159);
   U197 : AOI21_X1 port map( B1 => n219, B2 => A(3), A => B(3), ZN => n177);
   U214 : AOI21_X1 port map( B1 => n80, B2 => A(29), A => B(29), ZN => n143);
   U215 : INV_X1 port map( A => n83, ZN => n260);
   U216 : INV_X1 port map( A => n98, ZN => n265);
   U217 : NOR2_X1 port map( A1 => n122, A2 => n256, ZN => n160);
   U218 : OAI22_X1 port map( A1 => A(15), A2 => n272, B1 => n160, B2 => B(15), 
                           ZN => n119);
   U219 : INV_X1 port map( A => n230, ZN => n298);
   U220 : OAI21_X1 port map( B1 => A(2), B2 => n234, A => B(2), ZN => n178);
   U221 : OAI21_X1 port map( B1 => n278, B2 => A(4), A => B(4), ZN => n175);
   U222 : AOI21_X1 port map( B1 => n235, B2 => A(11), A => B(11), ZN => n165);
   U223 : OAI21_X1 port map( B1 => A(29), B2 => n206, A => n259, ZN => n141);
   U224 : INV_X1 port map( A => n178, ZN => n280);
   U225 : INV_X1 port map( A => n158, ZN => n270);
   U226 : INV_X1 port map( A => n122, ZN => n272);
   U227 : OAI21_X1 port map( B1 => A(3), B2 => n201, A => n279, ZN => n176);
   U228 : INV_X1 port map( A => n177, ZN => n279);
   U229 : AOI21_X1 port map( B1 => n258, B2 => A(30), A => B(30), ZN => n142);
   U230 : AOI21_X1 port map( B1 => n217, B2 => A(9), A => B(9), ZN => n168);
   U231 : INV_X1 port map( A => n167, ZN => n274);
   U232 : AOI21_X1 port map( B1 => n225, B2 => A(13), A => B(13), ZN => n162);
   U233 : AOI21_X1 port map( B1 => n220, B2 => A(7), A => B(7), ZN => n171);
   U234 : INV_X1 port map( A => n153, ZN => n268);
   U235 : OAI21_X1 port map( B1 => A(21), B2 => n267, A => B(21), ZN => n152);
   U236 : OAI21_X1 port map( B1 => A(24), B2 => n243, A => B(24), ZN => n148);
   U237 : INV_X1 port map( A => n143, ZN => n259);
   U238 : INV_X1 port map( A => n95, ZN => n264);
   U239 : OAI21_X1 port map( B1 => n151, B2 => n289, A => n152, ZN => n101);
   U240 : INV_X1 port map( A => n151, ZN => n267);
   U241 : AOI21_X1 port map( B1 => n106, B2 => A(20), A => n268, ZN => n151);
   U242 : OAI21_X1 port map( B1 => A(20), B2 => n106, A => B(20), ZN => n153);
   U243 : INV_X1 port map( A => n86, ZN => n261);
   U244 : INV_X1 port map( A => n170, ZN => n276);
   U245 : INV_X1 port map( A => n172, ZN => n277);
   U246 : INV_X1 port map( A => n156, ZN => n269);
   U247 : OR2_X1 port map( A1 => n212, A2 => A(31), ZN => n140);
   U248 : AOI21_X1 port map( B1 => n298, B2 => n299, A => n241, ZN => n137);
   U249 : OAI21_X1 port map( B1 => A(22), B2 => n239, A => B(22), ZN => n150);
   U250 : OAI21_X1 port map( B1 => A(26), B2 => n208, A => B(26), ZN => n146);
   U251 : AOI22_X1 port map( A1 => A(31), A2 => n212, B1 => n140, B2 => B(31), 
                           ZN => n139);
   U252 : XNOR2_X1 port map( A => n213, B => A(14), ZN => n124);
   U253 : INV_X1 port map( A => n141, ZN => n258);
   U254 : INV_X1 port map( A => n89, ZN => n262);
   U255 : OAI21_X1 port map( B1 => A(25), B2 => n207, A => B(25), ZN => n147);
   U256 : INV_X1 port map( A => n92, ZN => n263);
   U257 : INV_X1 port map( A => n101, ZN => n266);
   U258 : OAI21_X1 port map( B1 => A(18), B2 => n210, A => B(18), ZN => n156);
   U259 : OAI21_X1 port map( B1 => n119, B2 => n286, A => n159, ZN => n158);
   U260 : INV_X1 port map( A => n233, ZN => n271);
   U261 : OAI22_X1 port map( A1 => A(14), A2 => n213, B1 => n161, B2 => B(14), 
                           ZN => n122);
   U262 : AND2_X1 port map( A1 => n125, A2 => A(14), ZN => n161);
   U263 : AOI21_X1 port map( B1 => n131, B2 => A(12), A => B(12), ZN => n163);
   U264 : OAI21_X1 port map( B1 => n237, B2 => A(10), A => B(10), ZN => n166);
   U265 : OAI21_X1 port map( B1 => n204, B2 => A(8), A => B(8), ZN => n169);
   U266 : OAI21_X1 port map( B1 => n63, B2 => A(6), A => B(6), ZN => n172);
   U267 : OAI21_X1 port map( B1 => n241, B2 => n228, A => B(1), ZN => n180);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity writeBack_nbits32 is

   port( LMD_OUT, ALUREG_OUTPUT : in std_logic_vector (31 downto 0);  
         WB_MUX_SEL : in std_logic;  DATAIN_RF : out std_logic_vector (31 
         downto 0));

end writeBack_nbits32;

architecture SYN_STRUCTURAL of writeBack_nbits32 is

   component MUX21_GENERIC_bits32_1
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;

begin
   
   MUXWB : MUX21_GENERIC_bits32_1 port map( A(31) => ALUREG_OUTPUT(31), A(30) 
                           => ALUREG_OUTPUT(30), A(29) => ALUREG_OUTPUT(29), 
                           A(28) => ALUREG_OUTPUT(28), A(27) => 
                           ALUREG_OUTPUT(27), A(26) => ALUREG_OUTPUT(26), A(25)
                           => ALUREG_OUTPUT(25), A(24) => ALUREG_OUTPUT(24), 
                           A(23) => ALUREG_OUTPUT(23), A(22) => 
                           ALUREG_OUTPUT(22), A(21) => ALUREG_OUTPUT(21), A(20)
                           => ALUREG_OUTPUT(20), A(19) => ALUREG_OUTPUT(19), 
                           A(18) => ALUREG_OUTPUT(18), A(17) => 
                           ALUREG_OUTPUT(17), A(16) => ALUREG_OUTPUT(16), A(15)
                           => ALUREG_OUTPUT(15), A(14) => ALUREG_OUTPUT(14), 
                           A(13) => ALUREG_OUTPUT(13), A(12) => 
                           ALUREG_OUTPUT(12), A(11) => ALUREG_OUTPUT(11), A(10)
                           => ALUREG_OUTPUT(10), A(9) => ALUREG_OUTPUT(9), A(8)
                           => ALUREG_OUTPUT(8), A(7) => ALUREG_OUTPUT(7), A(6) 
                           => ALUREG_OUTPUT(6), A(5) => ALUREG_OUTPUT(5), A(4) 
                           => ALUREG_OUTPUT(4), A(3) => ALUREG_OUTPUT(3), A(2) 
                           => ALUREG_OUTPUT(2), A(1) => ALUREG_OUTPUT(1), A(0) 
                           => ALUREG_OUTPUT(0), B(31) => LMD_OUT(31), B(30) => 
                           LMD_OUT(30), B(29) => LMD_OUT(29), B(28) => 
                           LMD_OUT(28), B(27) => LMD_OUT(27), B(26) => 
                           LMD_OUT(26), B(25) => LMD_OUT(25), B(24) => 
                           LMD_OUT(24), B(23) => LMD_OUT(23), B(22) => 
                           LMD_OUT(22), B(21) => LMD_OUT(21), B(20) => 
                           LMD_OUT(20), B(19) => LMD_OUT(19), B(18) => 
                           LMD_OUT(18), B(17) => LMD_OUT(17), B(16) => 
                           LMD_OUT(16), B(15) => LMD_OUT(15), B(14) => 
                           LMD_OUT(14), B(13) => LMD_OUT(13), B(12) => 
                           LMD_OUT(12), B(11) => LMD_OUT(11), B(10) => 
                           LMD_OUT(10), B(9) => LMD_OUT(9), B(8) => LMD_OUT(8),
                           B(7) => LMD_OUT(7), B(6) => LMD_OUT(6), B(5) => 
                           LMD_OUT(5), B(4) => LMD_OUT(4), B(3) => LMD_OUT(3), 
                           B(2) => LMD_OUT(2), B(1) => LMD_OUT(1), B(0) => 
                           LMD_OUT(0), S => WB_MUX_SEL, Y(31) => DATAIN_RF(31),
                           Y(30) => DATAIN_RF(30), Y(29) => DATAIN_RF(29), 
                           Y(28) => DATAIN_RF(28), Y(27) => DATAIN_RF(27), 
                           Y(26) => DATAIN_RF(26), Y(25) => DATAIN_RF(25), 
                           Y(24) => DATAIN_RF(24), Y(23) => DATAIN_RF(23), 
                           Y(22) => DATAIN_RF(22), Y(21) => DATAIN_RF(21), 
                           Y(20) => DATAIN_RF(20), Y(19) => DATAIN_RF(19), 
                           Y(18) => DATAIN_RF(18), Y(17) => DATAIN_RF(17), 
                           Y(16) => DATAIN_RF(16), Y(15) => DATAIN_RF(15), 
                           Y(14) => DATAIN_RF(14), Y(13) => DATAIN_RF(13), 
                           Y(12) => DATAIN_RF(12), Y(11) => DATAIN_RF(11), 
                           Y(10) => DATAIN_RF(10), Y(9) => DATAIN_RF(9), Y(8) 
                           => DATAIN_RF(8), Y(7) => DATAIN_RF(7), Y(6) => 
                           DATAIN_RF(6), Y(5) => DATAIN_RF(5), Y(4) => 
                           DATAIN_RF(4), Y(3) => DATAIN_RF(3), Y(2) => 
                           DATAIN_RF(2), Y(1) => DATAIN_RF(1), Y(0) => 
                           DATAIN_RF(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity memoryUnit_nbits32 is

   port( clk, rst, LMD_LATCH_EN, JUMP_EN : in std_logic;  DRAM_DATA, 
         ALUREG_OUTPUT, NPC_OUT : in std_logic_vector (31 downto 0);  COND_OUT 
         : in std_logic;  DRAM_DATAout, TO_PC_OUT, ALU_OUT2 : out 
         std_logic_vector (31 downto 0);  IR_IN4 : in std_logic_vector (31 
         downto 0);  IR_OUT4 : out std_logic_vector (31 downto 0));

end memoryUnit_nbits32;

architecture SYN_STRUCTURAL of memoryUnit_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component register_generic_nbits32_1
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_2
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_bits32_2
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, muxjmp_to_mux, n3 : std_logic;

begin
   DRAM_DATAout <= ( DRAM_DATA(31), DRAM_DATA(30), DRAM_DATA(29), DRAM_DATA(28)
      , DRAM_DATA(27), DRAM_DATA(26), DRAM_DATA(25), DRAM_DATA(24), 
      DRAM_DATA(23), DRAM_DATA(22), DRAM_DATA(21), DRAM_DATA(20), DRAM_DATA(19)
      , DRAM_DATA(18), DRAM_DATA(17), DRAM_DATA(16), DRAM_DATA(15), 
      DRAM_DATA(14), DRAM_DATA(13), DRAM_DATA(12), DRAM_DATA(11), DRAM_DATA(10)
      , DRAM_DATA(9), DRAM_DATA(8), DRAM_DATA(7), DRAM_DATA(6), DRAM_DATA(5), 
      DRAM_DATA(4), DRAM_DATA(3), DRAM_DATA(2), DRAM_DATA(1), DRAM_DATA(0) );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   JUMPMUX : MUX21 port map( A => COND_OUT, B => X_Logic0_port, S => JUMP_EN, Y
                           => muxjmp_to_mux);
   MUX_PC : MUX21_GENERIC_bits32_2 port map( A(31) => ALUREG_OUTPUT(31), A(30) 
                           => ALUREG_OUTPUT(30), A(29) => ALUREG_OUTPUT(29), 
                           A(28) => ALUREG_OUTPUT(28), A(27) => 
                           ALUREG_OUTPUT(27), A(26) => ALUREG_OUTPUT(26), A(25)
                           => ALUREG_OUTPUT(25), A(24) => ALUREG_OUTPUT(24), 
                           A(23) => ALUREG_OUTPUT(23), A(22) => 
                           ALUREG_OUTPUT(22), A(21) => ALUREG_OUTPUT(21), A(20)
                           => ALUREG_OUTPUT(20), A(19) => ALUREG_OUTPUT(19), 
                           A(18) => ALUREG_OUTPUT(18), A(17) => 
                           ALUREG_OUTPUT(17), A(16) => ALUREG_OUTPUT(16), A(15)
                           => ALUREG_OUTPUT(15), A(14) => ALUREG_OUTPUT(14), 
                           A(13) => ALUREG_OUTPUT(13), A(12) => 
                           ALUREG_OUTPUT(12), A(11) => ALUREG_OUTPUT(11), A(10)
                           => ALUREG_OUTPUT(10), A(9) => ALUREG_OUTPUT(9), A(8)
                           => ALUREG_OUTPUT(8), A(7) => ALUREG_OUTPUT(7), A(6) 
                           => ALUREG_OUTPUT(6), A(5) => ALUREG_OUTPUT(5), A(4) 
                           => ALUREG_OUTPUT(4), A(3) => ALUREG_OUTPUT(3), A(2) 
                           => ALUREG_OUTPUT(2), A(1) => ALUREG_OUTPUT(1), A(0) 
                           => ALUREG_OUTPUT(0), B(31) => NPC_OUT(31), B(30) => 
                           NPC_OUT(30), B(29) => NPC_OUT(29), B(28) => 
                           NPC_OUT(28), B(27) => NPC_OUT(27), B(26) => 
                           NPC_OUT(26), B(25) => NPC_OUT(25), B(24) => 
                           NPC_OUT(24), B(23) => NPC_OUT(23), B(22) => 
                           NPC_OUT(22), B(21) => NPC_OUT(21), B(20) => 
                           NPC_OUT(20), B(19) => NPC_OUT(19), B(18) => 
                           NPC_OUT(18), B(17) => NPC_OUT(17), B(16) => 
                           NPC_OUT(16), B(15) => NPC_OUT(15), B(14) => 
                           NPC_OUT(14), B(13) => NPC_OUT(13), B(12) => 
                           NPC_OUT(12), B(11) => NPC_OUT(11), B(10) => 
                           NPC_OUT(10), B(9) => NPC_OUT(9), B(8) => NPC_OUT(8),
                           B(7) => NPC_OUT(7), B(6) => NPC_OUT(6), B(5) => 
                           NPC_OUT(5), B(4) => NPC_OUT(4), B(3) => NPC_OUT(3), 
                           B(2) => NPC_OUT(2), B(1) => NPC_OUT(1), B(0) => 
                           NPC_OUT(0), S => muxjmp_to_mux, Y(31) => 
                           TO_PC_OUT(31), Y(30) => TO_PC_OUT(30), Y(29) => 
                           TO_PC_OUT(29), Y(28) => TO_PC_OUT(28), Y(27) => 
                           TO_PC_OUT(27), Y(26) => TO_PC_OUT(26), Y(25) => 
                           TO_PC_OUT(25), Y(24) => TO_PC_OUT(24), Y(23) => 
                           TO_PC_OUT(23), Y(22) => TO_PC_OUT(22), Y(21) => 
                           TO_PC_OUT(21), Y(20) => TO_PC_OUT(20), Y(19) => 
                           TO_PC_OUT(19), Y(18) => TO_PC_OUT(18), Y(17) => 
                           TO_PC_OUT(17), Y(16) => TO_PC_OUT(16), Y(15) => 
                           TO_PC_OUT(15), Y(14) => TO_PC_OUT(14), Y(13) => 
                           TO_PC_OUT(13), Y(12) => TO_PC_OUT(12), Y(11) => 
                           TO_PC_OUT(11), Y(10) => TO_PC_OUT(10), Y(9) => 
                           TO_PC_OUT(9), Y(8) => TO_PC_OUT(8), Y(7) => 
                           TO_PC_OUT(7), Y(6) => TO_PC_OUT(6), Y(5) => 
                           TO_PC_OUT(5), Y(4) => TO_PC_OUT(4), Y(3) => 
                           TO_PC_OUT(3), Y(2) => TO_PC_OUT(2), Y(1) => 
                           TO_PC_OUT(1), Y(0) => TO_PC_OUT(0));
   ALU_OUT2r : register_generic_nbits32_2 port map( data_in(31) => 
                           ALUREG_OUTPUT(31), data_in(30) => ALUREG_OUTPUT(30),
                           data_in(29) => ALUREG_OUTPUT(29), data_in(28) => 
                           ALUREG_OUTPUT(28), data_in(27) => ALUREG_OUTPUT(27),
                           data_in(26) => ALUREG_OUTPUT(26), data_in(25) => 
                           ALUREG_OUTPUT(25), data_in(24) => ALUREG_OUTPUT(24),
                           data_in(23) => ALUREG_OUTPUT(23), data_in(22) => 
                           ALUREG_OUTPUT(22), data_in(21) => ALUREG_OUTPUT(21),
                           data_in(20) => ALUREG_OUTPUT(20), data_in(19) => 
                           ALUREG_OUTPUT(19), data_in(18) => ALUREG_OUTPUT(18),
                           data_in(17) => ALUREG_OUTPUT(17), data_in(16) => 
                           ALUREG_OUTPUT(16), data_in(15) => ALUREG_OUTPUT(15),
                           data_in(14) => ALUREG_OUTPUT(14), data_in(13) => 
                           ALUREG_OUTPUT(13), data_in(12) => ALUREG_OUTPUT(12),
                           data_in(11) => ALUREG_OUTPUT(11), data_in(10) => 
                           ALUREG_OUTPUT(10), data_in(9) => ALUREG_OUTPUT(9), 
                           data_in(8) => ALUREG_OUTPUT(8), data_in(7) => 
                           ALUREG_OUTPUT(7), data_in(6) => ALUREG_OUTPUT(6), 
                           data_in(5) => ALUREG_OUTPUT(5), data_in(4) => 
                           ALUREG_OUTPUT(4), data_in(3) => ALUREG_OUTPUT(3), 
                           data_in(2) => ALUREG_OUTPUT(2), data_in(1) => 
                           ALUREG_OUTPUT(1), data_in(0) => ALUREG_OUTPUT(0), CK
                           => clk, RESET => n3, ENABLE => X_Logic1_port, 
                           data_out(31) => ALU_OUT2(31), data_out(30) => 
                           ALU_OUT2(30), data_out(29) => ALU_OUT2(29), 
                           data_out(28) => ALU_OUT2(28), data_out(27) => 
                           ALU_OUT2(27), data_out(26) => ALU_OUT2(26), 
                           data_out(25) => ALU_OUT2(25), data_out(24) => 
                           ALU_OUT2(24), data_out(23) => ALU_OUT2(23), 
                           data_out(22) => ALU_OUT2(22), data_out(21) => 
                           ALU_OUT2(21), data_out(20) => ALU_OUT2(20), 
                           data_out(19) => ALU_OUT2(19), data_out(18) => 
                           ALU_OUT2(18), data_out(17) => ALU_OUT2(17), 
                           data_out(16) => ALU_OUT2(16), data_out(15) => 
                           ALU_OUT2(15), data_out(14) => ALU_OUT2(14), 
                           data_out(13) => ALU_OUT2(13), data_out(12) => 
                           ALU_OUT2(12), data_out(11) => ALU_OUT2(11), 
                           data_out(10) => ALU_OUT2(10), data_out(9) => 
                           ALU_OUT2(9), data_out(8) => ALU_OUT2(8), data_out(7)
                           => ALU_OUT2(7), data_out(6) => ALU_OUT2(6), 
                           data_out(5) => ALU_OUT2(5), data_out(4) => 
                           ALU_OUT2(4), data_out(3) => ALU_OUT2(3), data_out(2)
                           => ALU_OUT2(2), data_out(1) => ALU_OUT2(1), 
                           data_out(0) => ALU_OUT2(0));
   IR4 : register_generic_nbits32_1 port map( data_in(31) => IR_IN4(31), 
                           data_in(30) => IR_IN4(30), data_in(29) => IR_IN4(29)
                           , data_in(28) => IR_IN4(28), data_in(27) => 
                           IR_IN4(27), data_in(26) => IR_IN4(26), data_in(25) 
                           => IR_IN4(25), data_in(24) => IR_IN4(24), 
                           data_in(23) => IR_IN4(23), data_in(22) => IR_IN4(22)
                           , data_in(21) => IR_IN4(21), data_in(20) => 
                           IR_IN4(20), data_in(19) => IR_IN4(19), data_in(18) 
                           => IR_IN4(18), data_in(17) => IR_IN4(17), 
                           data_in(16) => IR_IN4(16), data_in(15) => IR_IN4(15)
                           , data_in(14) => IR_IN4(14), data_in(13) => 
                           IR_IN4(13), data_in(12) => IR_IN4(12), data_in(11) 
                           => IR_IN4(11), data_in(10) => IR_IN4(10), data_in(9)
                           => IR_IN4(9), data_in(8) => IR_IN4(8), data_in(7) =>
                           IR_IN4(7), data_in(6) => IR_IN4(6), data_in(5) => 
                           IR_IN4(5), data_in(4) => IR_IN4(4), data_in(3) => 
                           IR_IN4(3), data_in(2) => IR_IN4(2), data_in(1) => 
                           IR_IN4(1), data_in(0) => IR_IN4(0), CK => clk, RESET
                           => n3, ENABLE => X_Logic1_port, data_out(31) => 
                           IR_OUT4(31), data_out(30) => IR_OUT4(30), 
                           data_out(29) => IR_OUT4(29), data_out(28) => 
                           IR_OUT4(28), data_out(27) => IR_OUT4(27), 
                           data_out(26) => IR_OUT4(26), data_out(25) => 
                           IR_OUT4(25), data_out(24) => IR_OUT4(24), 
                           data_out(23) => IR_OUT4(23), data_out(22) => 
                           IR_OUT4(22), data_out(21) => IR_OUT4(21), 
                           data_out(20) => IR_OUT4(20), data_out(19) => 
                           IR_OUT4(19), data_out(18) => IR_OUT4(18), 
                           data_out(17) => IR_OUT4(17), data_out(16) => 
                           IR_OUT4(16), data_out(15) => IR_OUT4(15), 
                           data_out(14) => IR_OUT4(14), data_out(13) => 
                           IR_OUT4(13), data_out(12) => IR_OUT4(12), 
                           data_out(11) => IR_OUT4(11), data_out(10) => 
                           IR_OUT4(10), data_out(9) => IR_OUT4(9), data_out(8) 
                           => IR_OUT4(8), data_out(7) => IR_OUT4(7), 
                           data_out(6) => IR_OUT4(6), data_out(5) => IR_OUT4(5)
                           , data_out(4) => IR_OUT4(4), data_out(3) => 
                           IR_OUT4(3), data_out(2) => IR_OUT4(2), data_out(1) 
                           => IR_OUT4(1), data_out(0) => IR_OUT4(0));
   U3 : BUF_X1 port map( A => rst, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity executionUnit_nbits32 is

   port( clk, rst, ALU_OUTREG_ENABLE, MUXA_SEL, MUXB_SEL, COND_ENABLE : in 
         std_logic;  ALU_BITS : in std_logic_vector (0 to 3);  NPC_OUT, A_out, 
         B_out, Imm_out : in std_logic_vector (31 downto 0);  ALUREG_OUTPUT : 
         out std_logic_vector (31 downto 0);  COND_OUT : out std_logic;  IR_IN3
         : in std_logic_vector (31 downto 0);  IR_OUT3, B_outreg : out 
         std_logic_vector (31 downto 0));

end executionUnit_nbits32;

architecture SYN_STRUCTURAL of executionUnit_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_0
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component XNOR_logic
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component alu_nbits32
      port( FUNC : in std_logic_vector (0 to 3);  A, B : in std_logic_vector 
            (31 downto 0);  OUTALU : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_3
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_4
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_5
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_bits32_3
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_bits32_0
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component ZERO_DEC_bits32
      port( data : in std_logic_vector (31 downto 0);  zero_detect : out 
            std_logic);
   end component;
   
   signal X_Logic1_port, ZERO_DEC_OUT, MUX1_OUT_31_port, MUX1_OUT_30_port, 
      MUX1_OUT_29_port, MUX1_OUT_28_port, MUX1_OUT_27_port, MUX1_OUT_26_port, 
      MUX1_OUT_25_port, MUX1_OUT_24_port, MUX1_OUT_23_port, MUX1_OUT_22_port, 
      MUX1_OUT_21_port, MUX1_OUT_20_port, MUX1_OUT_19_port, MUX1_OUT_18_port, 
      MUX1_OUT_17_port, MUX1_OUT_16_port, MUX1_OUT_15_port, MUX1_OUT_14_port, 
      MUX1_OUT_13_port, MUX1_OUT_12_port, MUX1_OUT_11_port, MUX1_OUT_10_port, 
      MUX1_OUT_9_port, MUX1_OUT_8_port, MUX1_OUT_7_port, MUX1_OUT_6_port, 
      MUX1_OUT_5_port, MUX1_OUT_4_port, MUX1_OUT_3_port, MUX1_OUT_2_port, 
      MUX1_OUT_1_port, MUX1_OUT_0_port, MUX2_OUT_31_port, MUX2_OUT_30_port, 
      MUX2_OUT_29_port, MUX2_OUT_28_port, MUX2_OUT_27_port, MUX2_OUT_26_port, 
      MUX2_OUT_25_port, MUX2_OUT_24_port, MUX2_OUT_23_port, MUX2_OUT_22_port, 
      MUX2_OUT_21_port, MUX2_OUT_20_port, MUX2_OUT_19_port, MUX2_OUT_18_port, 
      MUX2_OUT_17_port, MUX2_OUT_16_port, MUX2_OUT_15_port, MUX2_OUT_14_port, 
      MUX2_OUT_13_port, MUX2_OUT_12_port, MUX2_OUT_11_port, MUX2_OUT_10_port, 
      MUX2_OUT_9_port, MUX2_OUT_8_port, MUX2_OUT_7_port, MUX2_OUT_6_port, 
      MUX2_OUT_5_port, MUX2_OUT_4_port, MUX2_OUT_3_port, MUX2_OUT_2_port, 
      MUX2_OUT_1_port, MUX2_OUT_0_port, ALU_output_31_port, ALU_output_30_port,
      ALU_output_29_port, ALU_output_28_port, ALU_output_27_port, 
      ALU_output_26_port, ALU_output_25_port, ALU_output_24_port, 
      ALU_output_23_port, ALU_output_22_port, ALU_output_21_port, 
      ALU_output_20_port, ALU_output_19_port, ALU_output_18_port, 
      ALU_output_17_port, ALU_output_16_port, ALU_output_15_port, 
      ALU_output_14_port, ALU_output_13_port, ALU_output_12_port, 
      ALU_output_11_port, ALU_output_10_port, ALU_output_9_port, 
      ALU_output_8_port, ALU_output_7_port, ALU_output_6_port, 
      ALU_output_5_port, ALU_output_4_port, ALU_output_3_port, 
      ALU_output_2_port, ALU_output_1_port, ALU_output_0_port, XNOR_OUT, n3 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   zerodec : ZERO_DEC_bits32 port map( data(31) => A_out(31), data(30) => 
                           A_out(30), data(29) => A_out(29), data(28) => 
                           A_out(28), data(27) => A_out(27), data(26) => 
                           A_out(26), data(25) => A_out(25), data(24) => 
                           A_out(24), data(23) => A_out(23), data(22) => 
                           A_out(22), data(21) => A_out(21), data(20) => 
                           A_out(20), data(19) => A_out(19), data(18) => 
                           A_out(18), data(17) => A_out(17), data(16) => 
                           A_out(16), data(15) => A_out(15), data(14) => 
                           A_out(14), data(13) => A_out(13), data(12) => 
                           A_out(12), data(11) => A_out(11), data(10) => 
                           A_out(10), data(9) => A_out(9), data(8) => A_out(8),
                           data(7) => A_out(7), data(6) => A_out(6), data(5) =>
                           A_out(5), data(4) => A_out(4), data(3) => A_out(3), 
                           data(2) => A_out(2), data(1) => A_out(1), data(0) =>
                           A_out(0), zero_detect => ZERO_DEC_OUT);
   mux1 : MUX21_GENERIC_bits32_0 port map( A(31) => A_out(31), A(30) => 
                           A_out(30), A(29) => A_out(29), A(28) => A_out(28), 
                           A(27) => A_out(27), A(26) => A_out(26), A(25) => 
                           A_out(25), A(24) => A_out(24), A(23) => A_out(23), 
                           A(22) => A_out(22), A(21) => A_out(21), A(20) => 
                           A_out(20), A(19) => A_out(19), A(18) => A_out(18), 
                           A(17) => A_out(17), A(16) => A_out(16), A(15) => 
                           A_out(15), A(14) => A_out(14), A(13) => A_out(13), 
                           A(12) => A_out(12), A(11) => A_out(11), A(10) => 
                           A_out(10), A(9) => A_out(9), A(8) => A_out(8), A(7) 
                           => A_out(7), A(6) => A_out(6), A(5) => A_out(5), 
                           A(4) => A_out(4), A(3) => A_out(3), A(2) => A_out(2)
                           , A(1) => A_out(1), A(0) => A_out(0), B(31) => 
                           NPC_OUT(31), B(30) => NPC_OUT(30), B(29) => 
                           NPC_OUT(29), B(28) => NPC_OUT(28), B(27) => 
                           NPC_OUT(27), B(26) => NPC_OUT(26), B(25) => 
                           NPC_OUT(25), B(24) => NPC_OUT(24), B(23) => 
                           NPC_OUT(23), B(22) => NPC_OUT(22), B(21) => 
                           NPC_OUT(21), B(20) => NPC_OUT(20), B(19) => 
                           NPC_OUT(19), B(18) => NPC_OUT(18), B(17) => 
                           NPC_OUT(17), B(16) => NPC_OUT(16), B(15) => 
                           NPC_OUT(15), B(14) => NPC_OUT(14), B(13) => 
                           NPC_OUT(13), B(12) => NPC_OUT(12), B(11) => 
                           NPC_OUT(11), B(10) => NPC_OUT(10), B(9) => 
                           NPC_OUT(9), B(8) => NPC_OUT(8), B(7) => NPC_OUT(7), 
                           B(6) => NPC_OUT(6), B(5) => NPC_OUT(5), B(4) => 
                           NPC_OUT(4), B(3) => NPC_OUT(3), B(2) => NPC_OUT(2), 
                           B(1) => NPC_OUT(1), B(0) => NPC_OUT(0), S => 
                           MUXA_SEL, Y(31) => MUX1_OUT_31_port, Y(30) => 
                           MUX1_OUT_30_port, Y(29) => MUX1_OUT_29_port, Y(28) 
                           => MUX1_OUT_28_port, Y(27) => MUX1_OUT_27_port, 
                           Y(26) => MUX1_OUT_26_port, Y(25) => MUX1_OUT_25_port
                           , Y(24) => MUX1_OUT_24_port, Y(23) => 
                           MUX1_OUT_23_port, Y(22) => MUX1_OUT_22_port, Y(21) 
                           => MUX1_OUT_21_port, Y(20) => MUX1_OUT_20_port, 
                           Y(19) => MUX1_OUT_19_port, Y(18) => MUX1_OUT_18_port
                           , Y(17) => MUX1_OUT_17_port, Y(16) => 
                           MUX1_OUT_16_port, Y(15) => MUX1_OUT_15_port, Y(14) 
                           => MUX1_OUT_14_port, Y(13) => MUX1_OUT_13_port, 
                           Y(12) => MUX1_OUT_12_port, Y(11) => MUX1_OUT_11_port
                           , Y(10) => MUX1_OUT_10_port, Y(9) => MUX1_OUT_9_port
                           , Y(8) => MUX1_OUT_8_port, Y(7) => MUX1_OUT_7_port, 
                           Y(6) => MUX1_OUT_6_port, Y(5) => MUX1_OUT_5_port, 
                           Y(4) => MUX1_OUT_4_port, Y(3) => MUX1_OUT_3_port, 
                           Y(2) => MUX1_OUT_2_port, Y(1) => MUX1_OUT_1_port, 
                           Y(0) => MUX1_OUT_0_port);
   mux2 : MUX21_GENERIC_bits32_3 port map( A(31) => Imm_out(31), A(30) => 
                           Imm_out(30), A(29) => Imm_out(29), A(28) => 
                           Imm_out(28), A(27) => Imm_out(27), A(26) => 
                           Imm_out(26), A(25) => Imm_out(25), A(24) => 
                           Imm_out(24), A(23) => Imm_out(23), A(22) => 
                           Imm_out(22), A(21) => Imm_out(21), A(20) => 
                           Imm_out(20), A(19) => Imm_out(19), A(18) => 
                           Imm_out(18), A(17) => Imm_out(17), A(16) => 
                           Imm_out(16), A(15) => Imm_out(15), A(14) => 
                           Imm_out(14), A(13) => Imm_out(13), A(12) => 
                           Imm_out(12), A(11) => Imm_out(11), A(10) => 
                           Imm_out(10), A(9) => Imm_out(9), A(8) => Imm_out(8),
                           A(7) => Imm_out(7), A(6) => Imm_out(6), A(5) => 
                           Imm_out(5), A(4) => Imm_out(4), A(3) => Imm_out(3), 
                           A(2) => Imm_out(2), A(1) => Imm_out(1), A(0) => 
                           Imm_out(0), B(31) => B_out(31), B(30) => B_out(30), 
                           B(29) => B_out(29), B(28) => B_out(28), B(27) => 
                           B_out(27), B(26) => B_out(26), B(25) => B_out(25), 
                           B(24) => B_out(24), B(23) => B_out(23), B(22) => 
                           B_out(22), B(21) => B_out(21), B(20) => B_out(20), 
                           B(19) => B_out(19), B(18) => B_out(18), B(17) => 
                           B_out(17), B(16) => B_out(16), B(15) => B_out(15), 
                           B(14) => B_out(14), B(13) => B_out(13), B(12) => 
                           B_out(12), B(11) => B_out(11), B(10) => B_out(10), 
                           B(9) => B_out(9), B(8) => B_out(8), B(7) => B_out(7)
                           , B(6) => B_out(6), B(5) => B_out(5), B(4) => 
                           B_out(4), B(3) => B_out(3), B(2) => B_out(2), B(1) 
                           => B_out(1), B(0) => B_out(0), S => MUXB_SEL, Y(31) 
                           => MUX2_OUT_31_port, Y(30) => MUX2_OUT_30_port, 
                           Y(29) => MUX2_OUT_29_port, Y(28) => MUX2_OUT_28_port
                           , Y(27) => MUX2_OUT_27_port, Y(26) => 
                           MUX2_OUT_26_port, Y(25) => MUX2_OUT_25_port, Y(24) 
                           => MUX2_OUT_24_port, Y(23) => MUX2_OUT_23_port, 
                           Y(22) => MUX2_OUT_22_port, Y(21) => MUX2_OUT_21_port
                           , Y(20) => MUX2_OUT_20_port, Y(19) => 
                           MUX2_OUT_19_port, Y(18) => MUX2_OUT_18_port, Y(17) 
                           => MUX2_OUT_17_port, Y(16) => MUX2_OUT_16_port, 
                           Y(15) => MUX2_OUT_15_port, Y(14) => MUX2_OUT_14_port
                           , Y(13) => MUX2_OUT_13_port, Y(12) => 
                           MUX2_OUT_12_port, Y(11) => MUX2_OUT_11_port, Y(10) 
                           => MUX2_OUT_10_port, Y(9) => MUX2_OUT_9_port, Y(8) 
                           => MUX2_OUT_8_port, Y(7) => MUX2_OUT_7_port, Y(6) =>
                           MUX2_OUT_6_port, Y(5) => MUX2_OUT_5_port, Y(4) => 
                           MUX2_OUT_4_port, Y(3) => MUX2_OUT_3_port, Y(2) => 
                           MUX2_OUT_2_port, Y(1) => MUX2_OUT_1_port, Y(0) => 
                           MUX2_OUT_0_port);
   ALUoutput : register_generic_nbits32_5 port map( data_in(31) => 
                           ALU_output_31_port, data_in(30) => 
                           ALU_output_30_port, data_in(29) => 
                           ALU_output_29_port, data_in(28) => 
                           ALU_output_28_port, data_in(27) => 
                           ALU_output_27_port, data_in(26) => 
                           ALU_output_26_port, data_in(25) => 
                           ALU_output_25_port, data_in(24) => 
                           ALU_output_24_port, data_in(23) => 
                           ALU_output_23_port, data_in(22) => 
                           ALU_output_22_port, data_in(21) => 
                           ALU_output_21_port, data_in(20) => 
                           ALU_output_20_port, data_in(19) => 
                           ALU_output_19_port, data_in(18) => 
                           ALU_output_18_port, data_in(17) => 
                           ALU_output_17_port, data_in(16) => 
                           ALU_output_16_port, data_in(15) => 
                           ALU_output_15_port, data_in(14) => 
                           ALU_output_14_port, data_in(13) => 
                           ALU_output_13_port, data_in(12) => 
                           ALU_output_12_port, data_in(11) => 
                           ALU_output_11_port, data_in(10) => 
                           ALU_output_10_port, data_in(9) => ALU_output_9_port,
                           data_in(8) => ALU_output_8_port, data_in(7) => 
                           ALU_output_7_port, data_in(6) => ALU_output_6_port, 
                           data_in(5) => ALU_output_5_port, data_in(4) => 
                           ALU_output_4_port, data_in(3) => ALU_output_3_port, 
                           data_in(2) => ALU_output_2_port, data_in(1) => 
                           ALU_output_1_port, data_in(0) => ALU_output_0_port, 
                           CK => clk, RESET => n3, ENABLE => ALU_OUTREG_ENABLE,
                           data_out(31) => ALUREG_OUTPUT(31), data_out(30) => 
                           ALUREG_OUTPUT(30), data_out(29) => ALUREG_OUTPUT(29)
                           , data_out(28) => ALUREG_OUTPUT(28), data_out(27) =>
                           ALUREG_OUTPUT(27), data_out(26) => ALUREG_OUTPUT(26)
                           , data_out(25) => ALUREG_OUTPUT(25), data_out(24) =>
                           ALUREG_OUTPUT(24), data_out(23) => ALUREG_OUTPUT(23)
                           , data_out(22) => ALUREG_OUTPUT(22), data_out(21) =>
                           ALUREG_OUTPUT(21), data_out(20) => ALUREG_OUTPUT(20)
                           , data_out(19) => ALUREG_OUTPUT(19), data_out(18) =>
                           ALUREG_OUTPUT(18), data_out(17) => ALUREG_OUTPUT(17)
                           , data_out(16) => ALUREG_OUTPUT(16), data_out(15) =>
                           ALUREG_OUTPUT(15), data_out(14) => ALUREG_OUTPUT(14)
                           , data_out(13) => ALUREG_OUTPUT(13), data_out(12) =>
                           ALUREG_OUTPUT(12), data_out(11) => ALUREG_OUTPUT(11)
                           , data_out(10) => ALUREG_OUTPUT(10), data_out(9) => 
                           ALUREG_OUTPUT(9), data_out(8) => ALUREG_OUTPUT(8), 
                           data_out(7) => ALUREG_OUTPUT(7), data_out(6) => 
                           ALUREG_OUTPUT(6), data_out(5) => ALUREG_OUTPUT(5), 
                           data_out(4) => ALUREG_OUTPUT(4), data_out(3) => 
                           ALUREG_OUTPUT(3), data_out(2) => ALUREG_OUTPUT(2), 
                           data_out(1) => ALUREG_OUTPUT(1), data_out(0) => 
                           ALUREG_OUTPUT(0));
   IR3 : register_generic_nbits32_4 port map( data_in(31) => IR_IN3(31), 
                           data_in(30) => IR_IN3(30), data_in(29) => IR_IN3(29)
                           , data_in(28) => IR_IN3(28), data_in(27) => 
                           IR_IN3(27), data_in(26) => IR_IN3(26), data_in(25) 
                           => IR_IN3(25), data_in(24) => IR_IN3(24), 
                           data_in(23) => IR_IN3(23), data_in(22) => IR_IN3(22)
                           , data_in(21) => IR_IN3(21), data_in(20) => 
                           IR_IN3(20), data_in(19) => IR_IN3(19), data_in(18) 
                           => IR_IN3(18), data_in(17) => IR_IN3(17), 
                           data_in(16) => IR_IN3(16), data_in(15) => IR_IN3(15)
                           , data_in(14) => IR_IN3(14), data_in(13) => 
                           IR_IN3(13), data_in(12) => IR_IN3(12), data_in(11) 
                           => IR_IN3(11), data_in(10) => IR_IN3(10), data_in(9)
                           => IR_IN3(9), data_in(8) => IR_IN3(8), data_in(7) =>
                           IR_IN3(7), data_in(6) => IR_IN3(6), data_in(5) => 
                           IR_IN3(5), data_in(4) => IR_IN3(4), data_in(3) => 
                           IR_IN3(3), data_in(2) => IR_IN3(2), data_in(1) => 
                           IR_IN3(1), data_in(0) => IR_IN3(0), CK => clk, RESET
                           => n3, ENABLE => X_Logic1_port, data_out(31) => 
                           IR_OUT3(31), data_out(30) => IR_OUT3(30), 
                           data_out(29) => IR_OUT3(29), data_out(28) => 
                           IR_OUT3(28), data_out(27) => IR_OUT3(27), 
                           data_out(26) => IR_OUT3(26), data_out(25) => 
                           IR_OUT3(25), data_out(24) => IR_OUT3(24), 
                           data_out(23) => IR_OUT3(23), data_out(22) => 
                           IR_OUT3(22), data_out(21) => IR_OUT3(21), 
                           data_out(20) => IR_OUT3(20), data_out(19) => 
                           IR_OUT3(19), data_out(18) => IR_OUT3(18), 
                           data_out(17) => IR_OUT3(17), data_out(16) => 
                           IR_OUT3(16), data_out(15) => IR_OUT3(15), 
                           data_out(14) => IR_OUT3(14), data_out(13) => 
                           IR_OUT3(13), data_out(12) => IR_OUT3(12), 
                           data_out(11) => IR_OUT3(11), data_out(10) => 
                           IR_OUT3(10), data_out(9) => IR_OUT3(9), data_out(8) 
                           => IR_OUT3(8), data_out(7) => IR_OUT3(7), 
                           data_out(6) => IR_OUT3(6), data_out(5) => IR_OUT3(5)
                           , data_out(4) => IR_OUT3(4), data_out(3) => 
                           IR_OUT3(3), data_out(2) => IR_OUT3(2), data_out(1) 
                           => IR_OUT3(1), data_out(0) => IR_OUT3(0));
   B_outregister : register_generic_nbits32_3 port map( data_in(31) => 
                           B_out(31), data_in(30) => B_out(30), data_in(29) => 
                           B_out(29), data_in(28) => B_out(28), data_in(27) => 
                           B_out(27), data_in(26) => B_out(26), data_in(25) => 
                           B_out(25), data_in(24) => B_out(24), data_in(23) => 
                           B_out(23), data_in(22) => B_out(22), data_in(21) => 
                           B_out(21), data_in(20) => B_out(20), data_in(19) => 
                           B_out(19), data_in(18) => B_out(18), data_in(17) => 
                           B_out(17), data_in(16) => B_out(16), data_in(15) => 
                           B_out(15), data_in(14) => B_out(14), data_in(13) => 
                           B_out(13), data_in(12) => B_out(12), data_in(11) => 
                           B_out(11), data_in(10) => B_out(10), data_in(9) => 
                           B_out(9), data_in(8) => B_out(8), data_in(7) => 
                           B_out(7), data_in(6) => B_out(6), data_in(5) => 
                           B_out(5), data_in(4) => B_out(4), data_in(3) => 
                           B_out(3), data_in(2) => B_out(2), data_in(1) => 
                           B_out(1), data_in(0) => B_out(0), CK => clk, RESET 
                           => n3, ENABLE => X_Logic1_port, data_out(31) => 
                           B_outreg(31), data_out(30) => B_outreg(30), 
                           data_out(29) => B_outreg(29), data_out(28) => 
                           B_outreg(28), data_out(27) => B_outreg(27), 
                           data_out(26) => B_outreg(26), data_out(25) => 
                           B_outreg(25), data_out(24) => B_outreg(24), 
                           data_out(23) => B_outreg(23), data_out(22) => 
                           B_outreg(22), data_out(21) => B_outreg(21), 
                           data_out(20) => B_outreg(20), data_out(19) => 
                           B_outreg(19), data_out(18) => B_outreg(18), 
                           data_out(17) => B_outreg(17), data_out(16) => 
                           B_outreg(16), data_out(15) => B_outreg(15), 
                           data_out(14) => B_outreg(14), data_out(13) => 
                           B_outreg(13), data_out(12) => B_outreg(12), 
                           data_out(11) => B_outreg(11), data_out(10) => 
                           B_outreg(10), data_out(9) => B_outreg(9), 
                           data_out(8) => B_outreg(8), data_out(7) => 
                           B_outreg(7), data_out(6) => B_outreg(6), data_out(5)
                           => B_outreg(5), data_out(4) => B_outreg(4), 
                           data_out(3) => B_outreg(3), data_out(2) => 
                           B_outreg(2), data_out(1) => B_outreg(1), data_out(0)
                           => B_outreg(0));
   alu1 : alu_nbits32 port map( FUNC(0) => ALU_BITS(0), FUNC(1) => ALU_BITS(1),
                           FUNC(2) => ALU_BITS(2), FUNC(3) => ALU_BITS(3), 
                           A(31) => MUX1_OUT_31_port, A(30) => MUX1_OUT_30_port
                           , A(29) => MUX1_OUT_29_port, A(28) => 
                           MUX1_OUT_28_port, A(27) => MUX1_OUT_27_port, A(26) 
                           => MUX1_OUT_26_port, A(25) => MUX1_OUT_25_port, 
                           A(24) => MUX1_OUT_24_port, A(23) => MUX1_OUT_23_port
                           , A(22) => MUX1_OUT_22_port, A(21) => 
                           MUX1_OUT_21_port, A(20) => MUX1_OUT_20_port, A(19) 
                           => MUX1_OUT_19_port, A(18) => MUX1_OUT_18_port, 
                           A(17) => MUX1_OUT_17_port, A(16) => MUX1_OUT_16_port
                           , A(15) => MUX1_OUT_15_port, A(14) => 
                           MUX1_OUT_14_port, A(13) => MUX1_OUT_13_port, A(12) 
                           => MUX1_OUT_12_port, A(11) => MUX1_OUT_11_port, 
                           A(10) => MUX1_OUT_10_port, A(9) => MUX1_OUT_9_port, 
                           A(8) => MUX1_OUT_8_port, A(7) => MUX1_OUT_7_port, 
                           A(6) => MUX1_OUT_6_port, A(5) => MUX1_OUT_5_port, 
                           A(4) => MUX1_OUT_4_port, A(3) => MUX1_OUT_3_port, 
                           A(2) => MUX1_OUT_2_port, A(1) => MUX1_OUT_1_port, 
                           A(0) => MUX1_OUT_0_port, B(31) => MUX2_OUT_31_port, 
                           B(30) => MUX2_OUT_30_port, B(29) => MUX2_OUT_29_port
                           , B(28) => MUX2_OUT_28_port, B(27) => 
                           MUX2_OUT_27_port, B(26) => MUX2_OUT_26_port, B(25) 
                           => MUX2_OUT_25_port, B(24) => MUX2_OUT_24_port, 
                           B(23) => MUX2_OUT_23_port, B(22) => MUX2_OUT_22_port
                           , B(21) => MUX2_OUT_21_port, B(20) => 
                           MUX2_OUT_20_port, B(19) => MUX2_OUT_19_port, B(18) 
                           => MUX2_OUT_18_port, B(17) => MUX2_OUT_17_port, 
                           B(16) => MUX2_OUT_16_port, B(15) => MUX2_OUT_15_port
                           , B(14) => MUX2_OUT_14_port, B(13) => 
                           MUX2_OUT_13_port, B(12) => MUX2_OUT_12_port, B(11) 
                           => MUX2_OUT_11_port, B(10) => MUX2_OUT_10_port, B(9)
                           => MUX2_OUT_9_port, B(8) => MUX2_OUT_8_port, B(7) =>
                           MUX2_OUT_7_port, B(6) => MUX2_OUT_6_port, B(5) => 
                           MUX2_OUT_5_port, B(4) => MUX2_OUT_4_port, B(3) => 
                           MUX2_OUT_3_port, B(2) => MUX2_OUT_2_port, B(1) => 
                           MUX2_OUT_1_port, B(0) => MUX2_OUT_0_port, OUTALU(31)
                           => ALU_output_31_port, OUTALU(30) => 
                           ALU_output_30_port, OUTALU(29) => ALU_output_29_port
                           , OUTALU(28) => ALU_output_28_port, OUTALU(27) => 
                           ALU_output_27_port, OUTALU(26) => ALU_output_26_port
                           , OUTALU(25) => ALU_output_25_port, OUTALU(24) => 
                           ALU_output_24_port, OUTALU(23) => ALU_output_23_port
                           , OUTALU(22) => ALU_output_22_port, OUTALU(21) => 
                           ALU_output_21_port, OUTALU(20) => ALU_output_20_port
                           , OUTALU(19) => ALU_output_19_port, OUTALU(18) => 
                           ALU_output_18_port, OUTALU(17) => ALU_output_17_port
                           , OUTALU(16) => ALU_output_16_port, OUTALU(15) => 
                           ALU_output_15_port, OUTALU(14) => ALU_output_14_port
                           , OUTALU(13) => ALU_output_13_port, OUTALU(12) => 
                           ALU_output_12_port, OUTALU(11) => ALU_output_11_port
                           , OUTALU(10) => ALU_output_10_port, OUTALU(9) => 
                           ALU_output_9_port, OUTALU(8) => ALU_output_8_port, 
                           OUTALU(7) => ALU_output_7_port, OUTALU(6) => 
                           ALU_output_6_port, OUTALU(5) => ALU_output_5_port, 
                           OUTALU(4) => ALU_output_4_port, OUTALU(3) => 
                           ALU_output_3_port, OUTALU(2) => ALU_output_2_port, 
                           OUTALU(1) => ALU_output_1_port, OUTALU(0) => 
                           ALU_output_0_port);
   XNOR_2 : XNOR_logic port map( A => ZERO_DEC_OUT, B => COND_ENABLE, Y => 
                           XNOR_OUT);
   COND : FD_0 port map( D => XNOR_OUT, CK => clk, RESET => n3, ENABLE => 
                           X_Logic1_port, Q => COND_OUT);
   U2 : BUF_X1 port map( A => rst, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity decodeUnit_nbits32 is

   port( clk, rst, RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE : in 
         std_logic;  DATAIN, IR_OUT : in std_logic_vector (31 downto 0);  A_out
         , B_out, Imm_out : out std_logic_vector (31 downto 0);  IR_IN2 : in 
         std_logic_vector (31 downto 0);  IR_OUT2 : out std_logic_vector (31 
         downto 0);  NPC_IN : in std_logic_vector (31 downto 0);  NPC2_OUT : 
         out std_logic_vector (31 downto 0));

end decodeUnit_nbits32;

architecture SYN_STRUCTURAL of decodeUnit_nbits32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component REGISTER_FILE_NBITS32_NREGISTERS32
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component SIGN_EXT_bits16
      port( inputt : in std_logic_vector (15 downto 0);  outputt : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_6
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_7
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_8
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic1_port, signExtOut_31_port, signExtOut_30_port, 
      signExtOut_29_port, signExtOut_28_port, signExtOut_27_port, 
      signExtOut_26_port, signExtOut_25_port, signExtOut_24_port, 
      signExtOut_23_port, signExtOut_22_port, signExtOut_21_port, 
      signExtOut_20_port, signExtOut_19_port, signExtOut_18_port, 
      signExtOut_17_port, signExtOut_16_port, signExtOut_15_port, 
      signExtOut_14_port, signExtOut_13_port, signExtOut_12_port, 
      signExtOut_11_port, signExtOut_10_port, signExtOut_9_port, 
      signExtOut_8_port, signExtOut_7_port, signExtOut_6_port, 
      signExtOut_5_port, signExtOut_4_port, signExtOut_3_port, 
      signExtOut_2_port, signExtOut_1_port, signExtOut_0_port, n7, n8, n9, n10,
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20 : std_logic;

begin
   
   X_Logic1_port <= '1';
   U7 : NOR4_X2 port map( A1 => IR_IN2(28), A2 => IR_IN2(27), A3 => IR_IN2(26),
                           A4 => n13, ZN => n8);
   NPC2 : register_generic_nbits32_8 port map( data_in(31) => NPC_IN(31), 
                           data_in(30) => NPC_IN(30), data_in(29) => NPC_IN(29)
                           , data_in(28) => NPC_IN(28), data_in(27) => 
                           NPC_IN(27), data_in(26) => NPC_IN(26), data_in(25) 
                           => NPC_IN(25), data_in(24) => NPC_IN(24), 
                           data_in(23) => NPC_IN(23), data_in(22) => NPC_IN(22)
                           , data_in(21) => NPC_IN(21), data_in(20) => 
                           NPC_IN(20), data_in(19) => NPC_IN(19), data_in(18) 
                           => NPC_IN(18), data_in(17) => NPC_IN(17), 
                           data_in(16) => NPC_IN(16), data_in(15) => NPC_IN(15)
                           , data_in(14) => NPC_IN(14), data_in(13) => 
                           NPC_IN(13), data_in(12) => NPC_IN(12), data_in(11) 
                           => NPC_IN(11), data_in(10) => NPC_IN(10), data_in(9)
                           => NPC_IN(9), data_in(8) => NPC_IN(8), data_in(7) =>
                           NPC_IN(7), data_in(6) => NPC_IN(6), data_in(5) => 
                           NPC_IN(5), data_in(4) => NPC_IN(4), data_in(3) => 
                           NPC_IN(3), data_in(2) => NPC_IN(2), data_in(1) => 
                           NPC_IN(1), data_in(0) => NPC_IN(0), CK => clk, RESET
                           => n14, ENABLE => X_Logic1_port, data_out(31) => 
                           NPC2_OUT(31), data_out(30) => NPC2_OUT(30), 
                           data_out(29) => NPC2_OUT(29), data_out(28) => 
                           NPC2_OUT(28), data_out(27) => NPC2_OUT(27), 
                           data_out(26) => NPC2_OUT(26), data_out(25) => 
                           NPC2_OUT(25), data_out(24) => NPC2_OUT(24), 
                           data_out(23) => NPC2_OUT(23), data_out(22) => 
                           NPC2_OUT(22), data_out(21) => NPC2_OUT(21), 
                           data_out(20) => NPC2_OUT(20), data_out(19) => 
                           NPC2_OUT(19), data_out(18) => NPC2_OUT(18), 
                           data_out(17) => NPC2_OUT(17), data_out(16) => 
                           NPC2_OUT(16), data_out(15) => NPC2_OUT(15), 
                           data_out(14) => NPC2_OUT(14), data_out(13) => 
                           NPC2_OUT(13), data_out(12) => NPC2_OUT(12), 
                           data_out(11) => NPC2_OUT(11), data_out(10) => 
                           NPC2_OUT(10), data_out(9) => NPC2_OUT(9), 
                           data_out(8) => NPC2_OUT(8), data_out(7) => 
                           NPC2_OUT(7), data_out(6) => NPC2_OUT(6), data_out(5)
                           => NPC2_OUT(5), data_out(4) => NPC2_OUT(4), 
                           data_out(3) => NPC2_OUT(3), data_out(2) => 
                           NPC2_OUT(2), data_out(1) => NPC2_OUT(1), data_out(0)
                           => NPC2_OUT(0));
   Imm : register_generic_nbits32_7 port map( data_in(31) => signExtOut_31_port
                           , data_in(30) => signExtOut_30_port, data_in(29) => 
                           signExtOut_29_port, data_in(28) => 
                           signExtOut_28_port, data_in(27) => 
                           signExtOut_27_port, data_in(26) => 
                           signExtOut_26_port, data_in(25) => 
                           signExtOut_25_port, data_in(24) => 
                           signExtOut_24_port, data_in(23) => 
                           signExtOut_23_port, data_in(22) => 
                           signExtOut_22_port, data_in(21) => 
                           signExtOut_21_port, data_in(20) => 
                           signExtOut_20_port, data_in(19) => 
                           signExtOut_19_port, data_in(18) => 
                           signExtOut_18_port, data_in(17) => 
                           signExtOut_17_port, data_in(16) => 
                           signExtOut_16_port, data_in(15) => 
                           signExtOut_15_port, data_in(14) => 
                           signExtOut_14_port, data_in(13) => 
                           signExtOut_13_port, data_in(12) => 
                           signExtOut_12_port, data_in(11) => 
                           signExtOut_11_port, data_in(10) => 
                           signExtOut_10_port, data_in(9) => signExtOut_9_port,
                           data_in(8) => signExtOut_8_port, data_in(7) => 
                           signExtOut_7_port, data_in(6) => signExtOut_6_port, 
                           data_in(5) => signExtOut_5_port, data_in(4) => 
                           signExtOut_4_port, data_in(3) => signExtOut_3_port, 
                           data_in(2) => signExtOut_2_port, data_in(1) => 
                           signExtOut_1_port, data_in(0) => signExtOut_0_port, 
                           CK => clk, RESET => n14, ENABLE => RegIMM_LATCH_EN, 
                           data_out(31) => Imm_out(31), data_out(30) => 
                           Imm_out(30), data_out(29) => Imm_out(29), 
                           data_out(28) => Imm_out(28), data_out(27) => 
                           Imm_out(27), data_out(26) => Imm_out(26), 
                           data_out(25) => Imm_out(25), data_out(24) => 
                           Imm_out(24), data_out(23) => Imm_out(23), 
                           data_out(22) => Imm_out(22), data_out(21) => 
                           Imm_out(21), data_out(20) => Imm_out(20), 
                           data_out(19) => Imm_out(19), data_out(18) => 
                           Imm_out(18), data_out(17) => Imm_out(17), 
                           data_out(16) => Imm_out(16), data_out(15) => 
                           Imm_out(15), data_out(14) => Imm_out(14), 
                           data_out(13) => Imm_out(13), data_out(12) => 
                           Imm_out(12), data_out(11) => Imm_out(11), 
                           data_out(10) => Imm_out(10), data_out(9) => 
                           Imm_out(9), data_out(8) => Imm_out(8), data_out(7) 
                           => Imm_out(7), data_out(6) => Imm_out(6), 
                           data_out(5) => Imm_out(5), data_out(4) => Imm_out(4)
                           , data_out(3) => Imm_out(3), data_out(2) => 
                           Imm_out(2), data_out(1) => Imm_out(1), data_out(0) 
                           => Imm_out(0));
   IR2 : register_generic_nbits32_6 port map( data_in(31) => IR_OUT(31), 
                           data_in(30) => IR_OUT(30), data_in(29) => IR_OUT(29)
                           , data_in(28) => IR_OUT(28), data_in(27) => 
                           IR_OUT(27), data_in(26) => IR_OUT(26), data_in(25) 
                           => IR_OUT(25), data_in(24) => IR_OUT(24), 
                           data_in(23) => IR_OUT(23), data_in(22) => IR_OUT(22)
                           , data_in(21) => IR_OUT(21), data_in(20) => 
                           IR_OUT(20), data_in(19) => IR_OUT(19), data_in(18) 
                           => IR_OUT(18), data_in(17) => IR_OUT(17), 
                           data_in(16) => IR_OUT(16), data_in(15) => IR_OUT(15)
                           , data_in(14) => IR_OUT(14), data_in(13) => 
                           IR_OUT(13), data_in(12) => IR_OUT(12), data_in(11) 
                           => IR_OUT(11), data_in(10) => IR_OUT(10), data_in(9)
                           => IR_OUT(9), data_in(8) => IR_OUT(8), data_in(7) =>
                           IR_OUT(7), data_in(6) => IR_OUT(6), data_in(5) => 
                           IR_OUT(5), data_in(4) => IR_OUT(4), data_in(3) => 
                           IR_OUT(3), data_in(2) => IR_OUT(2), data_in(1) => 
                           IR_OUT(1), data_in(0) => IR_OUT(0), CK => clk, RESET
                           => n14, ENABLE => X_Logic1_port, data_out(31) => 
                           IR_OUT2(31), data_out(30) => IR_OUT2(30), 
                           data_out(29) => IR_OUT2(29), data_out(28) => 
                           IR_OUT2(28), data_out(27) => IR_OUT2(27), 
                           data_out(26) => IR_OUT2(26), data_out(25) => 
                           IR_OUT2(25), data_out(24) => IR_OUT2(24), 
                           data_out(23) => IR_OUT2(23), data_out(22) => 
                           IR_OUT2(22), data_out(21) => IR_OUT2(21), 
                           data_out(20) => IR_OUT2(20), data_out(19) => 
                           IR_OUT2(19), data_out(18) => IR_OUT2(18), 
                           data_out(17) => IR_OUT2(17), data_out(16) => 
                           IR_OUT2(16), data_out(15) => IR_OUT2(15), 
                           data_out(14) => IR_OUT2(14), data_out(13) => 
                           IR_OUT2(13), data_out(12) => IR_OUT2(12), 
                           data_out(11) => IR_OUT2(11), data_out(10) => 
                           IR_OUT2(10), data_out(9) => IR_OUT2(9), data_out(8) 
                           => IR_OUT2(8), data_out(7) => IR_OUT2(7), 
                           data_out(6) => IR_OUT2(6), data_out(5) => IR_OUT2(5)
                           , data_out(4) => IR_OUT2(4), data_out(3) => 
                           IR_OUT2(3), data_out(2) => IR_OUT2(2), data_out(1) 
                           => IR_OUT2(1), data_out(0) => IR_OUT2(0));
   Signext : SIGN_EXT_bits16 port map( inputt(15) => IR_OUT(15), inputt(14) => 
                           IR_OUT(14), inputt(13) => IR_OUT(13), inputt(12) => 
                           IR_OUT(12), inputt(11) => IR_OUT(11), inputt(10) => 
                           IR_OUT(10), inputt(9) => IR_OUT(9), inputt(8) => 
                           IR_OUT(8), inputt(7) => IR_OUT(7), inputt(6) => 
                           IR_OUT(6), inputt(5) => IR_OUT(5), inputt(4) => 
                           IR_OUT(4), inputt(3) => IR_OUT(3), inputt(2) => 
                           IR_OUT(2), inputt(1) => IR_OUT(1), inputt(0) => 
                           IR_OUT(0), outputt(31) => signExtOut_31_port, 
                           outputt(30) => signExtOut_30_port, outputt(29) => 
                           signExtOut_29_port, outputt(28) => 
                           signExtOut_28_port, outputt(27) => 
                           signExtOut_27_port, outputt(26) => 
                           signExtOut_26_port, outputt(25) => 
                           signExtOut_25_port, outputt(24) => 
                           signExtOut_24_port, outputt(23) => 
                           signExtOut_23_port, outputt(22) => 
                           signExtOut_22_port, outputt(21) => 
                           signExtOut_21_port, outputt(20) => 
                           signExtOut_20_port, outputt(19) => 
                           signExtOut_19_port, outputt(18) => 
                           signExtOut_18_port, outputt(17) => 
                           signExtOut_17_port, outputt(16) => 
                           signExtOut_16_port, outputt(15) => 
                           signExtOut_15_port, outputt(14) => 
                           signExtOut_14_port, outputt(13) => 
                           signExtOut_13_port, outputt(12) => 
                           signExtOut_12_port, outputt(11) => 
                           signExtOut_11_port, outputt(10) => 
                           signExtOut_10_port, outputt(9) => signExtOut_9_port,
                           outputt(8) => signExtOut_8_port, outputt(7) => 
                           signExtOut_7_port, outputt(6) => signExtOut_6_port, 
                           outputt(5) => signExtOut_5_port, outputt(4) => 
                           signExtOut_4_port, outputt(3) => signExtOut_3_port, 
                           outputt(2) => signExtOut_2_port, outputt(1) => 
                           signExtOut_1_port, outputt(0) => signExtOut_0_port);
   RF : REGISTER_FILE_NBITS32_NREGISTERS32 port map( CLK => clk, RESET => n14, 
                           ENABLE => X_Logic1_port, RD1 => X_Logic1_port, RD2 
                           => X_Logic1_port, WR => RF_WE, ADD_WR(4) => n19, 
                           ADD_WR(3) => n18, ADD_WR(2) => n17, ADD_WR(1) => n16
                           , ADD_WR(0) => n15, ADD_RD1(4) => IR_OUT(25), 
                           ADD_RD1(3) => IR_OUT(24), ADD_RD1(2) => IR_OUT(23), 
                           ADD_RD1(1) => IR_OUT(22), ADD_RD1(0) => IR_OUT(21), 
                           ADD_RD2(4) => IR_OUT(20), ADD_RD2(3) => IR_OUT(19), 
                           ADD_RD2(2) => IR_OUT(18), ADD_RD2(1) => IR_OUT(17), 
                           ADD_RD2(0) => IR_OUT(16), DATAIN(31) => DATAIN(31), 
                           DATAIN(30) => DATAIN(30), DATAIN(29) => DATAIN(29), 
                           DATAIN(28) => DATAIN(28), DATAIN(27) => DATAIN(27), 
                           DATAIN(26) => DATAIN(26), DATAIN(25) => DATAIN(25), 
                           DATAIN(24) => DATAIN(24), DATAIN(23) => DATAIN(23), 
                           DATAIN(22) => DATAIN(22), DATAIN(21) => DATAIN(21), 
                           DATAIN(20) => DATAIN(20), DATAIN(19) => DATAIN(19), 
                           DATAIN(18) => DATAIN(18), DATAIN(17) => DATAIN(17), 
                           DATAIN(16) => DATAIN(16), DATAIN(15) => DATAIN(15), 
                           DATAIN(14) => DATAIN(14), DATAIN(13) => DATAIN(13), 
                           DATAIN(12) => DATAIN(12), DATAIN(11) => DATAIN(11), 
                           DATAIN(10) => DATAIN(10), DATAIN(9) => DATAIN(9), 
                           DATAIN(8) => DATAIN(8), DATAIN(7) => DATAIN(7), 
                           DATAIN(6) => DATAIN(6), DATAIN(5) => DATAIN(5), 
                           DATAIN(4) => DATAIN(4), DATAIN(3) => DATAIN(3), 
                           DATAIN(2) => DATAIN(2), DATAIN(1) => DATAIN(1), 
                           DATAIN(0) => DATAIN(0), OUT1(31) => A_out(31), 
                           OUT1(30) => A_out(30), OUT1(29) => A_out(29), 
                           OUT1(28) => A_out(28), OUT1(27) => A_out(27), 
                           OUT1(26) => A_out(26), OUT1(25) => A_out(25), 
                           OUT1(24) => A_out(24), OUT1(23) => A_out(23), 
                           OUT1(22) => A_out(22), OUT1(21) => A_out(21), 
                           OUT1(20) => A_out(20), OUT1(19) => A_out(19), 
                           OUT1(18) => A_out(18), OUT1(17) => A_out(17), 
                           OUT1(16) => A_out(16), OUT1(15) => A_out(15), 
                           OUT1(14) => A_out(14), OUT1(13) => A_out(13), 
                           OUT1(12) => A_out(12), OUT1(11) => A_out(11), 
                           OUT1(10) => A_out(10), OUT1(9) => A_out(9), OUT1(8) 
                           => A_out(8), OUT1(7) => A_out(7), OUT1(6) => 
                           A_out(6), OUT1(5) => A_out(5), OUT1(4) => A_out(4), 
                           OUT1(3) => A_out(3), OUT1(2) => A_out(2), OUT1(1) =>
                           A_out(1), OUT1(0) => A_out(0), OUT2(31) => B_out(31)
                           , OUT2(30) => B_out(30), OUT2(29) => B_out(29), 
                           OUT2(28) => B_out(28), OUT2(27) => B_out(27), 
                           OUT2(26) => B_out(26), OUT2(25) => B_out(25), 
                           OUT2(24) => B_out(24), OUT2(23) => B_out(23), 
                           OUT2(22) => B_out(22), OUT2(21) => B_out(21), 
                           OUT2(20) => B_out(20), OUT2(19) => B_out(19), 
                           OUT2(18) => B_out(18), OUT2(17) => B_out(17), 
                           OUT2(16) => B_out(16), OUT2(15) => B_out(15), 
                           OUT2(14) => B_out(14), OUT2(13) => B_out(13), 
                           OUT2(12) => B_out(12), OUT2(11) => B_out(11), 
                           OUT2(10) => B_out(10), OUT2(9) => B_out(9), OUT2(8) 
                           => B_out(8), OUT2(7) => B_out(7), OUT2(6) => 
                           B_out(6), OUT2(5) => B_out(5), OUT2(4) => B_out(4), 
                           OUT2(3) => B_out(3), OUT2(2) => B_out(2), OUT2(1) =>
                           B_out(1), OUT2(0) => B_out(0));
   U2 : BUF_X1 port map( A => rst, Z => n14);
   U3 : INV_X1 port map( A => n8, ZN => n20);
   U4 : OR3_X1 port map( A1 => IR_IN2(31), A2 => IR_IN2(30), A3 => IR_IN2(29), 
                           ZN => n13);
   U5 : INV_X1 port map( A => n10, ZN => n17);
   U6 : AOI22_X1 port map( A1 => IR_IN2(18), A2 => n20, B1 => IR_IN2(13), B2 =>
                           n8, ZN => n10);
   U8 : INV_X1 port map( A => n12, ZN => n15);
   U9 : AOI22_X1 port map( A1 => IR_IN2(16), A2 => n20, B1 => IR_IN2(11), B2 =>
                           n8, ZN => n12);
   U10 : INV_X1 port map( A => n7, ZN => n19);
   U11 : AOI22_X1 port map( A1 => IR_IN2(20), A2 => n20, B1 => IR_IN2(15), B2 
                           => n8, ZN => n7);
   U12 : INV_X1 port map( A => n9, ZN => n18);
   U13 : AOI22_X1 port map( A1 => IR_IN2(19), A2 => n20, B1 => IR_IN2(14), B2 
                           => n8, ZN => n9);
   U14 : INV_X1 port map( A => n11, ZN => n16);
   U15 : AOI22_X1 port map( A1 => IR_IN2(17), A2 => n20, B1 => IR_IN2(12), B2 
                           => n8, ZN => n11);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity fetchUnit_nbits32 is

   port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 downto 
         0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN : in std_logic;  PC_IN : 
         in std_logic_vector (31 downto 0);  ADDRESS_IRAM, NPC_OUT, IR_OUT, 
         ADDERPC_OUT : out std_logic_vector (31 downto 0));

end fetchUnit_nbits32;

architecture SYN_STRUCTURAL of fetchUnit_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component register_generic_nbits32_9
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_10
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_0
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component RCA_NBITS32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ADDRESS_IRAM_31_port, 
      ADDRESS_IRAM_30_port, ADDRESS_IRAM_29_port, ADDRESS_IRAM_28_port, 
      ADDRESS_IRAM_27_port, ADDRESS_IRAM_26_port, ADDRESS_IRAM_25_port, 
      ADDRESS_IRAM_24_port, ADDRESS_IRAM_23_port, ADDRESS_IRAM_22_port, 
      ADDRESS_IRAM_21_port, ADDRESS_IRAM_20_port, ADDRESS_IRAM_19_port, 
      ADDRESS_IRAM_18_port, ADDRESS_IRAM_17_port, ADDRESS_IRAM_16_port, 
      ADDRESS_IRAM_15_port, ADDRESS_IRAM_14_port, ADDRESS_IRAM_13_port, 
      ADDRESS_IRAM_12_port, ADDRESS_IRAM_11_port, ADDRESS_IRAM_10_port, 
      ADDRESS_IRAM_9_port, ADDRESS_IRAM_8_port, ADDRESS_IRAM_7_port, 
      ADDRESS_IRAM_6_port, ADDRESS_IRAM_5_port, ADDRESS_IRAM_4_port, 
      ADDRESS_IRAM_3_port, ADDRESS_IRAM_2_port, ADDRESS_IRAM_1_port, 
      ADDRESS_IRAM_0_port, ADDERPC_OUT_31_port, ADDERPC_OUT_30_port, 
      ADDERPC_OUT_29_port, ADDERPC_OUT_28_port, ADDERPC_OUT_27_port, 
      ADDERPC_OUT_26_port, ADDERPC_OUT_25_port, ADDERPC_OUT_24_port, 
      ADDERPC_OUT_23_port, ADDERPC_OUT_22_port, ADDERPC_OUT_21_port, 
      ADDERPC_OUT_20_port, ADDERPC_OUT_19_port, ADDERPC_OUT_18_port, 
      ADDERPC_OUT_17_port, ADDERPC_OUT_16_port, ADDERPC_OUT_15_port, 
      ADDERPC_OUT_14_port, ADDERPC_OUT_13_port, ADDERPC_OUT_12_port, 
      ADDERPC_OUT_11_port, ADDERPC_OUT_10_port, ADDERPC_OUT_9_port, 
      ADDERPC_OUT_8_port, ADDERPC_OUT_7_port, ADDERPC_OUT_6_port, 
      ADDERPC_OUT_5_port, ADDERPC_OUT_4_port, ADDERPC_OUT_3_port, 
      ADDERPC_OUT_2_port, ADDERPC_OUT_1_port, ADDERPC_OUT_0_port, n3, n4, 
      n_1755 : std_logic;

begin
   ADDRESS_IRAM <= ( ADDRESS_IRAM_31_port, ADDRESS_IRAM_30_port, 
      ADDRESS_IRAM_29_port, ADDRESS_IRAM_28_port, ADDRESS_IRAM_27_port, 
      ADDRESS_IRAM_26_port, ADDRESS_IRAM_25_port, ADDRESS_IRAM_24_port, 
      ADDRESS_IRAM_23_port, ADDRESS_IRAM_22_port, ADDRESS_IRAM_21_port, 
      ADDRESS_IRAM_20_port, ADDRESS_IRAM_19_port, ADDRESS_IRAM_18_port, 
      ADDRESS_IRAM_17_port, ADDRESS_IRAM_16_port, ADDRESS_IRAM_15_port, 
      ADDRESS_IRAM_14_port, ADDRESS_IRAM_13_port, ADDRESS_IRAM_12_port, 
      ADDRESS_IRAM_11_port, ADDRESS_IRAM_10_port, ADDRESS_IRAM_9_port, 
      ADDRESS_IRAM_8_port, ADDRESS_IRAM_7_port, ADDRESS_IRAM_6_port, 
      ADDRESS_IRAM_5_port, ADDRESS_IRAM_4_port, ADDRESS_IRAM_3_port, 
      ADDRESS_IRAM_2_port, ADDRESS_IRAM_1_port, ADDRESS_IRAM_0_port );
   ADDERPC_OUT <= ( ADDERPC_OUT_31_port, ADDERPC_OUT_30_port, 
      ADDERPC_OUT_29_port, ADDERPC_OUT_28_port, ADDERPC_OUT_27_port, 
      ADDERPC_OUT_26_port, ADDERPC_OUT_25_port, ADDERPC_OUT_24_port, 
      ADDERPC_OUT_23_port, ADDERPC_OUT_22_port, ADDERPC_OUT_21_port, 
      ADDERPC_OUT_20_port, ADDERPC_OUT_19_port, ADDERPC_OUT_18_port, 
      ADDERPC_OUT_17_port, ADDERPC_OUT_16_port, ADDERPC_OUT_15_port, 
      ADDERPC_OUT_14_port, ADDERPC_OUT_13_port, ADDERPC_OUT_12_port, 
      ADDERPC_OUT_11_port, ADDERPC_OUT_10_port, ADDERPC_OUT_9_port, 
      ADDERPC_OUT_8_port, ADDERPC_OUT_7_port, ADDERPC_OUT_6_port, 
      ADDERPC_OUT_5_port, ADDERPC_OUT_4_port, ADDERPC_OUT_3_port, 
      ADDERPC_OUT_2_port, ADDERPC_OUT_1_port, ADDERPC_OUT_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADD : RCA_NBITS32 port map( A(31) => ADDRESS_IRAM_31_port, A(30) => 
                           ADDRESS_IRAM_30_port, A(29) => ADDRESS_IRAM_29_port,
                           A(28) => ADDRESS_IRAM_28_port, A(27) => 
                           ADDRESS_IRAM_27_port, A(26) => ADDRESS_IRAM_26_port,
                           A(25) => ADDRESS_IRAM_25_port, A(24) => 
                           ADDRESS_IRAM_24_port, A(23) => ADDRESS_IRAM_23_port,
                           A(22) => ADDRESS_IRAM_22_port, A(21) => 
                           ADDRESS_IRAM_21_port, A(20) => ADDRESS_IRAM_20_port,
                           A(19) => ADDRESS_IRAM_19_port, A(18) => 
                           ADDRESS_IRAM_18_port, A(17) => ADDRESS_IRAM_17_port,
                           A(16) => ADDRESS_IRAM_16_port, A(15) => 
                           ADDRESS_IRAM_15_port, A(14) => ADDRESS_IRAM_14_port,
                           A(13) => ADDRESS_IRAM_13_port, A(12) => 
                           ADDRESS_IRAM_12_port, A(11) => ADDRESS_IRAM_11_port,
                           A(10) => ADDRESS_IRAM_10_port, A(9) => 
                           ADDRESS_IRAM_9_port, A(8) => ADDRESS_IRAM_8_port, 
                           A(7) => ADDRESS_IRAM_7_port, A(6) => 
                           ADDRESS_IRAM_6_port, A(5) => ADDRESS_IRAM_5_port, 
                           A(4) => ADDRESS_IRAM_4_port, A(3) => 
                           ADDRESS_IRAM_3_port, A(2) => ADDRESS_IRAM_2_port, 
                           A(1) => ADDRESS_IRAM_1_port, A(0) => 
                           ADDRESS_IRAM_0_port, B(31) => X_Logic0_port, B(30) 
                           => X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic1_port, Ci => X_Logic0_port, S(31) => 
                           ADDERPC_OUT_31_port, S(30) => ADDERPC_OUT_30_port, 
                           S(29) => ADDERPC_OUT_29_port, S(28) => 
                           ADDERPC_OUT_28_port, S(27) => ADDERPC_OUT_27_port, 
                           S(26) => ADDERPC_OUT_26_port, S(25) => 
                           ADDERPC_OUT_25_port, S(24) => ADDERPC_OUT_24_port, 
                           S(23) => ADDERPC_OUT_23_port, S(22) => 
                           ADDERPC_OUT_22_port, S(21) => ADDERPC_OUT_21_port, 
                           S(20) => ADDERPC_OUT_20_port, S(19) => 
                           ADDERPC_OUT_19_port, S(18) => ADDERPC_OUT_18_port, 
                           S(17) => ADDERPC_OUT_17_port, S(16) => 
                           ADDERPC_OUT_16_port, S(15) => ADDERPC_OUT_15_port, 
                           S(14) => ADDERPC_OUT_14_port, S(13) => 
                           ADDERPC_OUT_13_port, S(12) => ADDERPC_OUT_12_port, 
                           S(11) => ADDERPC_OUT_11_port, S(10) => 
                           ADDERPC_OUT_10_port, S(9) => ADDERPC_OUT_9_port, 
                           S(8) => ADDERPC_OUT_8_port, S(7) => 
                           ADDERPC_OUT_7_port, S(6) => ADDERPC_OUT_6_port, S(5)
                           => ADDERPC_OUT_5_port, S(4) => ADDERPC_OUT_4_port, 
                           S(3) => ADDERPC_OUT_3_port, S(2) => 
                           ADDERPC_OUT_2_port, S(1) => ADDERPC_OUT_1_port, S(0)
                           => ADDERPC_OUT_0_port, Co => n_1755);
   PC : register_generic_nbits32_0 port map( data_in(31) => PC_IN(31), 
                           data_in(30) => PC_IN(30), data_in(29) => PC_IN(29), 
                           data_in(28) => PC_IN(28), data_in(27) => PC_IN(27), 
                           data_in(26) => PC_IN(26), data_in(25) => PC_IN(25), 
                           data_in(24) => PC_IN(24), data_in(23) => PC_IN(23), 
                           data_in(22) => PC_IN(22), data_in(21) => PC_IN(21), 
                           data_in(20) => PC_IN(20), data_in(19) => PC_IN(19), 
                           data_in(18) => PC_IN(18), data_in(17) => PC_IN(17), 
                           data_in(16) => PC_IN(16), data_in(15) => PC_IN(15), 
                           data_in(14) => PC_IN(14), data_in(13) => PC_IN(13), 
                           data_in(12) => PC_IN(12), data_in(11) => PC_IN(11), 
                           data_in(10) => PC_IN(10), data_in(9) => PC_IN(9), 
                           data_in(8) => PC_IN(8), data_in(7) => PC_IN(7), 
                           data_in(6) => PC_IN(6), data_in(5) => PC_IN(5), 
                           data_in(4) => PC_IN(4), data_in(3) => PC_IN(3), 
                           data_in(2) => PC_IN(2), data_in(1) => PC_IN(1), 
                           data_in(0) => PC_IN(0), CK => clk, RESET => n4, 
                           ENABLE => PC_LATCH_EN, data_out(31) => 
                           ADDRESS_IRAM_31_port, data_out(30) => 
                           ADDRESS_IRAM_30_port, data_out(29) => 
                           ADDRESS_IRAM_29_port, data_out(28) => 
                           ADDRESS_IRAM_28_port, data_out(27) => 
                           ADDRESS_IRAM_27_port, data_out(26) => 
                           ADDRESS_IRAM_26_port, data_out(25) => 
                           ADDRESS_IRAM_25_port, data_out(24) => 
                           ADDRESS_IRAM_24_port, data_out(23) => 
                           ADDRESS_IRAM_23_port, data_out(22) => 
                           ADDRESS_IRAM_22_port, data_out(21) => 
                           ADDRESS_IRAM_21_port, data_out(20) => 
                           ADDRESS_IRAM_20_port, data_out(19) => 
                           ADDRESS_IRAM_19_port, data_out(18) => 
                           ADDRESS_IRAM_18_port, data_out(17) => 
                           ADDRESS_IRAM_17_port, data_out(16) => 
                           ADDRESS_IRAM_16_port, data_out(15) => 
                           ADDRESS_IRAM_15_port, data_out(14) => 
                           ADDRESS_IRAM_14_port, data_out(13) => 
                           ADDRESS_IRAM_13_port, data_out(12) => 
                           ADDRESS_IRAM_12_port, data_out(11) => 
                           ADDRESS_IRAM_11_port, data_out(10) => 
                           ADDRESS_IRAM_10_port, data_out(9) => 
                           ADDRESS_IRAM_9_port, data_out(8) => 
                           ADDRESS_IRAM_8_port, data_out(7) => 
                           ADDRESS_IRAM_7_port, data_out(6) => 
                           ADDRESS_IRAM_6_port, data_out(5) => 
                           ADDRESS_IRAM_5_port, data_out(4) => 
                           ADDRESS_IRAM_4_port, data_out(3) => 
                           ADDRESS_IRAM_3_port, data_out(2) => 
                           ADDRESS_IRAM_2_port, data_out(1) => 
                           ADDRESS_IRAM_1_port, data_out(0) => 
                           ADDRESS_IRAM_0_port);
   IR : register_generic_nbits32_10 port map( data_in(31) => DATA_IRAM(31), 
                           data_in(30) => DATA_IRAM(30), data_in(29) => 
                           DATA_IRAM(29), data_in(28) => DATA_IRAM(28), 
                           data_in(27) => DATA_IRAM(27), data_in(26) => 
                           DATA_IRAM(26), data_in(25) => DATA_IRAM(25), 
                           data_in(24) => DATA_IRAM(24), data_in(23) => 
                           DATA_IRAM(23), data_in(22) => DATA_IRAM(22), 
                           data_in(21) => DATA_IRAM(21), data_in(20) => 
                           DATA_IRAM(20), data_in(19) => DATA_IRAM(19), 
                           data_in(18) => DATA_IRAM(18), data_in(17) => 
                           DATA_IRAM(17), data_in(16) => DATA_IRAM(16), 
                           data_in(15) => DATA_IRAM(15), data_in(14) => 
                           DATA_IRAM(14), data_in(13) => DATA_IRAM(13), 
                           data_in(12) => DATA_IRAM(12), data_in(11) => 
                           DATA_IRAM(11), data_in(10) => DATA_IRAM(10), 
                           data_in(9) => DATA_IRAM(9), data_in(8) => 
                           DATA_IRAM(8), data_in(7) => DATA_IRAM(7), data_in(6)
                           => DATA_IRAM(6), data_in(5) => DATA_IRAM(5), 
                           data_in(4) => DATA_IRAM(4), data_in(3) => 
                           DATA_IRAM(3), data_in(2) => DATA_IRAM(2), data_in(1)
                           => DATA_IRAM(1), data_in(0) => DATA_IRAM(0), CK => 
                           clk, RESET => n4, ENABLE => IR_LATCH_EN, 
                           data_out(31) => IR_OUT(31), data_out(30) => 
                           IR_OUT(30), data_out(29) => IR_OUT(29), data_out(28)
                           => IR_OUT(28), data_out(27) => IR_OUT(27), 
                           data_out(26) => IR_OUT(26), data_out(25) => 
                           IR_OUT(25), data_out(24) => IR_OUT(24), data_out(23)
                           => IR_OUT(23), data_out(22) => IR_OUT(22), 
                           data_out(21) => IR_OUT(21), data_out(20) => 
                           IR_OUT(20), data_out(19) => IR_OUT(19), data_out(18)
                           => IR_OUT(18), data_out(17) => IR_OUT(17), 
                           data_out(16) => IR_OUT(16), data_out(15) => 
                           IR_OUT(15), data_out(14) => IR_OUT(14), data_out(13)
                           => IR_OUT(13), data_out(12) => IR_OUT(12), 
                           data_out(11) => IR_OUT(11), data_out(10) => 
                           IR_OUT(10), data_out(9) => IR_OUT(9), data_out(8) =>
                           IR_OUT(8), data_out(7) => IR_OUT(7), data_out(6) => 
                           IR_OUT(6), data_out(5) => IR_OUT(5), data_out(4) => 
                           IR_OUT(4), data_out(3) => IR_OUT(3), data_out(2) => 
                           IR_OUT(2), data_out(1) => IR_OUT(1), data_out(0) => 
                           IR_OUT(0));
   NPC : register_generic_nbits32_9 port map( data_in(31) => n3, data_in(30) =>
                           ADDERPC_OUT_30_port, data_in(29) => 
                           ADDERPC_OUT_29_port, data_in(28) => 
                           ADDERPC_OUT_28_port, data_in(27) => 
                           ADDERPC_OUT_27_port, data_in(26) => 
                           ADDERPC_OUT_26_port, data_in(25) => 
                           ADDERPC_OUT_25_port, data_in(24) => 
                           ADDERPC_OUT_24_port, data_in(23) => 
                           ADDERPC_OUT_23_port, data_in(22) => 
                           ADDERPC_OUT_22_port, data_in(21) => 
                           ADDERPC_OUT_21_port, data_in(20) => 
                           ADDERPC_OUT_20_port, data_in(19) => 
                           ADDERPC_OUT_19_port, data_in(18) => 
                           ADDERPC_OUT_18_port, data_in(17) => 
                           ADDERPC_OUT_17_port, data_in(16) => 
                           ADDERPC_OUT_16_port, data_in(15) => 
                           ADDERPC_OUT_15_port, data_in(14) => 
                           ADDERPC_OUT_14_port, data_in(13) => 
                           ADDERPC_OUT_13_port, data_in(12) => 
                           ADDERPC_OUT_12_port, data_in(11) => 
                           ADDERPC_OUT_11_port, data_in(10) => 
                           ADDERPC_OUT_10_port, data_in(9) => 
                           ADDERPC_OUT_9_port, data_in(8) => ADDERPC_OUT_8_port
                           , data_in(7) => ADDERPC_OUT_7_port, data_in(6) => 
                           ADDERPC_OUT_6_port, data_in(5) => ADDERPC_OUT_5_port
                           , data_in(4) => ADDERPC_OUT_4_port, data_in(3) => 
                           ADDERPC_OUT_3_port, data_in(2) => ADDERPC_OUT_2_port
                           , data_in(1) => ADDERPC_OUT_1_port, data_in(0) => 
                           ADDERPC_OUT_0_port, CK => clk, RESET => n4, ENABLE 
                           => NPC_LATCH_EN, data_out(31) => NPC_OUT(31), 
                           data_out(30) => NPC_OUT(30), data_out(29) => 
                           NPC_OUT(29), data_out(28) => NPC_OUT(28), 
                           data_out(27) => NPC_OUT(27), data_out(26) => 
                           NPC_OUT(26), data_out(25) => NPC_OUT(25), 
                           data_out(24) => NPC_OUT(24), data_out(23) => 
                           NPC_OUT(23), data_out(22) => NPC_OUT(22), 
                           data_out(21) => NPC_OUT(21), data_out(20) => 
                           NPC_OUT(20), data_out(19) => NPC_OUT(19), 
                           data_out(18) => NPC_OUT(18), data_out(17) => 
                           NPC_OUT(17), data_out(16) => NPC_OUT(16), 
                           data_out(15) => NPC_OUT(15), data_out(14) => 
                           NPC_OUT(14), data_out(13) => NPC_OUT(13), 
                           data_out(12) => NPC_OUT(12), data_out(11) => 
                           NPC_OUT(11), data_out(10) => NPC_OUT(10), 
                           data_out(9) => NPC_OUT(9), data_out(8) => NPC_OUT(8)
                           , data_out(7) => NPC_OUT(7), data_out(6) => 
                           NPC_OUT(6), data_out(5) => NPC_OUT(5), data_out(4) 
                           => NPC_OUT(4), data_out(3) => NPC_OUT(3), 
                           data_out(2) => NPC_OUT(2), data_out(1) => NPC_OUT(1)
                           , data_out(0) => NPC_OUT(0));
   U3 : CLKBUF_X1 port map( A => ADDERPC_OUT_31_port, Z => n3);
   U4 : BUF_X1 port map( A => rst, Z => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity datapath_nbits32 is

   port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 downto 
         0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN, RegA_LATCH_EN, 
         RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE, MUXA_SEL, MUXB_SEL, 
         ALU_OUTREG_EN, EQ_COND : in std_logic;  ALU_OPCODE : in 
         std_logic_vector (0 to 3);  DRAM_DATA : in std_logic_vector (31 downto
         0);  LMD_LATCH_EN, JUMP_EN, WB_MUX_SEL : in std_logic;  B, ALU_OUT, 
         ADDRESS_IRAM, IR_OUT : out std_logic_vector (31 downto 0));

end datapath_nbits32;

architecture SYN_STRUCTURAL of datapath_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component writeBack_nbits32
      port( LMD_OUT, ALUREG_OUTPUT : in std_logic_vector (31 downto 0);  
            WB_MUX_SEL : in std_logic;  DATAIN_RF : out std_logic_vector (31 
            downto 0));
   end component;
   
   component memoryUnit_nbits32
      port( clk, rst, LMD_LATCH_EN, JUMP_EN : in std_logic;  DRAM_DATA, 
            ALUREG_OUTPUT, NPC_OUT : in std_logic_vector (31 downto 0);  
            COND_OUT : in std_logic;  DRAM_DATAout, TO_PC_OUT, ALU_OUT2 : out 
            std_logic_vector (31 downto 0);  IR_IN4 : in std_logic_vector (31 
            downto 0);  IR_OUT4 : out std_logic_vector (31 downto 0));
   end component;
   
   component executionUnit_nbits32
      port( clk, rst, ALU_OUTREG_ENABLE, MUXA_SEL, MUXB_SEL, COND_ENABLE : in 
            std_logic;  ALU_BITS : in std_logic_vector (0 to 3);  NPC_OUT, 
            A_out, B_out, Imm_out : in std_logic_vector (31 downto 0);  
            ALUREG_OUTPUT : out std_logic_vector (31 downto 0);  COND_OUT : out
            std_logic;  IR_IN3 : in std_logic_vector (31 downto 0);  IR_OUT3, 
            B_outreg : out std_logic_vector (31 downto 0));
   end component;
   
   component decodeUnit_nbits32
      port( clk, rst, RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE : in
            std_logic;  DATAIN, IR_OUT : in std_logic_vector (31 downto 0);  
            A_out, B_out, Imm_out : out std_logic_vector (31 downto 0);  IR_IN2
            : in std_logic_vector (31 downto 0);  IR_OUT2 : out 
            std_logic_vector (31 downto 0);  NPC_IN : in std_logic_vector (31 
            downto 0);  NPC2_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component fetchUnit_nbits32
      port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 
            downto 0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN : in std_logic; 
            PC_IN : in std_logic_vector (31 downto 0);  ADDRESS_IRAM, NPC_OUT, 
            IR_OUT, ADDERPC_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal ALU_OUT_31_port, ALU_OUT_30_port, ALU_OUT_29_port, ALU_OUT_28_port, 
      ALU_OUT_27_port, ALU_OUT_26_port, ALU_OUT_25_port, ALU_OUT_24_port, 
      ALU_OUT_23_port, ALU_OUT_22_port, ALU_OUT_21_port, ALU_OUT_20_port, 
      ALU_OUT_19_port, ALU_OUT_18_port, ALU_OUT_17_port, ALU_OUT_16_port, 
      ALU_OUT_15_port, ALU_OUT_14_port, ALU_OUT_13_port, ALU_OUT_12_port, 
      ALU_OUT_11_port, ALU_OUT_10_port, ALU_OUT_9_port, ALU_OUT_8_port, 
      ALU_OUT_7_port, ALU_OUT_6_port, ALU_OUT_5_port, ALU_OUT_4_port, 
      ALU_OUT_3_port, ALU_OUT_2_port, ALU_OUT_1_port, ALU_OUT_0_port, 
      IR_OUT_31_port, IR_OUT_30_port, IR_OUT_29_port, IR_OUT_28_port, 
      IR_OUT_27_port, IR_OUT_26_port, IR_OUT_25_port, IR_OUT_24_port, 
      IR_OUT_23_port, IR_OUT_22_port, IR_OUT_21_port, IR_OUT_20_port, 
      IR_OUT_19_port, IR_OUT_18_port, IR_OUT_17_port, IR_OUT_16_port, 
      IR_OUT_15_port, IR_OUT_14_port, IR_OUT_13_port, IR_OUT_12_port, 
      IR_OUT_11_port, IR_OUT_10_port, IR_OUT_9_port, IR_OUT_8_port, 
      IR_OUT_7_port, IR_OUT_6_port, IR_OUT_5_port, IR_OUT_4_port, IR_OUT_3_port
      , IR_OUT_2_port, IR_OUT_1_port, IR_OUT_0_port, TO_PC_OUTs_31_port, 
      TO_PC_OUTs_30_port, TO_PC_OUTs_29_port, TO_PC_OUTs_28_port, 
      TO_PC_OUTs_27_port, TO_PC_OUTs_26_port, TO_PC_OUTs_25_port, 
      TO_PC_OUTs_24_port, TO_PC_OUTs_23_port, TO_PC_OUTs_22_port, 
      TO_PC_OUTs_21_port, TO_PC_OUTs_20_port, TO_PC_OUTs_19_port, 
      TO_PC_OUTs_18_port, TO_PC_OUTs_17_port, TO_PC_OUTs_16_port, 
      TO_PC_OUTs_15_port, TO_PC_OUTs_14_port, TO_PC_OUTs_13_port, 
      TO_PC_OUTs_12_port, TO_PC_OUTs_11_port, TO_PC_OUTs_10_port, 
      TO_PC_OUTs_9_port, TO_PC_OUTs_8_port, TO_PC_OUTs_7_port, 
      TO_PC_OUTs_6_port, TO_PC_OUTs_5_port, TO_PC_OUTs_4_port, 
      TO_PC_OUTs_3_port, TO_PC_OUTs_2_port, TO_PC_OUTs_1_port, 
      TO_PC_OUTs_0_port, NPC_OUTs_31_port, NPC_OUTs_30_port, NPC_OUTs_29_port, 
      NPC_OUTs_28_port, NPC_OUTs_27_port, NPC_OUTs_26_port, NPC_OUTs_25_port, 
      NPC_OUTs_24_port, NPC_OUTs_23_port, NPC_OUTs_22_port, NPC_OUTs_21_port, 
      NPC_OUTs_20_port, NPC_OUTs_19_port, NPC_OUTs_18_port, NPC_OUTs_17_port, 
      NPC_OUTs_16_port, NPC_OUTs_15_port, NPC_OUTs_14_port, NPC_OUTs_13_port, 
      NPC_OUTs_12_port, NPC_OUTs_11_port, NPC_OUTs_10_port, NPC_OUTs_9_port, 
      NPC_OUTs_8_port, NPC_OUTs_7_port, NPC_OUTs_6_port, NPC_OUTs_5_port, 
      NPC_OUTs_4_port, NPC_OUTs_3_port, NPC_OUTs_2_port, NPC_OUTs_1_port, 
      NPC_OUTs_0_port, ADDERPC_OUTs_31_port, ADDERPC_OUTs_30_port, 
      ADDERPC_OUTs_29_port, ADDERPC_OUTs_28_port, ADDERPC_OUTs_27_port, 
      ADDERPC_OUTs_26_port, ADDERPC_OUTs_25_port, ADDERPC_OUTs_24_port, 
      ADDERPC_OUTs_23_port, ADDERPC_OUTs_22_port, ADDERPC_OUTs_21_port, 
      ADDERPC_OUTs_20_port, ADDERPC_OUTs_19_port, ADDERPC_OUTs_18_port, 
      ADDERPC_OUTs_17_port, ADDERPC_OUTs_16_port, ADDERPC_OUTs_15_port, 
      ADDERPC_OUTs_14_port, ADDERPC_OUTs_13_port, ADDERPC_OUTs_12_port, 
      ADDERPC_OUTs_11_port, ADDERPC_OUTs_10_port, ADDERPC_OUTs_9_port, 
      ADDERPC_OUTs_8_port, ADDERPC_OUTs_7_port, ADDERPC_OUTs_6_port, 
      ADDERPC_OUTs_5_port, ADDERPC_OUTs_4_port, ADDERPC_OUTs_3_port, 
      ADDERPC_OUTs_2_port, ADDERPC_OUTs_1_port, ADDERPC_OUTs_0_port, 
      DATAIN_RFs_31_port, DATAIN_RFs_30_port, DATAIN_RFs_29_port, 
      DATAIN_RFs_28_port, DATAIN_RFs_27_port, DATAIN_RFs_26_port, 
      DATAIN_RFs_25_port, DATAIN_RFs_24_port, DATAIN_RFs_23_port, 
      DATAIN_RFs_22_port, DATAIN_RFs_21_port, DATAIN_RFs_20_port, 
      DATAIN_RFs_19_port, DATAIN_RFs_18_port, DATAIN_RFs_17_port, 
      DATAIN_RFs_16_port, DATAIN_RFs_15_port, DATAIN_RFs_14_port, 
      DATAIN_RFs_13_port, DATAIN_RFs_12_port, DATAIN_RFs_11_port, 
      DATAIN_RFs_10_port, DATAIN_RFs_9_port, DATAIN_RFs_8_port, 
      DATAIN_RFs_7_port, DATAIN_RFs_6_port, DATAIN_RFs_5_port, 
      DATAIN_RFs_4_port, DATAIN_RFs_3_port, DATAIN_RFs_2_port, 
      DATAIN_RFs_1_port, DATAIN_RFs_0_port, A_outs_31_port, A_outs_30_port, 
      A_outs_29_port, A_outs_28_port, A_outs_27_port, A_outs_26_port, 
      A_outs_25_port, A_outs_24_port, A_outs_23_port, A_outs_22_port, 
      A_outs_21_port, A_outs_20_port, A_outs_19_port, A_outs_18_port, 
      A_outs_17_port, A_outs_16_port, A_outs_15_port, A_outs_14_port, 
      A_outs_13_port, A_outs_12_port, A_outs_11_port, A_outs_10_port, 
      A_outs_9_port, A_outs_8_port, A_outs_7_port, A_outs_6_port, A_outs_5_port
      , A_outs_4_port, A_outs_3_port, A_outs_2_port, A_outs_1_port, 
      A_outs_0_port, B_outs_31_port, B_outs_30_port, B_outs_29_port, 
      B_outs_28_port, B_outs_27_port, B_outs_26_port, B_outs_25_port, 
      B_outs_24_port, B_outs_23_port, B_outs_22_port, B_outs_21_port, 
      B_outs_20_port, B_outs_19_port, B_outs_18_port, B_outs_17_port, 
      B_outs_16_port, B_outs_15_port, B_outs_14_port, B_outs_13_port, 
      B_outs_12_port, B_outs_11_port, B_outs_10_port, B_outs_9_port, 
      B_outs_8_port, B_outs_7_port, B_outs_6_port, B_outs_5_port, B_outs_4_port
      , B_outs_3_port, B_outs_2_port, B_outs_1_port, B_outs_0_port, 
      Imm_outs_31_port, Imm_outs_30_port, Imm_outs_29_port, Imm_outs_28_port, 
      Imm_outs_27_port, Imm_outs_26_port, Imm_outs_25_port, Imm_outs_24_port, 
      Imm_outs_23_port, Imm_outs_22_port, Imm_outs_21_port, Imm_outs_20_port, 
      Imm_outs_19_port, Imm_outs_18_port, Imm_outs_17_port, Imm_outs_16_port, 
      Imm_outs_15_port, Imm_outs_14_port, Imm_outs_13_port, Imm_outs_12_port, 
      Imm_outs_11_port, Imm_outs_10_port, Imm_outs_9_port, Imm_outs_8_port, 
      Imm_outs_7_port, Imm_outs_6_port, Imm_outs_5_port, Imm_outs_4_port, 
      Imm_outs_3_port, Imm_outs_2_port, Imm_outs_1_port, Imm_outs_0_port, 
      IR_OUT4s_31_port, IR_OUT4s_30_port, IR_OUT4s_29_port, IR_OUT4s_28_port, 
      IR_OUT4s_27_port, IR_OUT4s_26_port, IR_OUT4s_25_port, IR_OUT4s_24_port, 
      IR_OUT4s_23_port, IR_OUT4s_22_port, IR_OUT4s_21_port, IR_OUT4s_20_port, 
      IR_OUT4s_19_port, IR_OUT4s_18_port, IR_OUT4s_17_port, IR_OUT4s_16_port, 
      IR_OUT4s_15_port, IR_OUT4s_14_port, IR_OUT4s_13_port, IR_OUT4s_12_port, 
      IR_OUT4s_11_port, IR_OUT4s_10_port, IR_OUT4s_9_port, IR_OUT4s_8_port, 
      IR_OUT4s_7_port, IR_OUT4s_6_port, IR_OUT4s_5_port, IR_OUT4s_4_port, 
      IR_OUT4s_3_port, IR_OUT4s_2_port, IR_OUT4s_1_port, IR_OUT4s_0_port, 
      IR_OUT2s_31_port, IR_OUT2s_30_port, IR_OUT2s_29_port, IR_OUT2s_28_port, 
      IR_OUT2s_27_port, IR_OUT2s_26_port, IR_OUT2s_25_port, IR_OUT2s_24_port, 
      IR_OUT2s_23_port, IR_OUT2s_22_port, IR_OUT2s_21_port, IR_OUT2s_20_port, 
      IR_OUT2s_19_port, IR_OUT2s_18_port, IR_OUT2s_17_port, IR_OUT2s_16_port, 
      IR_OUT2s_15_port, IR_OUT2s_14_port, IR_OUT2s_13_port, IR_OUT2s_12_port, 
      IR_OUT2s_11_port, IR_OUT2s_10_port, IR_OUT2s_9_port, IR_OUT2s_8_port, 
      IR_OUT2s_7_port, IR_OUT2s_6_port, IR_OUT2s_5_port, IR_OUT2s_4_port, 
      IR_OUT2s_3_port, IR_OUT2s_2_port, IR_OUT2s_1_port, IR_OUT2s_0_port, 
      NPC2_OUTs_31_port, NPC2_OUTs_30_port, NPC2_OUTs_29_port, 
      NPC2_OUTs_28_port, NPC2_OUTs_27_port, NPC2_OUTs_26_port, 
      NPC2_OUTs_25_port, NPC2_OUTs_24_port, NPC2_OUTs_23_port, 
      NPC2_OUTs_22_port, NPC2_OUTs_21_port, NPC2_OUTs_20_port, 
      NPC2_OUTs_19_port, NPC2_OUTs_18_port, NPC2_OUTs_17_port, 
      NPC2_OUTs_16_port, NPC2_OUTs_15_port, NPC2_OUTs_14_port, 
      NPC2_OUTs_13_port, NPC2_OUTs_12_port, NPC2_OUTs_11_port, 
      NPC2_OUTs_10_port, NPC2_OUTs_9_port, NPC2_OUTs_8_port, NPC2_OUTs_7_port, 
      NPC2_OUTs_6_port, NPC2_OUTs_5_port, NPC2_OUTs_4_port, NPC2_OUTs_3_port, 
      NPC2_OUTs_2_port, NPC2_OUTs_1_port, NPC2_OUTs_0_port, COND_OUTs, 
      IR_OUT3s_31_port, IR_OUT3s_30_port, IR_OUT3s_29_port, IR_OUT3s_28_port, 
      IR_OUT3s_27_port, IR_OUT3s_26_port, IR_OUT3s_25_port, IR_OUT3s_24_port, 
      IR_OUT3s_23_port, IR_OUT3s_22_port, IR_OUT3s_21_port, IR_OUT3s_20_port, 
      IR_OUT3s_19_port, IR_OUT3s_18_port, IR_OUT3s_17_port, IR_OUT3s_16_port, 
      IR_OUT3s_15_port, IR_OUT3s_14_port, IR_OUT3s_13_port, IR_OUT3s_12_port, 
      IR_OUT3s_11_port, IR_OUT3s_10_port, IR_OUT3s_9_port, IR_OUT3s_8_port, 
      IR_OUT3s_7_port, IR_OUT3s_6_port, IR_OUT3s_5_port, IR_OUT3s_4_port, 
      IR_OUT3s_3_port, IR_OUT3s_2_port, IR_OUT3s_1_port, IR_OUT3s_0_port, 
      LMD_OUTs_31_port, LMD_OUTs_30_port, LMD_OUTs_29_port, LMD_OUTs_28_port, 
      LMD_OUTs_27_port, LMD_OUTs_26_port, LMD_OUTs_25_port, LMD_OUTs_24_port, 
      LMD_OUTs_23_port, LMD_OUTs_22_port, LMD_OUTs_21_port, LMD_OUTs_20_port, 
      LMD_OUTs_19_port, LMD_OUTs_18_port, LMD_OUTs_17_port, LMD_OUTs_16_port, 
      LMD_OUTs_15_port, LMD_OUTs_14_port, LMD_OUTs_13_port, LMD_OUTs_12_port, 
      LMD_OUTs_11_port, LMD_OUTs_10_port, LMD_OUTs_9_port, LMD_OUTs_8_port, 
      LMD_OUTs_7_port, LMD_OUTs_6_port, LMD_OUTs_5_port, LMD_OUTs_4_port, 
      LMD_OUTs_3_port, LMD_OUTs_2_port, LMD_OUTs_1_port, LMD_OUTs_0_port, 
      ALU_OUT2s_31_port, ALU_OUT2s_30_port, ALU_OUT2s_29_port, 
      ALU_OUT2s_28_port, ALU_OUT2s_27_port, ALU_OUT2s_26_port, 
      ALU_OUT2s_25_port, ALU_OUT2s_24_port, ALU_OUT2s_23_port, 
      ALU_OUT2s_22_port, ALU_OUT2s_21_port, ALU_OUT2s_20_port, 
      ALU_OUT2s_19_port, ALU_OUT2s_18_port, ALU_OUT2s_17_port, 
      ALU_OUT2s_16_port, ALU_OUT2s_15_port, ALU_OUT2s_14_port, 
      ALU_OUT2s_13_port, ALU_OUT2s_12_port, ALU_OUT2s_11_port, 
      ALU_OUT2s_10_port, ALU_OUT2s_9_port, ALU_OUT2s_8_port, ALU_OUT2s_7_port, 
      ALU_OUT2s_6_port, ALU_OUT2s_5_port, ALU_OUT2s_4_port, ALU_OUT2s_3_port, 
      ALU_OUT2s_2_port, ALU_OUT2s_1_port, ALU_OUT2s_0_port, n3 : std_logic;

begin
   ALU_OUT <= ( ALU_OUT_31_port, ALU_OUT_30_port, ALU_OUT_29_port, 
      ALU_OUT_28_port, ALU_OUT_27_port, ALU_OUT_26_port, ALU_OUT_25_port, 
      ALU_OUT_24_port, ALU_OUT_23_port, ALU_OUT_22_port, ALU_OUT_21_port, 
      ALU_OUT_20_port, ALU_OUT_19_port, ALU_OUT_18_port, ALU_OUT_17_port, 
      ALU_OUT_16_port, ALU_OUT_15_port, ALU_OUT_14_port, ALU_OUT_13_port, 
      ALU_OUT_12_port, ALU_OUT_11_port, ALU_OUT_10_port, ALU_OUT_9_port, 
      ALU_OUT_8_port, ALU_OUT_7_port, ALU_OUT_6_port, ALU_OUT_5_port, 
      ALU_OUT_4_port, ALU_OUT_3_port, ALU_OUT_2_port, ALU_OUT_1_port, 
      ALU_OUT_0_port );
   IR_OUT <= ( IR_OUT_31_port, IR_OUT_30_port, IR_OUT_29_port, IR_OUT_28_port, 
      IR_OUT_27_port, IR_OUT_26_port, IR_OUT_25_port, IR_OUT_24_port, 
      IR_OUT_23_port, IR_OUT_22_port, IR_OUT_21_port, IR_OUT_20_port, 
      IR_OUT_19_port, IR_OUT_18_port, IR_OUT_17_port, IR_OUT_16_port, 
      IR_OUT_15_port, IR_OUT_14_port, IR_OUT_13_port, IR_OUT_12_port, 
      IR_OUT_11_port, IR_OUT_10_port, IR_OUT_9_port, IR_OUT_8_port, 
      IR_OUT_7_port, IR_OUT_6_port, IR_OUT_5_port, IR_OUT_4_port, IR_OUT_3_port
      , IR_OUT_2_port, IR_OUT_1_port, IR_OUT_0_port );
   
   FETCH : fetchUnit_nbits32 port map( clk => clk, rst => n3, DATA_IRAM(31) => 
                           DATA_IRAM(31), DATA_IRAM(30) => DATA_IRAM(30), 
                           DATA_IRAM(29) => DATA_IRAM(29), DATA_IRAM(28) => 
                           DATA_IRAM(28), DATA_IRAM(27) => DATA_IRAM(27), 
                           DATA_IRAM(26) => DATA_IRAM(26), DATA_IRAM(25) => 
                           DATA_IRAM(25), DATA_IRAM(24) => DATA_IRAM(24), 
                           DATA_IRAM(23) => DATA_IRAM(23), DATA_IRAM(22) => 
                           DATA_IRAM(22), DATA_IRAM(21) => DATA_IRAM(21), 
                           DATA_IRAM(20) => DATA_IRAM(20), DATA_IRAM(19) => 
                           DATA_IRAM(19), DATA_IRAM(18) => DATA_IRAM(18), 
                           DATA_IRAM(17) => DATA_IRAM(17), DATA_IRAM(16) => 
                           DATA_IRAM(16), DATA_IRAM(15) => DATA_IRAM(15), 
                           DATA_IRAM(14) => DATA_IRAM(14), DATA_IRAM(13) => 
                           DATA_IRAM(13), DATA_IRAM(12) => DATA_IRAM(12), 
                           DATA_IRAM(11) => DATA_IRAM(11), DATA_IRAM(10) => 
                           DATA_IRAM(10), DATA_IRAM(9) => DATA_IRAM(9), 
                           DATA_IRAM(8) => DATA_IRAM(8), DATA_IRAM(7) => 
                           DATA_IRAM(7), DATA_IRAM(6) => DATA_IRAM(6), 
                           DATA_IRAM(5) => DATA_IRAM(5), DATA_IRAM(4) => 
                           DATA_IRAM(4), DATA_IRAM(3) => DATA_IRAM(3), 
                           DATA_IRAM(2) => DATA_IRAM(2), DATA_IRAM(1) => 
                           DATA_IRAM(1), DATA_IRAM(0) => DATA_IRAM(0), 
                           IR_LATCH_EN => IR_LATCH_EN, NPC_LATCH_EN => 
                           NPC_LATCH_EN, PC_LATCH_EN => PC_LATCH_EN, PC_IN(31) 
                           => TO_PC_OUTs_31_port, PC_IN(30) => 
                           TO_PC_OUTs_30_port, PC_IN(29) => TO_PC_OUTs_29_port,
                           PC_IN(28) => TO_PC_OUTs_28_port, PC_IN(27) => 
                           TO_PC_OUTs_27_port, PC_IN(26) => TO_PC_OUTs_26_port,
                           PC_IN(25) => TO_PC_OUTs_25_port, PC_IN(24) => 
                           TO_PC_OUTs_24_port, PC_IN(23) => TO_PC_OUTs_23_port,
                           PC_IN(22) => TO_PC_OUTs_22_port, PC_IN(21) => 
                           TO_PC_OUTs_21_port, PC_IN(20) => TO_PC_OUTs_20_port,
                           PC_IN(19) => TO_PC_OUTs_19_port, PC_IN(18) => 
                           TO_PC_OUTs_18_port, PC_IN(17) => TO_PC_OUTs_17_port,
                           PC_IN(16) => TO_PC_OUTs_16_port, PC_IN(15) => 
                           TO_PC_OUTs_15_port, PC_IN(14) => TO_PC_OUTs_14_port,
                           PC_IN(13) => TO_PC_OUTs_13_port, PC_IN(12) => 
                           TO_PC_OUTs_12_port, PC_IN(11) => TO_PC_OUTs_11_port,
                           PC_IN(10) => TO_PC_OUTs_10_port, PC_IN(9) => 
                           TO_PC_OUTs_9_port, PC_IN(8) => TO_PC_OUTs_8_port, 
                           PC_IN(7) => TO_PC_OUTs_7_port, PC_IN(6) => 
                           TO_PC_OUTs_6_port, PC_IN(5) => TO_PC_OUTs_5_port, 
                           PC_IN(4) => TO_PC_OUTs_4_port, PC_IN(3) => 
                           TO_PC_OUTs_3_port, PC_IN(2) => TO_PC_OUTs_2_port, 
                           PC_IN(1) => TO_PC_OUTs_1_port, PC_IN(0) => 
                           TO_PC_OUTs_0_port, ADDRESS_IRAM(31) => 
                           ADDRESS_IRAM(31), ADDRESS_IRAM(30) => 
                           ADDRESS_IRAM(30), ADDRESS_IRAM(29) => 
                           ADDRESS_IRAM(29), ADDRESS_IRAM(28) => 
                           ADDRESS_IRAM(28), ADDRESS_IRAM(27) => 
                           ADDRESS_IRAM(27), ADDRESS_IRAM(26) => 
                           ADDRESS_IRAM(26), ADDRESS_IRAM(25) => 
                           ADDRESS_IRAM(25), ADDRESS_IRAM(24) => 
                           ADDRESS_IRAM(24), ADDRESS_IRAM(23) => 
                           ADDRESS_IRAM(23), ADDRESS_IRAM(22) => 
                           ADDRESS_IRAM(22), ADDRESS_IRAM(21) => 
                           ADDRESS_IRAM(21), ADDRESS_IRAM(20) => 
                           ADDRESS_IRAM(20), ADDRESS_IRAM(19) => 
                           ADDRESS_IRAM(19), ADDRESS_IRAM(18) => 
                           ADDRESS_IRAM(18), ADDRESS_IRAM(17) => 
                           ADDRESS_IRAM(17), ADDRESS_IRAM(16) => 
                           ADDRESS_IRAM(16), ADDRESS_IRAM(15) => 
                           ADDRESS_IRAM(15), ADDRESS_IRAM(14) => 
                           ADDRESS_IRAM(14), ADDRESS_IRAM(13) => 
                           ADDRESS_IRAM(13), ADDRESS_IRAM(12) => 
                           ADDRESS_IRAM(12), ADDRESS_IRAM(11) => 
                           ADDRESS_IRAM(11), ADDRESS_IRAM(10) => 
                           ADDRESS_IRAM(10), ADDRESS_IRAM(9) => ADDRESS_IRAM(9)
                           , ADDRESS_IRAM(8) => ADDRESS_IRAM(8), 
                           ADDRESS_IRAM(7) => ADDRESS_IRAM(7), ADDRESS_IRAM(6) 
                           => ADDRESS_IRAM(6), ADDRESS_IRAM(5) => 
                           ADDRESS_IRAM(5), ADDRESS_IRAM(4) => ADDRESS_IRAM(4),
                           ADDRESS_IRAM(3) => ADDRESS_IRAM(3), ADDRESS_IRAM(2) 
                           => ADDRESS_IRAM(2), ADDRESS_IRAM(1) => 
                           ADDRESS_IRAM(1), ADDRESS_IRAM(0) => ADDRESS_IRAM(0),
                           NPC_OUT(31) => NPC_OUTs_31_port, NPC_OUT(30) => 
                           NPC_OUTs_30_port, NPC_OUT(29) => NPC_OUTs_29_port, 
                           NPC_OUT(28) => NPC_OUTs_28_port, NPC_OUT(27) => 
                           NPC_OUTs_27_port, NPC_OUT(26) => NPC_OUTs_26_port, 
                           NPC_OUT(25) => NPC_OUTs_25_port, NPC_OUT(24) => 
                           NPC_OUTs_24_port, NPC_OUT(23) => NPC_OUTs_23_port, 
                           NPC_OUT(22) => NPC_OUTs_22_port, NPC_OUT(21) => 
                           NPC_OUTs_21_port, NPC_OUT(20) => NPC_OUTs_20_port, 
                           NPC_OUT(19) => NPC_OUTs_19_port, NPC_OUT(18) => 
                           NPC_OUTs_18_port, NPC_OUT(17) => NPC_OUTs_17_port, 
                           NPC_OUT(16) => NPC_OUTs_16_port, NPC_OUT(15) => 
                           NPC_OUTs_15_port, NPC_OUT(14) => NPC_OUTs_14_port, 
                           NPC_OUT(13) => NPC_OUTs_13_port, NPC_OUT(12) => 
                           NPC_OUTs_12_port, NPC_OUT(11) => NPC_OUTs_11_port, 
                           NPC_OUT(10) => NPC_OUTs_10_port, NPC_OUT(9) => 
                           NPC_OUTs_9_port, NPC_OUT(8) => NPC_OUTs_8_port, 
                           NPC_OUT(7) => NPC_OUTs_7_port, NPC_OUT(6) => 
                           NPC_OUTs_6_port, NPC_OUT(5) => NPC_OUTs_5_port, 
                           NPC_OUT(4) => NPC_OUTs_4_port, NPC_OUT(3) => 
                           NPC_OUTs_3_port, NPC_OUT(2) => NPC_OUTs_2_port, 
                           NPC_OUT(1) => NPC_OUTs_1_port, NPC_OUT(0) => 
                           NPC_OUTs_0_port, IR_OUT(31) => IR_OUT_31_port, 
                           IR_OUT(30) => IR_OUT_30_port, IR_OUT(29) => 
                           IR_OUT_29_port, IR_OUT(28) => IR_OUT_28_port, 
                           IR_OUT(27) => IR_OUT_27_port, IR_OUT(26) => 
                           IR_OUT_26_port, IR_OUT(25) => IR_OUT_25_port, 
                           IR_OUT(24) => IR_OUT_24_port, IR_OUT(23) => 
                           IR_OUT_23_port, IR_OUT(22) => IR_OUT_22_port, 
                           IR_OUT(21) => IR_OUT_21_port, IR_OUT(20) => 
                           IR_OUT_20_port, IR_OUT(19) => IR_OUT_19_port, 
                           IR_OUT(18) => IR_OUT_18_port, IR_OUT(17) => 
                           IR_OUT_17_port, IR_OUT(16) => IR_OUT_16_port, 
                           IR_OUT(15) => IR_OUT_15_port, IR_OUT(14) => 
                           IR_OUT_14_port, IR_OUT(13) => IR_OUT_13_port, 
                           IR_OUT(12) => IR_OUT_12_port, IR_OUT(11) => 
                           IR_OUT_11_port, IR_OUT(10) => IR_OUT_10_port, 
                           IR_OUT(9) => IR_OUT_9_port, IR_OUT(8) => 
                           IR_OUT_8_port, IR_OUT(7) => IR_OUT_7_port, IR_OUT(6)
                           => IR_OUT_6_port, IR_OUT(5) => IR_OUT_5_port, 
                           IR_OUT(4) => IR_OUT_4_port, IR_OUT(3) => 
                           IR_OUT_3_port, IR_OUT(2) => IR_OUT_2_port, IR_OUT(1)
                           => IR_OUT_1_port, IR_OUT(0) => IR_OUT_0_port, 
                           ADDERPC_OUT(31) => ADDERPC_OUTs_31_port, 
                           ADDERPC_OUT(30) => ADDERPC_OUTs_30_port, 
                           ADDERPC_OUT(29) => ADDERPC_OUTs_29_port, 
                           ADDERPC_OUT(28) => ADDERPC_OUTs_28_port, 
                           ADDERPC_OUT(27) => ADDERPC_OUTs_27_port, 
                           ADDERPC_OUT(26) => ADDERPC_OUTs_26_port, 
                           ADDERPC_OUT(25) => ADDERPC_OUTs_25_port, 
                           ADDERPC_OUT(24) => ADDERPC_OUTs_24_port, 
                           ADDERPC_OUT(23) => ADDERPC_OUTs_23_port, 
                           ADDERPC_OUT(22) => ADDERPC_OUTs_22_port, 
                           ADDERPC_OUT(21) => ADDERPC_OUTs_21_port, 
                           ADDERPC_OUT(20) => ADDERPC_OUTs_20_port, 
                           ADDERPC_OUT(19) => ADDERPC_OUTs_19_port, 
                           ADDERPC_OUT(18) => ADDERPC_OUTs_18_port, 
                           ADDERPC_OUT(17) => ADDERPC_OUTs_17_port, 
                           ADDERPC_OUT(16) => ADDERPC_OUTs_16_port, 
                           ADDERPC_OUT(15) => ADDERPC_OUTs_15_port, 
                           ADDERPC_OUT(14) => ADDERPC_OUTs_14_port, 
                           ADDERPC_OUT(13) => ADDERPC_OUTs_13_port, 
                           ADDERPC_OUT(12) => ADDERPC_OUTs_12_port, 
                           ADDERPC_OUT(11) => ADDERPC_OUTs_11_port, 
                           ADDERPC_OUT(10) => ADDERPC_OUTs_10_port, 
                           ADDERPC_OUT(9) => ADDERPC_OUTs_9_port, 
                           ADDERPC_OUT(8) => ADDERPC_OUTs_8_port, 
                           ADDERPC_OUT(7) => ADDERPC_OUTs_7_port, 
                           ADDERPC_OUT(6) => ADDERPC_OUTs_6_port, 
                           ADDERPC_OUT(5) => ADDERPC_OUTs_5_port, 
                           ADDERPC_OUT(4) => ADDERPC_OUTs_4_port, 
                           ADDERPC_OUT(3) => ADDERPC_OUTs_3_port, 
                           ADDERPC_OUT(2) => ADDERPC_OUTs_2_port, 
                           ADDERPC_OUT(1) => ADDERPC_OUTs_1_port, 
                           ADDERPC_OUT(0) => ADDERPC_OUTs_0_port);
   DECODE : decodeUnit_nbits32 port map( clk => clk, rst => n3, RegA_LATCH_EN 
                           => RegA_LATCH_EN, RegB_LATCH_EN => RegB_LATCH_EN, 
                           RegIMM_LATCH_EN => RegIMM_LATCH_EN, RF_WE => RF_WE, 
                           DATAIN(31) => DATAIN_RFs_31_port, DATAIN(30) => 
                           DATAIN_RFs_30_port, DATAIN(29) => DATAIN_RFs_29_port
                           , DATAIN(28) => DATAIN_RFs_28_port, DATAIN(27) => 
                           DATAIN_RFs_27_port, DATAIN(26) => DATAIN_RFs_26_port
                           , DATAIN(25) => DATAIN_RFs_25_port, DATAIN(24) => 
                           DATAIN_RFs_24_port, DATAIN(23) => DATAIN_RFs_23_port
                           , DATAIN(22) => DATAIN_RFs_22_port, DATAIN(21) => 
                           DATAIN_RFs_21_port, DATAIN(20) => DATAIN_RFs_20_port
                           , DATAIN(19) => DATAIN_RFs_19_port, DATAIN(18) => 
                           DATAIN_RFs_18_port, DATAIN(17) => DATAIN_RFs_17_port
                           , DATAIN(16) => DATAIN_RFs_16_port, DATAIN(15) => 
                           DATAIN_RFs_15_port, DATAIN(14) => DATAIN_RFs_14_port
                           , DATAIN(13) => DATAIN_RFs_13_port, DATAIN(12) => 
                           DATAIN_RFs_12_port, DATAIN(11) => DATAIN_RFs_11_port
                           , DATAIN(10) => DATAIN_RFs_10_port, DATAIN(9) => 
                           DATAIN_RFs_9_port, DATAIN(8) => DATAIN_RFs_8_port, 
                           DATAIN(7) => DATAIN_RFs_7_port, DATAIN(6) => 
                           DATAIN_RFs_6_port, DATAIN(5) => DATAIN_RFs_5_port, 
                           DATAIN(4) => DATAIN_RFs_4_port, DATAIN(3) => 
                           DATAIN_RFs_3_port, DATAIN(2) => DATAIN_RFs_2_port, 
                           DATAIN(1) => DATAIN_RFs_1_port, DATAIN(0) => 
                           DATAIN_RFs_0_port, IR_OUT(31) => IR_OUT_31_port, 
                           IR_OUT(30) => IR_OUT_30_port, IR_OUT(29) => 
                           IR_OUT_29_port, IR_OUT(28) => IR_OUT_28_port, 
                           IR_OUT(27) => IR_OUT_27_port, IR_OUT(26) => 
                           IR_OUT_26_port, IR_OUT(25) => IR_OUT_25_port, 
                           IR_OUT(24) => IR_OUT_24_port, IR_OUT(23) => 
                           IR_OUT_23_port, IR_OUT(22) => IR_OUT_22_port, 
                           IR_OUT(21) => IR_OUT_21_port, IR_OUT(20) => 
                           IR_OUT_20_port, IR_OUT(19) => IR_OUT_19_port, 
                           IR_OUT(18) => IR_OUT_18_port, IR_OUT(17) => 
                           IR_OUT_17_port, IR_OUT(16) => IR_OUT_16_port, 
                           IR_OUT(15) => IR_OUT_15_port, IR_OUT(14) => 
                           IR_OUT_14_port, IR_OUT(13) => IR_OUT_13_port, 
                           IR_OUT(12) => IR_OUT_12_port, IR_OUT(11) => 
                           IR_OUT_11_port, IR_OUT(10) => IR_OUT_10_port, 
                           IR_OUT(9) => IR_OUT_9_port, IR_OUT(8) => 
                           IR_OUT_8_port, IR_OUT(7) => IR_OUT_7_port, IR_OUT(6)
                           => IR_OUT_6_port, IR_OUT(5) => IR_OUT_5_port, 
                           IR_OUT(4) => IR_OUT_4_port, IR_OUT(3) => 
                           IR_OUT_3_port, IR_OUT(2) => IR_OUT_2_port, IR_OUT(1)
                           => IR_OUT_1_port, IR_OUT(0) => IR_OUT_0_port, 
                           A_out(31) => A_outs_31_port, A_out(30) => 
                           A_outs_30_port, A_out(29) => A_outs_29_port, 
                           A_out(28) => A_outs_28_port, A_out(27) => 
                           A_outs_27_port, A_out(26) => A_outs_26_port, 
                           A_out(25) => A_outs_25_port, A_out(24) => 
                           A_outs_24_port, A_out(23) => A_outs_23_port, 
                           A_out(22) => A_outs_22_port, A_out(21) => 
                           A_outs_21_port, A_out(20) => A_outs_20_port, 
                           A_out(19) => A_outs_19_port, A_out(18) => 
                           A_outs_18_port, A_out(17) => A_outs_17_port, 
                           A_out(16) => A_outs_16_port, A_out(15) => 
                           A_outs_15_port, A_out(14) => A_outs_14_port, 
                           A_out(13) => A_outs_13_port, A_out(12) => 
                           A_outs_12_port, A_out(11) => A_outs_11_port, 
                           A_out(10) => A_outs_10_port, A_out(9) => 
                           A_outs_9_port, A_out(8) => A_outs_8_port, A_out(7) 
                           => A_outs_7_port, A_out(6) => A_outs_6_port, 
                           A_out(5) => A_outs_5_port, A_out(4) => A_outs_4_port
                           , A_out(3) => A_outs_3_port, A_out(2) => 
                           A_outs_2_port, A_out(1) => A_outs_1_port, A_out(0) 
                           => A_outs_0_port, B_out(31) => B_outs_31_port, 
                           B_out(30) => B_outs_30_port, B_out(29) => 
                           B_outs_29_port, B_out(28) => B_outs_28_port, 
                           B_out(27) => B_outs_27_port, B_out(26) => 
                           B_outs_26_port, B_out(25) => B_outs_25_port, 
                           B_out(24) => B_outs_24_port, B_out(23) => 
                           B_outs_23_port, B_out(22) => B_outs_22_port, 
                           B_out(21) => B_outs_21_port, B_out(20) => 
                           B_outs_20_port, B_out(19) => B_outs_19_port, 
                           B_out(18) => B_outs_18_port, B_out(17) => 
                           B_outs_17_port, B_out(16) => B_outs_16_port, 
                           B_out(15) => B_outs_15_port, B_out(14) => 
                           B_outs_14_port, B_out(13) => B_outs_13_port, 
                           B_out(12) => B_outs_12_port, B_out(11) => 
                           B_outs_11_port, B_out(10) => B_outs_10_port, 
                           B_out(9) => B_outs_9_port, B_out(8) => B_outs_8_port
                           , B_out(7) => B_outs_7_port, B_out(6) => 
                           B_outs_6_port, B_out(5) => B_outs_5_port, B_out(4) 
                           => B_outs_4_port, B_out(3) => B_outs_3_port, 
                           B_out(2) => B_outs_2_port, B_out(1) => B_outs_1_port
                           , B_out(0) => B_outs_0_port, Imm_out(31) => 
                           Imm_outs_31_port, Imm_out(30) => Imm_outs_30_port, 
                           Imm_out(29) => Imm_outs_29_port, Imm_out(28) => 
                           Imm_outs_28_port, Imm_out(27) => Imm_outs_27_port, 
                           Imm_out(26) => Imm_outs_26_port, Imm_out(25) => 
                           Imm_outs_25_port, Imm_out(24) => Imm_outs_24_port, 
                           Imm_out(23) => Imm_outs_23_port, Imm_out(22) => 
                           Imm_outs_22_port, Imm_out(21) => Imm_outs_21_port, 
                           Imm_out(20) => Imm_outs_20_port, Imm_out(19) => 
                           Imm_outs_19_port, Imm_out(18) => Imm_outs_18_port, 
                           Imm_out(17) => Imm_outs_17_port, Imm_out(16) => 
                           Imm_outs_16_port, Imm_out(15) => Imm_outs_15_port, 
                           Imm_out(14) => Imm_outs_14_port, Imm_out(13) => 
                           Imm_outs_13_port, Imm_out(12) => Imm_outs_12_port, 
                           Imm_out(11) => Imm_outs_11_port, Imm_out(10) => 
                           Imm_outs_10_port, Imm_out(9) => Imm_outs_9_port, 
                           Imm_out(8) => Imm_outs_8_port, Imm_out(7) => 
                           Imm_outs_7_port, Imm_out(6) => Imm_outs_6_port, 
                           Imm_out(5) => Imm_outs_5_port, Imm_out(4) => 
                           Imm_outs_4_port, Imm_out(3) => Imm_outs_3_port, 
                           Imm_out(2) => Imm_outs_2_port, Imm_out(1) => 
                           Imm_outs_1_port, Imm_out(0) => Imm_outs_0_port, 
                           IR_IN2(31) => IR_OUT4s_31_port, IR_IN2(30) => 
                           IR_OUT4s_30_port, IR_IN2(29) => IR_OUT4s_29_port, 
                           IR_IN2(28) => IR_OUT4s_28_port, IR_IN2(27) => 
                           IR_OUT4s_27_port, IR_IN2(26) => IR_OUT4s_26_port, 
                           IR_IN2(25) => IR_OUT4s_25_port, IR_IN2(24) => 
                           IR_OUT4s_24_port, IR_IN2(23) => IR_OUT4s_23_port, 
                           IR_IN2(22) => IR_OUT4s_22_port, IR_IN2(21) => 
                           IR_OUT4s_21_port, IR_IN2(20) => IR_OUT4s_20_port, 
                           IR_IN2(19) => IR_OUT4s_19_port, IR_IN2(18) => 
                           IR_OUT4s_18_port, IR_IN2(17) => IR_OUT4s_17_port, 
                           IR_IN2(16) => IR_OUT4s_16_port, IR_IN2(15) => 
                           IR_OUT4s_15_port, IR_IN2(14) => IR_OUT4s_14_port, 
                           IR_IN2(13) => IR_OUT4s_13_port, IR_IN2(12) => 
                           IR_OUT4s_12_port, IR_IN2(11) => IR_OUT4s_11_port, 
                           IR_IN2(10) => IR_OUT4s_10_port, IR_IN2(9) => 
                           IR_OUT4s_9_port, IR_IN2(8) => IR_OUT4s_8_port, 
                           IR_IN2(7) => IR_OUT4s_7_port, IR_IN2(6) => 
                           IR_OUT4s_6_port, IR_IN2(5) => IR_OUT4s_5_port, 
                           IR_IN2(4) => IR_OUT4s_4_port, IR_IN2(3) => 
                           IR_OUT4s_3_port, IR_IN2(2) => IR_OUT4s_2_port, 
                           IR_IN2(1) => IR_OUT4s_1_port, IR_IN2(0) => 
                           IR_OUT4s_0_port, IR_OUT2(31) => IR_OUT2s_31_port, 
                           IR_OUT2(30) => IR_OUT2s_30_port, IR_OUT2(29) => 
                           IR_OUT2s_29_port, IR_OUT2(28) => IR_OUT2s_28_port, 
                           IR_OUT2(27) => IR_OUT2s_27_port, IR_OUT2(26) => 
                           IR_OUT2s_26_port, IR_OUT2(25) => IR_OUT2s_25_port, 
                           IR_OUT2(24) => IR_OUT2s_24_port, IR_OUT2(23) => 
                           IR_OUT2s_23_port, IR_OUT2(22) => IR_OUT2s_22_port, 
                           IR_OUT2(21) => IR_OUT2s_21_port, IR_OUT2(20) => 
                           IR_OUT2s_20_port, IR_OUT2(19) => IR_OUT2s_19_port, 
                           IR_OUT2(18) => IR_OUT2s_18_port, IR_OUT2(17) => 
                           IR_OUT2s_17_port, IR_OUT2(16) => IR_OUT2s_16_port, 
                           IR_OUT2(15) => IR_OUT2s_15_port, IR_OUT2(14) => 
                           IR_OUT2s_14_port, IR_OUT2(13) => IR_OUT2s_13_port, 
                           IR_OUT2(12) => IR_OUT2s_12_port, IR_OUT2(11) => 
                           IR_OUT2s_11_port, IR_OUT2(10) => IR_OUT2s_10_port, 
                           IR_OUT2(9) => IR_OUT2s_9_port, IR_OUT2(8) => 
                           IR_OUT2s_8_port, IR_OUT2(7) => IR_OUT2s_7_port, 
                           IR_OUT2(6) => IR_OUT2s_6_port, IR_OUT2(5) => 
                           IR_OUT2s_5_port, IR_OUT2(4) => IR_OUT2s_4_port, 
                           IR_OUT2(3) => IR_OUT2s_3_port, IR_OUT2(2) => 
                           IR_OUT2s_2_port, IR_OUT2(1) => IR_OUT2s_1_port, 
                           IR_OUT2(0) => IR_OUT2s_0_port, NPC_IN(31) => 
                           NPC_OUTs_31_port, NPC_IN(30) => NPC_OUTs_30_port, 
                           NPC_IN(29) => NPC_OUTs_29_port, NPC_IN(28) => 
                           NPC_OUTs_28_port, NPC_IN(27) => NPC_OUTs_27_port, 
                           NPC_IN(26) => NPC_OUTs_26_port, NPC_IN(25) => 
                           NPC_OUTs_25_port, NPC_IN(24) => NPC_OUTs_24_port, 
                           NPC_IN(23) => NPC_OUTs_23_port, NPC_IN(22) => 
                           NPC_OUTs_22_port, NPC_IN(21) => NPC_OUTs_21_port, 
                           NPC_IN(20) => NPC_OUTs_20_port, NPC_IN(19) => 
                           NPC_OUTs_19_port, NPC_IN(18) => NPC_OUTs_18_port, 
                           NPC_IN(17) => NPC_OUTs_17_port, NPC_IN(16) => 
                           NPC_OUTs_16_port, NPC_IN(15) => NPC_OUTs_15_port, 
                           NPC_IN(14) => NPC_OUTs_14_port, NPC_IN(13) => 
                           NPC_OUTs_13_port, NPC_IN(12) => NPC_OUTs_12_port, 
                           NPC_IN(11) => NPC_OUTs_11_port, NPC_IN(10) => 
                           NPC_OUTs_10_port, NPC_IN(9) => NPC_OUTs_9_port, 
                           NPC_IN(8) => NPC_OUTs_8_port, NPC_IN(7) => 
                           NPC_OUTs_7_port, NPC_IN(6) => NPC_OUTs_6_port, 
                           NPC_IN(5) => NPC_OUTs_5_port, NPC_IN(4) => 
                           NPC_OUTs_4_port, NPC_IN(3) => NPC_OUTs_3_port, 
                           NPC_IN(2) => NPC_OUTs_2_port, NPC_IN(1) => 
                           NPC_OUTs_1_port, NPC_IN(0) => NPC_OUTs_0_port, 
                           NPC2_OUT(31) => NPC2_OUTs_31_port, NPC2_OUT(30) => 
                           NPC2_OUTs_30_port, NPC2_OUT(29) => NPC2_OUTs_29_port
                           , NPC2_OUT(28) => NPC2_OUTs_28_port, NPC2_OUT(27) =>
                           NPC2_OUTs_27_port, NPC2_OUT(26) => NPC2_OUTs_26_port
                           , NPC2_OUT(25) => NPC2_OUTs_25_port, NPC2_OUT(24) =>
                           NPC2_OUTs_24_port, NPC2_OUT(23) => NPC2_OUTs_23_port
                           , NPC2_OUT(22) => NPC2_OUTs_22_port, NPC2_OUT(21) =>
                           NPC2_OUTs_21_port, NPC2_OUT(20) => NPC2_OUTs_20_port
                           , NPC2_OUT(19) => NPC2_OUTs_19_port, NPC2_OUT(18) =>
                           NPC2_OUTs_18_port, NPC2_OUT(17) => NPC2_OUTs_17_port
                           , NPC2_OUT(16) => NPC2_OUTs_16_port, NPC2_OUT(15) =>
                           NPC2_OUTs_15_port, NPC2_OUT(14) => NPC2_OUTs_14_port
                           , NPC2_OUT(13) => NPC2_OUTs_13_port, NPC2_OUT(12) =>
                           NPC2_OUTs_12_port, NPC2_OUT(11) => NPC2_OUTs_11_port
                           , NPC2_OUT(10) => NPC2_OUTs_10_port, NPC2_OUT(9) => 
                           NPC2_OUTs_9_port, NPC2_OUT(8) => NPC2_OUTs_8_port, 
                           NPC2_OUT(7) => NPC2_OUTs_7_port, NPC2_OUT(6) => 
                           NPC2_OUTs_6_port, NPC2_OUT(5) => NPC2_OUTs_5_port, 
                           NPC2_OUT(4) => NPC2_OUTs_4_port, NPC2_OUT(3) => 
                           NPC2_OUTs_3_port, NPC2_OUT(2) => NPC2_OUTs_2_port, 
                           NPC2_OUT(1) => NPC2_OUTs_1_port, NPC2_OUT(0) => 
                           NPC2_OUTs_0_port);
   EXECUTE : executionUnit_nbits32 port map( clk => clk, rst => n3, 
                           ALU_OUTREG_ENABLE => ALU_OUTREG_EN, MUXA_SEL => 
                           MUXA_SEL, MUXB_SEL => MUXB_SEL, COND_ENABLE => 
                           EQ_COND, ALU_BITS(0) => ALU_OPCODE(0), ALU_BITS(1) 
                           => ALU_OPCODE(1), ALU_BITS(2) => ALU_OPCODE(2), 
                           ALU_BITS(3) => ALU_OPCODE(3), NPC_OUT(31) => 
                           NPC2_OUTs_31_port, NPC_OUT(30) => NPC2_OUTs_30_port,
                           NPC_OUT(29) => NPC2_OUTs_29_port, NPC_OUT(28) => 
                           NPC2_OUTs_28_port, NPC_OUT(27) => NPC2_OUTs_27_port,
                           NPC_OUT(26) => NPC2_OUTs_26_port, NPC_OUT(25) => 
                           NPC2_OUTs_25_port, NPC_OUT(24) => NPC2_OUTs_24_port,
                           NPC_OUT(23) => NPC2_OUTs_23_port, NPC_OUT(22) => 
                           NPC2_OUTs_22_port, NPC_OUT(21) => NPC2_OUTs_21_port,
                           NPC_OUT(20) => NPC2_OUTs_20_port, NPC_OUT(19) => 
                           NPC2_OUTs_19_port, NPC_OUT(18) => NPC2_OUTs_18_port,
                           NPC_OUT(17) => NPC2_OUTs_17_port, NPC_OUT(16) => 
                           NPC2_OUTs_16_port, NPC_OUT(15) => NPC2_OUTs_15_port,
                           NPC_OUT(14) => NPC2_OUTs_14_port, NPC_OUT(13) => 
                           NPC2_OUTs_13_port, NPC_OUT(12) => NPC2_OUTs_12_port,
                           NPC_OUT(11) => NPC2_OUTs_11_port, NPC_OUT(10) => 
                           NPC2_OUTs_10_port, NPC_OUT(9) => NPC2_OUTs_9_port, 
                           NPC_OUT(8) => NPC2_OUTs_8_port, NPC_OUT(7) => 
                           NPC2_OUTs_7_port, NPC_OUT(6) => NPC2_OUTs_6_port, 
                           NPC_OUT(5) => NPC2_OUTs_5_port, NPC_OUT(4) => 
                           NPC2_OUTs_4_port, NPC_OUT(3) => NPC2_OUTs_3_port, 
                           NPC_OUT(2) => NPC2_OUTs_2_port, NPC_OUT(1) => 
                           NPC2_OUTs_1_port, NPC_OUT(0) => NPC2_OUTs_0_port, 
                           A_out(31) => A_outs_31_port, A_out(30) => 
                           A_outs_30_port, A_out(29) => A_outs_29_port, 
                           A_out(28) => A_outs_28_port, A_out(27) => 
                           A_outs_27_port, A_out(26) => A_outs_26_port, 
                           A_out(25) => A_outs_25_port, A_out(24) => 
                           A_outs_24_port, A_out(23) => A_outs_23_port, 
                           A_out(22) => A_outs_22_port, A_out(21) => 
                           A_outs_21_port, A_out(20) => A_outs_20_port, 
                           A_out(19) => A_outs_19_port, A_out(18) => 
                           A_outs_18_port, A_out(17) => A_outs_17_port, 
                           A_out(16) => A_outs_16_port, A_out(15) => 
                           A_outs_15_port, A_out(14) => A_outs_14_port, 
                           A_out(13) => A_outs_13_port, A_out(12) => 
                           A_outs_12_port, A_out(11) => A_outs_11_port, 
                           A_out(10) => A_outs_10_port, A_out(9) => 
                           A_outs_9_port, A_out(8) => A_outs_8_port, A_out(7) 
                           => A_outs_7_port, A_out(6) => A_outs_6_port, 
                           A_out(5) => A_outs_5_port, A_out(4) => A_outs_4_port
                           , A_out(3) => A_outs_3_port, A_out(2) => 
                           A_outs_2_port, A_out(1) => A_outs_1_port, A_out(0) 
                           => A_outs_0_port, B_out(31) => B_outs_31_port, 
                           B_out(30) => B_outs_30_port, B_out(29) => 
                           B_outs_29_port, B_out(28) => B_outs_28_port, 
                           B_out(27) => B_outs_27_port, B_out(26) => 
                           B_outs_26_port, B_out(25) => B_outs_25_port, 
                           B_out(24) => B_outs_24_port, B_out(23) => 
                           B_outs_23_port, B_out(22) => B_outs_22_port, 
                           B_out(21) => B_outs_21_port, B_out(20) => 
                           B_outs_20_port, B_out(19) => B_outs_19_port, 
                           B_out(18) => B_outs_18_port, B_out(17) => 
                           B_outs_17_port, B_out(16) => B_outs_16_port, 
                           B_out(15) => B_outs_15_port, B_out(14) => 
                           B_outs_14_port, B_out(13) => B_outs_13_port, 
                           B_out(12) => B_outs_12_port, B_out(11) => 
                           B_outs_11_port, B_out(10) => B_outs_10_port, 
                           B_out(9) => B_outs_9_port, B_out(8) => B_outs_8_port
                           , B_out(7) => B_outs_7_port, B_out(6) => 
                           B_outs_6_port, B_out(5) => B_outs_5_port, B_out(4) 
                           => B_outs_4_port, B_out(3) => B_outs_3_port, 
                           B_out(2) => B_outs_2_port, B_out(1) => B_outs_1_port
                           , B_out(0) => B_outs_0_port, Imm_out(31) => 
                           Imm_outs_31_port, Imm_out(30) => Imm_outs_30_port, 
                           Imm_out(29) => Imm_outs_29_port, Imm_out(28) => 
                           Imm_outs_28_port, Imm_out(27) => Imm_outs_27_port, 
                           Imm_out(26) => Imm_outs_26_port, Imm_out(25) => 
                           Imm_outs_25_port, Imm_out(24) => Imm_outs_24_port, 
                           Imm_out(23) => Imm_outs_23_port, Imm_out(22) => 
                           Imm_outs_22_port, Imm_out(21) => Imm_outs_21_port, 
                           Imm_out(20) => Imm_outs_20_port, Imm_out(19) => 
                           Imm_outs_19_port, Imm_out(18) => Imm_outs_18_port, 
                           Imm_out(17) => Imm_outs_17_port, Imm_out(16) => 
                           Imm_outs_16_port, Imm_out(15) => Imm_outs_15_port, 
                           Imm_out(14) => Imm_outs_14_port, Imm_out(13) => 
                           Imm_outs_13_port, Imm_out(12) => Imm_outs_12_port, 
                           Imm_out(11) => Imm_outs_11_port, Imm_out(10) => 
                           Imm_outs_10_port, Imm_out(9) => Imm_outs_9_port, 
                           Imm_out(8) => Imm_outs_8_port, Imm_out(7) => 
                           Imm_outs_7_port, Imm_out(6) => Imm_outs_6_port, 
                           Imm_out(5) => Imm_outs_5_port, Imm_out(4) => 
                           Imm_outs_4_port, Imm_out(3) => Imm_outs_3_port, 
                           Imm_out(2) => Imm_outs_2_port, Imm_out(1) => 
                           Imm_outs_1_port, Imm_out(0) => Imm_outs_0_port, 
                           ALUREG_OUTPUT(31) => ALU_OUT_31_port, 
                           ALUREG_OUTPUT(30) => ALU_OUT_30_port, 
                           ALUREG_OUTPUT(29) => ALU_OUT_29_port, 
                           ALUREG_OUTPUT(28) => ALU_OUT_28_port, 
                           ALUREG_OUTPUT(27) => ALU_OUT_27_port, 
                           ALUREG_OUTPUT(26) => ALU_OUT_26_port, 
                           ALUREG_OUTPUT(25) => ALU_OUT_25_port, 
                           ALUREG_OUTPUT(24) => ALU_OUT_24_port, 
                           ALUREG_OUTPUT(23) => ALU_OUT_23_port, 
                           ALUREG_OUTPUT(22) => ALU_OUT_22_port, 
                           ALUREG_OUTPUT(21) => ALU_OUT_21_port, 
                           ALUREG_OUTPUT(20) => ALU_OUT_20_port, 
                           ALUREG_OUTPUT(19) => ALU_OUT_19_port, 
                           ALUREG_OUTPUT(18) => ALU_OUT_18_port, 
                           ALUREG_OUTPUT(17) => ALU_OUT_17_port, 
                           ALUREG_OUTPUT(16) => ALU_OUT_16_port, 
                           ALUREG_OUTPUT(15) => ALU_OUT_15_port, 
                           ALUREG_OUTPUT(14) => ALU_OUT_14_port, 
                           ALUREG_OUTPUT(13) => ALU_OUT_13_port, 
                           ALUREG_OUTPUT(12) => ALU_OUT_12_port, 
                           ALUREG_OUTPUT(11) => ALU_OUT_11_port, 
                           ALUREG_OUTPUT(10) => ALU_OUT_10_port, 
                           ALUREG_OUTPUT(9) => ALU_OUT_9_port, ALUREG_OUTPUT(8)
                           => ALU_OUT_8_port, ALUREG_OUTPUT(7) => 
                           ALU_OUT_7_port, ALUREG_OUTPUT(6) => ALU_OUT_6_port, 
                           ALUREG_OUTPUT(5) => ALU_OUT_5_port, ALUREG_OUTPUT(4)
                           => ALU_OUT_4_port, ALUREG_OUTPUT(3) => 
                           ALU_OUT_3_port, ALUREG_OUTPUT(2) => ALU_OUT_2_port, 
                           ALUREG_OUTPUT(1) => ALU_OUT_1_port, ALUREG_OUTPUT(0)
                           => ALU_OUT_0_port, COND_OUT => COND_OUTs, IR_IN3(31)
                           => IR_OUT2s_31_port, IR_IN3(30) => IR_OUT2s_30_port,
                           IR_IN3(29) => IR_OUT2s_29_port, IR_IN3(28) => 
                           IR_OUT2s_28_port, IR_IN3(27) => IR_OUT2s_27_port, 
                           IR_IN3(26) => IR_OUT2s_26_port, IR_IN3(25) => 
                           IR_OUT2s_25_port, IR_IN3(24) => IR_OUT2s_24_port, 
                           IR_IN3(23) => IR_OUT2s_23_port, IR_IN3(22) => 
                           IR_OUT2s_22_port, IR_IN3(21) => IR_OUT2s_21_port, 
                           IR_IN3(20) => IR_OUT2s_20_port, IR_IN3(19) => 
                           IR_OUT2s_19_port, IR_IN3(18) => IR_OUT2s_18_port, 
                           IR_IN3(17) => IR_OUT2s_17_port, IR_IN3(16) => 
                           IR_OUT2s_16_port, IR_IN3(15) => IR_OUT2s_15_port, 
                           IR_IN3(14) => IR_OUT2s_14_port, IR_IN3(13) => 
                           IR_OUT2s_13_port, IR_IN3(12) => IR_OUT2s_12_port, 
                           IR_IN3(11) => IR_OUT2s_11_port, IR_IN3(10) => 
                           IR_OUT2s_10_port, IR_IN3(9) => IR_OUT2s_9_port, 
                           IR_IN3(8) => IR_OUT2s_8_port, IR_IN3(7) => 
                           IR_OUT2s_7_port, IR_IN3(6) => IR_OUT2s_6_port, 
                           IR_IN3(5) => IR_OUT2s_5_port, IR_IN3(4) => 
                           IR_OUT2s_4_port, IR_IN3(3) => IR_OUT2s_3_port, 
                           IR_IN3(2) => IR_OUT2s_2_port, IR_IN3(1) => 
                           IR_OUT2s_1_port, IR_IN3(0) => IR_OUT2s_0_port, 
                           IR_OUT3(31) => IR_OUT3s_31_port, IR_OUT3(30) => 
                           IR_OUT3s_30_port, IR_OUT3(29) => IR_OUT3s_29_port, 
                           IR_OUT3(28) => IR_OUT3s_28_port, IR_OUT3(27) => 
                           IR_OUT3s_27_port, IR_OUT3(26) => IR_OUT3s_26_port, 
                           IR_OUT3(25) => IR_OUT3s_25_port, IR_OUT3(24) => 
                           IR_OUT3s_24_port, IR_OUT3(23) => IR_OUT3s_23_port, 
                           IR_OUT3(22) => IR_OUT3s_22_port, IR_OUT3(21) => 
                           IR_OUT3s_21_port, IR_OUT3(20) => IR_OUT3s_20_port, 
                           IR_OUT3(19) => IR_OUT3s_19_port, IR_OUT3(18) => 
                           IR_OUT3s_18_port, IR_OUT3(17) => IR_OUT3s_17_port, 
                           IR_OUT3(16) => IR_OUT3s_16_port, IR_OUT3(15) => 
                           IR_OUT3s_15_port, IR_OUT3(14) => IR_OUT3s_14_port, 
                           IR_OUT3(13) => IR_OUT3s_13_port, IR_OUT3(12) => 
                           IR_OUT3s_12_port, IR_OUT3(11) => IR_OUT3s_11_port, 
                           IR_OUT3(10) => IR_OUT3s_10_port, IR_OUT3(9) => 
                           IR_OUT3s_9_port, IR_OUT3(8) => IR_OUT3s_8_port, 
                           IR_OUT3(7) => IR_OUT3s_7_port, IR_OUT3(6) => 
                           IR_OUT3s_6_port, IR_OUT3(5) => IR_OUT3s_5_port, 
                           IR_OUT3(4) => IR_OUT3s_4_port, IR_OUT3(3) => 
                           IR_OUT3s_3_port, IR_OUT3(2) => IR_OUT3s_2_port, 
                           IR_OUT3(1) => IR_OUT3s_1_port, IR_OUT3(0) => 
                           IR_OUT3s_0_port, B_outreg(31) => B(31), B_outreg(30)
                           => B(30), B_outreg(29) => B(29), B_outreg(28) => 
                           B(28), B_outreg(27) => B(27), B_outreg(26) => B(26),
                           B_outreg(25) => B(25), B_outreg(24) => B(24), 
                           B_outreg(23) => B(23), B_outreg(22) => B(22), 
                           B_outreg(21) => B(21), B_outreg(20) => B(20), 
                           B_outreg(19) => B(19), B_outreg(18) => B(18), 
                           B_outreg(17) => B(17), B_outreg(16) => B(16), 
                           B_outreg(15) => B(15), B_outreg(14) => B(14), 
                           B_outreg(13) => B(13), B_outreg(12) => B(12), 
                           B_outreg(11) => B(11), B_outreg(10) => B(10), 
                           B_outreg(9) => B(9), B_outreg(8) => B(8), 
                           B_outreg(7) => B(7), B_outreg(6) => B(6), 
                           B_outreg(5) => B(5), B_outreg(4) => B(4), 
                           B_outreg(3) => B(3), B_outreg(2) => B(2), 
                           B_outreg(1) => B(1), B_outreg(0) => B(0));
   MEMORY : memoryUnit_nbits32 port map( clk => clk, rst => n3, LMD_LATCH_EN =>
                           LMD_LATCH_EN, JUMP_EN => JUMP_EN, DRAM_DATA(31) => 
                           DRAM_DATA(31), DRAM_DATA(30) => DRAM_DATA(30), 
                           DRAM_DATA(29) => DRAM_DATA(29), DRAM_DATA(28) => 
                           DRAM_DATA(28), DRAM_DATA(27) => DRAM_DATA(27), 
                           DRAM_DATA(26) => DRAM_DATA(26), DRAM_DATA(25) => 
                           DRAM_DATA(25), DRAM_DATA(24) => DRAM_DATA(24), 
                           DRAM_DATA(23) => DRAM_DATA(23), DRAM_DATA(22) => 
                           DRAM_DATA(22), DRAM_DATA(21) => DRAM_DATA(21), 
                           DRAM_DATA(20) => DRAM_DATA(20), DRAM_DATA(19) => 
                           DRAM_DATA(19), DRAM_DATA(18) => DRAM_DATA(18), 
                           DRAM_DATA(17) => DRAM_DATA(17), DRAM_DATA(16) => 
                           DRAM_DATA(16), DRAM_DATA(15) => DRAM_DATA(15), 
                           DRAM_DATA(14) => DRAM_DATA(14), DRAM_DATA(13) => 
                           DRAM_DATA(13), DRAM_DATA(12) => DRAM_DATA(12), 
                           DRAM_DATA(11) => DRAM_DATA(11), DRAM_DATA(10) => 
                           DRAM_DATA(10), DRAM_DATA(9) => DRAM_DATA(9), 
                           DRAM_DATA(8) => DRAM_DATA(8), DRAM_DATA(7) => 
                           DRAM_DATA(7), DRAM_DATA(6) => DRAM_DATA(6), 
                           DRAM_DATA(5) => DRAM_DATA(5), DRAM_DATA(4) => 
                           DRAM_DATA(4), DRAM_DATA(3) => DRAM_DATA(3), 
                           DRAM_DATA(2) => DRAM_DATA(2), DRAM_DATA(1) => 
                           DRAM_DATA(1), DRAM_DATA(0) => DRAM_DATA(0), 
                           ALUREG_OUTPUT(31) => ALU_OUT_31_port, 
                           ALUREG_OUTPUT(30) => ALU_OUT_30_port, 
                           ALUREG_OUTPUT(29) => ALU_OUT_29_port, 
                           ALUREG_OUTPUT(28) => ALU_OUT_28_port, 
                           ALUREG_OUTPUT(27) => ALU_OUT_27_port, 
                           ALUREG_OUTPUT(26) => ALU_OUT_26_port, 
                           ALUREG_OUTPUT(25) => ALU_OUT_25_port, 
                           ALUREG_OUTPUT(24) => ALU_OUT_24_port, 
                           ALUREG_OUTPUT(23) => ALU_OUT_23_port, 
                           ALUREG_OUTPUT(22) => ALU_OUT_22_port, 
                           ALUREG_OUTPUT(21) => ALU_OUT_21_port, 
                           ALUREG_OUTPUT(20) => ALU_OUT_20_port, 
                           ALUREG_OUTPUT(19) => ALU_OUT_19_port, 
                           ALUREG_OUTPUT(18) => ALU_OUT_18_port, 
                           ALUREG_OUTPUT(17) => ALU_OUT_17_port, 
                           ALUREG_OUTPUT(16) => ALU_OUT_16_port, 
                           ALUREG_OUTPUT(15) => ALU_OUT_15_port, 
                           ALUREG_OUTPUT(14) => ALU_OUT_14_port, 
                           ALUREG_OUTPUT(13) => ALU_OUT_13_port, 
                           ALUREG_OUTPUT(12) => ALU_OUT_12_port, 
                           ALUREG_OUTPUT(11) => ALU_OUT_11_port, 
                           ALUREG_OUTPUT(10) => ALU_OUT_10_port, 
                           ALUREG_OUTPUT(9) => ALU_OUT_9_port, ALUREG_OUTPUT(8)
                           => ALU_OUT_8_port, ALUREG_OUTPUT(7) => 
                           ALU_OUT_7_port, ALUREG_OUTPUT(6) => ALU_OUT_6_port, 
                           ALUREG_OUTPUT(5) => ALU_OUT_5_port, ALUREG_OUTPUT(4)
                           => ALU_OUT_4_port, ALUREG_OUTPUT(3) => 
                           ALU_OUT_3_port, ALUREG_OUTPUT(2) => ALU_OUT_2_port, 
                           ALUREG_OUTPUT(1) => ALU_OUT_1_port, ALUREG_OUTPUT(0)
                           => ALU_OUT_0_port, NPC_OUT(31) => 
                           ADDERPC_OUTs_31_port, NPC_OUT(30) => 
                           ADDERPC_OUTs_30_port, NPC_OUT(29) => 
                           ADDERPC_OUTs_29_port, NPC_OUT(28) => 
                           ADDERPC_OUTs_28_port, NPC_OUT(27) => 
                           ADDERPC_OUTs_27_port, NPC_OUT(26) => 
                           ADDERPC_OUTs_26_port, NPC_OUT(25) => 
                           ADDERPC_OUTs_25_port, NPC_OUT(24) => 
                           ADDERPC_OUTs_24_port, NPC_OUT(23) => 
                           ADDERPC_OUTs_23_port, NPC_OUT(22) => 
                           ADDERPC_OUTs_22_port, NPC_OUT(21) => 
                           ADDERPC_OUTs_21_port, NPC_OUT(20) => 
                           ADDERPC_OUTs_20_port, NPC_OUT(19) => 
                           ADDERPC_OUTs_19_port, NPC_OUT(18) => 
                           ADDERPC_OUTs_18_port, NPC_OUT(17) => 
                           ADDERPC_OUTs_17_port, NPC_OUT(16) => 
                           ADDERPC_OUTs_16_port, NPC_OUT(15) => 
                           ADDERPC_OUTs_15_port, NPC_OUT(14) => 
                           ADDERPC_OUTs_14_port, NPC_OUT(13) => 
                           ADDERPC_OUTs_13_port, NPC_OUT(12) => 
                           ADDERPC_OUTs_12_port, NPC_OUT(11) => 
                           ADDERPC_OUTs_11_port, NPC_OUT(10) => 
                           ADDERPC_OUTs_10_port, NPC_OUT(9) => 
                           ADDERPC_OUTs_9_port, NPC_OUT(8) => 
                           ADDERPC_OUTs_8_port, NPC_OUT(7) => 
                           ADDERPC_OUTs_7_port, NPC_OUT(6) => 
                           ADDERPC_OUTs_6_port, NPC_OUT(5) => 
                           ADDERPC_OUTs_5_port, NPC_OUT(4) => 
                           ADDERPC_OUTs_4_port, NPC_OUT(3) => 
                           ADDERPC_OUTs_3_port, NPC_OUT(2) => 
                           ADDERPC_OUTs_2_port, NPC_OUT(1) => 
                           ADDERPC_OUTs_1_port, NPC_OUT(0) => 
                           ADDERPC_OUTs_0_port, COND_OUT => COND_OUTs, 
                           DRAM_DATAout(31) => LMD_OUTs_31_port, 
                           DRAM_DATAout(30) => LMD_OUTs_30_port, 
                           DRAM_DATAout(29) => LMD_OUTs_29_port, 
                           DRAM_DATAout(28) => LMD_OUTs_28_port, 
                           DRAM_DATAout(27) => LMD_OUTs_27_port, 
                           DRAM_DATAout(26) => LMD_OUTs_26_port, 
                           DRAM_DATAout(25) => LMD_OUTs_25_port, 
                           DRAM_DATAout(24) => LMD_OUTs_24_port, 
                           DRAM_DATAout(23) => LMD_OUTs_23_port, 
                           DRAM_DATAout(22) => LMD_OUTs_22_port, 
                           DRAM_DATAout(21) => LMD_OUTs_21_port, 
                           DRAM_DATAout(20) => LMD_OUTs_20_port, 
                           DRAM_DATAout(19) => LMD_OUTs_19_port, 
                           DRAM_DATAout(18) => LMD_OUTs_18_port, 
                           DRAM_DATAout(17) => LMD_OUTs_17_port, 
                           DRAM_DATAout(16) => LMD_OUTs_16_port, 
                           DRAM_DATAout(15) => LMD_OUTs_15_port, 
                           DRAM_DATAout(14) => LMD_OUTs_14_port, 
                           DRAM_DATAout(13) => LMD_OUTs_13_port, 
                           DRAM_DATAout(12) => LMD_OUTs_12_port, 
                           DRAM_DATAout(11) => LMD_OUTs_11_port, 
                           DRAM_DATAout(10) => LMD_OUTs_10_port, 
                           DRAM_DATAout(9) => LMD_OUTs_9_port, DRAM_DATAout(8) 
                           => LMD_OUTs_8_port, DRAM_DATAout(7) => 
                           LMD_OUTs_7_port, DRAM_DATAout(6) => LMD_OUTs_6_port,
                           DRAM_DATAout(5) => LMD_OUTs_5_port, DRAM_DATAout(4) 
                           => LMD_OUTs_4_port, DRAM_DATAout(3) => 
                           LMD_OUTs_3_port, DRAM_DATAout(2) => LMD_OUTs_2_port,
                           DRAM_DATAout(1) => LMD_OUTs_1_port, DRAM_DATAout(0) 
                           => LMD_OUTs_0_port, TO_PC_OUT(31) => 
                           TO_PC_OUTs_31_port, TO_PC_OUT(30) => 
                           TO_PC_OUTs_30_port, TO_PC_OUT(29) => 
                           TO_PC_OUTs_29_port, TO_PC_OUT(28) => 
                           TO_PC_OUTs_28_port, TO_PC_OUT(27) => 
                           TO_PC_OUTs_27_port, TO_PC_OUT(26) => 
                           TO_PC_OUTs_26_port, TO_PC_OUT(25) => 
                           TO_PC_OUTs_25_port, TO_PC_OUT(24) => 
                           TO_PC_OUTs_24_port, TO_PC_OUT(23) => 
                           TO_PC_OUTs_23_port, TO_PC_OUT(22) => 
                           TO_PC_OUTs_22_port, TO_PC_OUT(21) => 
                           TO_PC_OUTs_21_port, TO_PC_OUT(20) => 
                           TO_PC_OUTs_20_port, TO_PC_OUT(19) => 
                           TO_PC_OUTs_19_port, TO_PC_OUT(18) => 
                           TO_PC_OUTs_18_port, TO_PC_OUT(17) => 
                           TO_PC_OUTs_17_port, TO_PC_OUT(16) => 
                           TO_PC_OUTs_16_port, TO_PC_OUT(15) => 
                           TO_PC_OUTs_15_port, TO_PC_OUT(14) => 
                           TO_PC_OUTs_14_port, TO_PC_OUT(13) => 
                           TO_PC_OUTs_13_port, TO_PC_OUT(12) => 
                           TO_PC_OUTs_12_port, TO_PC_OUT(11) => 
                           TO_PC_OUTs_11_port, TO_PC_OUT(10) => 
                           TO_PC_OUTs_10_port, TO_PC_OUT(9) => 
                           TO_PC_OUTs_9_port, TO_PC_OUT(8) => TO_PC_OUTs_8_port
                           , TO_PC_OUT(7) => TO_PC_OUTs_7_port, TO_PC_OUT(6) =>
                           TO_PC_OUTs_6_port, TO_PC_OUT(5) => TO_PC_OUTs_5_port
                           , TO_PC_OUT(4) => TO_PC_OUTs_4_port, TO_PC_OUT(3) =>
                           TO_PC_OUTs_3_port, TO_PC_OUT(2) => TO_PC_OUTs_2_port
                           , TO_PC_OUT(1) => TO_PC_OUTs_1_port, TO_PC_OUT(0) =>
                           TO_PC_OUTs_0_port, ALU_OUT2(31) => ALU_OUT2s_31_port
                           , ALU_OUT2(30) => ALU_OUT2s_30_port, ALU_OUT2(29) =>
                           ALU_OUT2s_29_port, ALU_OUT2(28) => ALU_OUT2s_28_port
                           , ALU_OUT2(27) => ALU_OUT2s_27_port, ALU_OUT2(26) =>
                           ALU_OUT2s_26_port, ALU_OUT2(25) => ALU_OUT2s_25_port
                           , ALU_OUT2(24) => ALU_OUT2s_24_port, ALU_OUT2(23) =>
                           ALU_OUT2s_23_port, ALU_OUT2(22) => ALU_OUT2s_22_port
                           , ALU_OUT2(21) => ALU_OUT2s_21_port, ALU_OUT2(20) =>
                           ALU_OUT2s_20_port, ALU_OUT2(19) => ALU_OUT2s_19_port
                           , ALU_OUT2(18) => ALU_OUT2s_18_port, ALU_OUT2(17) =>
                           ALU_OUT2s_17_port, ALU_OUT2(16) => ALU_OUT2s_16_port
                           , ALU_OUT2(15) => ALU_OUT2s_15_port, ALU_OUT2(14) =>
                           ALU_OUT2s_14_port, ALU_OUT2(13) => ALU_OUT2s_13_port
                           , ALU_OUT2(12) => ALU_OUT2s_12_port, ALU_OUT2(11) =>
                           ALU_OUT2s_11_port, ALU_OUT2(10) => ALU_OUT2s_10_port
                           , ALU_OUT2(9) => ALU_OUT2s_9_port, ALU_OUT2(8) => 
                           ALU_OUT2s_8_port, ALU_OUT2(7) => ALU_OUT2s_7_port, 
                           ALU_OUT2(6) => ALU_OUT2s_6_port, ALU_OUT2(5) => 
                           ALU_OUT2s_5_port, ALU_OUT2(4) => ALU_OUT2s_4_port, 
                           ALU_OUT2(3) => ALU_OUT2s_3_port, ALU_OUT2(2) => 
                           ALU_OUT2s_2_port, ALU_OUT2(1) => ALU_OUT2s_1_port, 
                           ALU_OUT2(0) => ALU_OUT2s_0_port, IR_IN4(31) => 
                           IR_OUT3s_31_port, IR_IN4(30) => IR_OUT3s_30_port, 
                           IR_IN4(29) => IR_OUT3s_29_port, IR_IN4(28) => 
                           IR_OUT3s_28_port, IR_IN4(27) => IR_OUT3s_27_port, 
                           IR_IN4(26) => IR_OUT3s_26_port, IR_IN4(25) => 
                           IR_OUT3s_25_port, IR_IN4(24) => IR_OUT3s_24_port, 
                           IR_IN4(23) => IR_OUT3s_23_port, IR_IN4(22) => 
                           IR_OUT3s_22_port, IR_IN4(21) => IR_OUT3s_21_port, 
                           IR_IN4(20) => IR_OUT3s_20_port, IR_IN4(19) => 
                           IR_OUT3s_19_port, IR_IN4(18) => IR_OUT3s_18_port, 
                           IR_IN4(17) => IR_OUT3s_17_port, IR_IN4(16) => 
                           IR_OUT3s_16_port, IR_IN4(15) => IR_OUT3s_15_port, 
                           IR_IN4(14) => IR_OUT3s_14_port, IR_IN4(13) => 
                           IR_OUT3s_13_port, IR_IN4(12) => IR_OUT3s_12_port, 
                           IR_IN4(11) => IR_OUT3s_11_port, IR_IN4(10) => 
                           IR_OUT3s_10_port, IR_IN4(9) => IR_OUT3s_9_port, 
                           IR_IN4(8) => IR_OUT3s_8_port, IR_IN4(7) => 
                           IR_OUT3s_7_port, IR_IN4(6) => IR_OUT3s_6_port, 
                           IR_IN4(5) => IR_OUT3s_5_port, IR_IN4(4) => 
                           IR_OUT3s_4_port, IR_IN4(3) => IR_OUT3s_3_port, 
                           IR_IN4(2) => IR_OUT3s_2_port, IR_IN4(1) => 
                           IR_OUT3s_1_port, IR_IN4(0) => IR_OUT3s_0_port, 
                           IR_OUT4(31) => IR_OUT4s_31_port, IR_OUT4(30) => 
                           IR_OUT4s_30_port, IR_OUT4(29) => IR_OUT4s_29_port, 
                           IR_OUT4(28) => IR_OUT4s_28_port, IR_OUT4(27) => 
                           IR_OUT4s_27_port, IR_OUT4(26) => IR_OUT4s_26_port, 
                           IR_OUT4(25) => IR_OUT4s_25_port, IR_OUT4(24) => 
                           IR_OUT4s_24_port, IR_OUT4(23) => IR_OUT4s_23_port, 
                           IR_OUT4(22) => IR_OUT4s_22_port, IR_OUT4(21) => 
                           IR_OUT4s_21_port, IR_OUT4(20) => IR_OUT4s_20_port, 
                           IR_OUT4(19) => IR_OUT4s_19_port, IR_OUT4(18) => 
                           IR_OUT4s_18_port, IR_OUT4(17) => IR_OUT4s_17_port, 
                           IR_OUT4(16) => IR_OUT4s_16_port, IR_OUT4(15) => 
                           IR_OUT4s_15_port, IR_OUT4(14) => IR_OUT4s_14_port, 
                           IR_OUT4(13) => IR_OUT4s_13_port, IR_OUT4(12) => 
                           IR_OUT4s_12_port, IR_OUT4(11) => IR_OUT4s_11_port, 
                           IR_OUT4(10) => IR_OUT4s_10_port, IR_OUT4(9) => 
                           IR_OUT4s_9_port, IR_OUT4(8) => IR_OUT4s_8_port, 
                           IR_OUT4(7) => IR_OUT4s_7_port, IR_OUT4(6) => 
                           IR_OUT4s_6_port, IR_OUT4(5) => IR_OUT4s_5_port, 
                           IR_OUT4(4) => IR_OUT4s_4_port, IR_OUT4(3) => 
                           IR_OUT4s_3_port, IR_OUT4(2) => IR_OUT4s_2_port, 
                           IR_OUT4(1) => IR_OUT4s_1_port, IR_OUT4(0) => 
                           IR_OUT4s_0_port);
   WB : writeBack_nbits32 port map( LMD_OUT(31) => LMD_OUTs_31_port, 
                           LMD_OUT(30) => LMD_OUTs_30_port, LMD_OUT(29) => 
                           LMD_OUTs_29_port, LMD_OUT(28) => LMD_OUTs_28_port, 
                           LMD_OUT(27) => LMD_OUTs_27_port, LMD_OUT(26) => 
                           LMD_OUTs_26_port, LMD_OUT(25) => LMD_OUTs_25_port, 
                           LMD_OUT(24) => LMD_OUTs_24_port, LMD_OUT(23) => 
                           LMD_OUTs_23_port, LMD_OUT(22) => LMD_OUTs_22_port, 
                           LMD_OUT(21) => LMD_OUTs_21_port, LMD_OUT(20) => 
                           LMD_OUTs_20_port, LMD_OUT(19) => LMD_OUTs_19_port, 
                           LMD_OUT(18) => LMD_OUTs_18_port, LMD_OUT(17) => 
                           LMD_OUTs_17_port, LMD_OUT(16) => LMD_OUTs_16_port, 
                           LMD_OUT(15) => LMD_OUTs_15_port, LMD_OUT(14) => 
                           LMD_OUTs_14_port, LMD_OUT(13) => LMD_OUTs_13_port, 
                           LMD_OUT(12) => LMD_OUTs_12_port, LMD_OUT(11) => 
                           LMD_OUTs_11_port, LMD_OUT(10) => LMD_OUTs_10_port, 
                           LMD_OUT(9) => LMD_OUTs_9_port, LMD_OUT(8) => 
                           LMD_OUTs_8_port, LMD_OUT(7) => LMD_OUTs_7_port, 
                           LMD_OUT(6) => LMD_OUTs_6_port, LMD_OUT(5) => 
                           LMD_OUTs_5_port, LMD_OUT(4) => LMD_OUTs_4_port, 
                           LMD_OUT(3) => LMD_OUTs_3_port, LMD_OUT(2) => 
                           LMD_OUTs_2_port, LMD_OUT(1) => LMD_OUTs_1_port, 
                           LMD_OUT(0) => LMD_OUTs_0_port, ALUREG_OUTPUT(31) => 
                           ALU_OUT2s_31_port, ALUREG_OUTPUT(30) => 
                           ALU_OUT2s_30_port, ALUREG_OUTPUT(29) => 
                           ALU_OUT2s_29_port, ALUREG_OUTPUT(28) => 
                           ALU_OUT2s_28_port, ALUREG_OUTPUT(27) => 
                           ALU_OUT2s_27_port, ALUREG_OUTPUT(26) => 
                           ALU_OUT2s_26_port, ALUREG_OUTPUT(25) => 
                           ALU_OUT2s_25_port, ALUREG_OUTPUT(24) => 
                           ALU_OUT2s_24_port, ALUREG_OUTPUT(23) => 
                           ALU_OUT2s_23_port, ALUREG_OUTPUT(22) => 
                           ALU_OUT2s_22_port, ALUREG_OUTPUT(21) => 
                           ALU_OUT2s_21_port, ALUREG_OUTPUT(20) => 
                           ALU_OUT2s_20_port, ALUREG_OUTPUT(19) => 
                           ALU_OUT2s_19_port, ALUREG_OUTPUT(18) => 
                           ALU_OUT2s_18_port, ALUREG_OUTPUT(17) => 
                           ALU_OUT2s_17_port, ALUREG_OUTPUT(16) => 
                           ALU_OUT2s_16_port, ALUREG_OUTPUT(15) => 
                           ALU_OUT2s_15_port, ALUREG_OUTPUT(14) => 
                           ALU_OUT2s_14_port, ALUREG_OUTPUT(13) => 
                           ALU_OUT2s_13_port, ALUREG_OUTPUT(12) => 
                           ALU_OUT2s_12_port, ALUREG_OUTPUT(11) => 
                           ALU_OUT2s_11_port, ALUREG_OUTPUT(10) => 
                           ALU_OUT2s_10_port, ALUREG_OUTPUT(9) => 
                           ALU_OUT2s_9_port, ALUREG_OUTPUT(8) => 
                           ALU_OUT2s_8_port, ALUREG_OUTPUT(7) => 
                           ALU_OUT2s_7_port, ALUREG_OUTPUT(6) => 
                           ALU_OUT2s_6_port, ALUREG_OUTPUT(5) => 
                           ALU_OUT2s_5_port, ALUREG_OUTPUT(4) => 
                           ALU_OUT2s_4_port, ALUREG_OUTPUT(3) => 
                           ALU_OUT2s_3_port, ALUREG_OUTPUT(2) => 
                           ALU_OUT2s_2_port, ALUREG_OUTPUT(1) => 
                           ALU_OUT2s_1_port, ALUREG_OUTPUT(0) => 
                           ALU_OUT2s_0_port, WB_MUX_SEL => WB_MUX_SEL, 
                           DATAIN_RF(31) => DATAIN_RFs_31_port, DATAIN_RF(30) 
                           => DATAIN_RFs_30_port, DATAIN_RF(29) => 
                           DATAIN_RFs_29_port, DATAIN_RF(28) => 
                           DATAIN_RFs_28_port, DATAIN_RF(27) => 
                           DATAIN_RFs_27_port, DATAIN_RF(26) => 
                           DATAIN_RFs_26_port, DATAIN_RF(25) => 
                           DATAIN_RFs_25_port, DATAIN_RF(24) => 
                           DATAIN_RFs_24_port, DATAIN_RF(23) => 
                           DATAIN_RFs_23_port, DATAIN_RF(22) => 
                           DATAIN_RFs_22_port, DATAIN_RF(21) => 
                           DATAIN_RFs_21_port, DATAIN_RF(20) => 
                           DATAIN_RFs_20_port, DATAIN_RF(19) => 
                           DATAIN_RFs_19_port, DATAIN_RF(18) => 
                           DATAIN_RFs_18_port, DATAIN_RF(17) => 
                           DATAIN_RFs_17_port, DATAIN_RF(16) => 
                           DATAIN_RFs_16_port, DATAIN_RF(15) => 
                           DATAIN_RFs_15_port, DATAIN_RF(14) => 
                           DATAIN_RFs_14_port, DATAIN_RF(13) => 
                           DATAIN_RFs_13_port, DATAIN_RF(12) => 
                           DATAIN_RFs_12_port, DATAIN_RF(11) => 
                           DATAIN_RFs_11_port, DATAIN_RF(10) => 
                           DATAIN_RFs_10_port, DATAIN_RF(9) => 
                           DATAIN_RFs_9_port, DATAIN_RF(8) => DATAIN_RFs_8_port
                           , DATAIN_RF(7) => DATAIN_RFs_7_port, DATAIN_RF(6) =>
                           DATAIN_RFs_6_port, DATAIN_RF(5) => DATAIN_RFs_5_port
                           , DATAIN_RF(4) => DATAIN_RFs_4_port, DATAIN_RF(3) =>
                           DATAIN_RFs_3_port, DATAIN_RF(2) => DATAIN_RFs_2_port
                           , DATAIN_RF(1) => DATAIN_RFs_1_port, DATAIN_RF(0) =>
                           DATAIN_RFs_0_port);
   U1 : BUF_X1 port map( A => rst, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
         std_logic;  ALU_OPCODE : out std_logic_vector (0 to 3);  DRAM_WE, 
         LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, WB_MUX_SEL, RF_WE : out std_logic
         );

end dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, cw_8_port, cw_7_port, cw_1, cw1_5_port, cw1_4_port, 
      cw1_3_port, cw1_1, cw1_0, cw2_1_port, cw2_0_port, aluOpcode_i_3_port, 
      aluOpcode_i_2_port, aluOpcode_i_1_port, aluOpcode_i_0_port, n2, n105, 
      n106, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      RegA_LATCH_EN_port, n98, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n_1756, n_1757, n_1758, n_1759, 
      n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, 
      n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775 : std_logic;

begin
   IR_LATCH_EN <= X_Logic1_port;
   NPC_LATCH_EN <= X_Logic1_port;
   RegA_LATCH_EN <= RegA_LATCH_EN_port;
   RegIMM_LATCH_EN <= cw_8_port;
   PC_LATCH_EN <= X_Logic1_port;
   
   X_Logic1_port <= '1';
   cw1_reg_7_inst : DFFR_X1 port map( D => cw_7_port, CK => Clk, RN => n107, Q 
                           => ALU_OUTREG_EN, QN => n_1756);
   cw1_reg_6_inst : DFFR_X1 port map( D => n98, CK => Clk, RN => n107, Q => 
                           EQ_COND, QN => n_1757);
   cw1_reg_5_inst : DFFR_X1 port map( D => n106, CK => Clk, RN => n107, Q => 
                           cw1_5_port, QN => n_1758);
   cw1_reg_4_inst : SDFFR_X1 port map( D => IR_IN(31), SI => n2, SE => n105, CK
                           => Clk, RN => n107, Q => cw1_4_port, QN => n_1759);
   cw1_reg_3_inst : DFFR_X1 port map( D => n116, CK => Clk, RN => n107, Q => 
                           cw1_3_port, QN => n_1760);
   cw1_reg_1_inst : DFFR_X1 port map( D => cw_1, CK => Clk, RN => n107, Q => 
                           cw1_1, QN => n_1761);
   cw1_reg_0_inst : DFFR_X1 port map( D => n110, CK => Clk, RN => n107, Q => 
                           cw1_0, QN => n_1762);
   cw2_reg_5_inst : DFFR_X1 port map( D => cw1_5_port, CK => Clk, RN => n107, Q
                           => DRAM_WE, QN => n_1763);
   cw2_reg_4_inst : DFFR_X1 port map( D => cw1_4_port, CK => Clk, RN => n107, Q
                           => LMD_LATCH_EN, QN => n_1764);
   cw2_reg_3_inst : DFFR_X1 port map( D => cw1_3_port, CK => Clk, RN => n107, Q
                           => JUMP_EN, QN => n_1765);
   cw2_reg_1_inst : DFFR_X1 port map( D => cw1_1, CK => Clk, RN => n107, Q => 
                           cw2_1_port, QN => n_1766);
   cw2_reg_0_inst : DFFR_X1 port map( D => cw1_0, CK => Clk, RN => n107, Q => 
                           cw2_0_port, QN => n_1767);
   cw3_reg_0_inst : DFFR_X1 port map( D => cw2_0_port, CK => Clk, RN => n107, Q
                           => RF_WE, QN => n_1768);
   aluOpcode1_reg_3_inst : DFFS_X1 port map( D => aluOpcode_i_3_port, CK => Clk
                           , SN => n107, Q => ALU_OPCODE(0), QN => n_1769);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => aluOpcode_i_2_port, CK => Clk
                           , RN => n107, Q => ALU_OPCODE(1), QN => n_1770);
   aluOpcode1_reg_1_inst : DFFS_X1 port map( D => aluOpcode_i_1_port, CK => Clk
                           , SN => n107, Q => ALU_OPCODE(2), QN => n_1771);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => aluOpcode_i_0_port, CK => Clk
                           , RN => n107, Q => ALU_OPCODE(3), QN => n_1772);
   n2 <= '0';
   U96 : NAND3_X1 port map( A1 => n27, A2 => n119, A3 => n28, ZN => 
                           RegA_LATCH_EN_port);
   U97 : NAND3_X1 port map( A1 => n29, A2 => n125, A3 => n30, ZN => cw_8_port);
   U98 : NAND3_X1 port map( A1 => n27, A2 => n119, A3 => n33, ZN => cw_7_port);
   U99 : NAND3_X1 port map( A1 => n43, A2 => IR_IN(30), A3 => n44, ZN => n36);
   U100 : NAND3_X1 port map( A1 => IR_IN(3), A2 => n124, A3 => IR_IN(2), ZN => 
                           n45);
   U101 : NAND3_X1 port map( A1 => n51, A2 => n118, A3 => n52, ZN => 
                           aluOpcode_i_2_port);
   U102 : NAND3_X1 port map( A1 => n55, A2 => n56, A3 => n124, ZN => n51);
   U103 : OAI33_X1 port map( A1 => n114, A2 => IR_IN(3), A3 => n57, B1 => n58, 
                           B2 => n109, B3 => n113, ZN => n56);
   U104 : XOR2_X1 port map( A => IR_IN(0), B => IR_IN(3), Z => n73);
   U105 : NAND3_X1 port map( A1 => n55, A2 => n79, A3 => n124, ZN => n78);
   U106 : OAI33_X1 port map( A1 => n113, A2 => n80, A3 => n109, B1 => n81, B2 
                           => IR_IN(3), B3 => IR_IN(0), ZN => n79);
   U107 : XOR2_X1 port map( A => IR_IN(5), B => IR_IN(2), Z => n82);
   U108 : NAND3_X1 port map( A1 => n43, A2 => n131, A3 => n44, ZN => n76);
   U109 : NAND3_X1 port map( A1 => n55, A2 => n80, A3 => n93, ZN => n91);
   cw1_reg_8_inst : DFFR_X1 port map( D => cw_8_port, CK => Clk, RN => n107, Q 
                           => MUXB_SEL, QN => n_1773);
   cw3_reg_1_inst : DFFR_X1 port map( D => cw2_1_port, CK => Clk, RN => n107, Q
                           => WB_MUX_SEL, QN => n_1774);
   cw1_reg_9_inst : DFFR_X1 port map( D => RegA_LATCH_EN_port, CK => Clk, RN =>
                           n107, Q => MUXA_SEL, QN => n_1775);
   U3 : BUF_X1 port map( A => Rst, Z => n108);
   U5 : INV_X1 port map( A => n60, ZN => n126);
   U6 : NAND2_X1 port map( A1 => n76, A2 => n28, ZN => n98);
   U7 : INV_X1 port map( A => n27, ZN => n110);
   U8 : INV_X1 port map( A => n33, ZN => n116);
   U9 : INV_X1 port map( A => n106, ZN => n119);
   U10 : INV_X1 port map( A => n35, ZN => n124);
   U11 : NOR3_X1 port map( A1 => n31, A2 => n98, A3 => n106, ZN => n30);
   U12 : INV_X1 port map( A => n32, ZN => n125);
   U13 : NOR4_X1 port map( A1 => n53, A2 => n75, A3 => n126, A4 => n83, ZN => 
                           n37);
   U14 : OR2_X1 port map( A1 => n48, A2 => n84, ZN => n83);
   U15 : NOR3_X1 port map( A1 => n128, A2 => n74, A3 => n131, ZN => n84);
   U16 : NOR3_X1 port map( A1 => n70, A2 => n49, A3 => n131, ZN => n85);
   U17 : NAND2_X1 port map( A1 => n85, A2 => n129, ZN => n60);
   U18 : INV_X1 port map( A => n43, ZN => n128);
   U19 : NOR3_X1 port map( A1 => n130, A2 => n105, A3 => n132, ZN => n106);
   U20 : NAND2_X1 port map( A1 => n65, A2 => n131, ZN => n105);
   U21 : NOR4_X1 port map( A1 => n123, A2 => n131, A3 => n129, A4 => n49, ZN =>
                           n42);
   U22 : NOR3_X1 port map( A1 => n54, A2 => n49, A3 => n70, ZN => n53);
   U23 : NOR3_X1 port map( A1 => n49, A2 => n74, A3 => n54, ZN => n41);
   U24 : NOR3_X1 port map( A1 => n54, A2 => n49, A3 => n123, ZN => n40);
   U25 : INV_X1 port map( A => n44, ZN => n123);
   U26 : NAND2_X1 port map( A1 => n77, A2 => n117, ZN => n28);
   U27 : INV_X1 port map( A => n74, ZN => n117);
   U28 : NOR2_X1 port map( A1 => n31, A2 => cw_1, ZN => n27);
   U29 : OAI21_X1 port map( B1 => n34, B2 => n35, A => n29, ZN => cw_1);
   U30 : NAND4_X1 port map( A1 => n60, A2 => n120, A3 => n61, A4 => n62, ZN => 
                           aluOpcode_i_1_port);
   U31 : INV_X1 port map( A => n31, ZN => n120);
   U32 : NOR3_X1 port map( A1 => n75, A2 => n106, A3 => n116, ZN => n61);
   U33 : NOR4_X1 port map( A1 => n41, A2 => n39, A3 => n63, A4 => n50, ZN => 
                           n62);
   U34 : NOR3_X1 port map( A1 => n47, A2 => n98, A3 => n32, ZN => n33);
   U35 : INV_X1 port map( A => n59, ZN => n113);
   U36 : NAND2_X1 port map( A1 => n77, A2 => n44, ZN => n35);
   U37 : INV_X1 port map( A => n41, ZN => n118);
   U38 : NOR3_X1 port map( A1 => n126, A2 => n53, A3 => n40, ZN => n52);
   U39 : NOR3_X1 port map( A1 => n32, A2 => n106, A3 => n47, ZN => n86);
   U40 : OAI211_X1 port map( C1 => n34, C2 => n35, A => n76, B => n86, ZN => 
                           RegB_LATCH_EN);
   U41 : INV_X1 port map( A => n108, ZN => n107);
   U42 : NAND2_X1 port map( A1 => IR_IN(29), A2 => n132, ZN => n49);
   U43 : INV_X1 port map( A => IR_IN(31), ZN => n132);
   U44 : AND2_X1 port map( A1 => n85, A2 => IR_IN(28), ZN => n48);
   U45 : AND4_X1 port map( A1 => n36, A2 => n122, A3 => n37, A4 => n38, ZN => 
                           n29);
   U46 : NOR3_X1 port map( A1 => n39, A2 => n40, A3 => n41, ZN => n38);
   U47 : INV_X1 port map( A => n42, ZN => n122);
   U48 : NAND2_X1 port map( A1 => IR_IN(26), A2 => n127, ZN => n70);
   U49 : INV_X1 port map( A => IR_IN(27), ZN => n127);
   U50 : NOR3_X1 port map( A1 => IR_IN(29), A2 => IR_IN(31), A3 => n129, ZN => 
                           n43);
   U51 : INV_X1 port map( A => IR_IN(28), ZN => n129);
   U52 : INV_X1 port map( A => IR_IN(30), ZN => n131);
   U53 : NAND2_X1 port map( A1 => IR_IN(27), A2 => n121, ZN => n74);
   U54 : INV_X1 port map( A => IR_IN(26), ZN => n121);
   U55 : NOR3_X1 port map( A1 => n70, A2 => IR_IN(30), A3 => n128, ZN => n32);
   U56 : NOR3_X1 port map( A1 => n121, A2 => IR_IN(28), A3 => n127, ZN => n65);
   U57 : NOR4_X1 port map( A1 => n49, A2 => n74, A3 => IR_IN(28), A4 => 
                           IR_IN(30), ZN => n75);
   U58 : NAND2_X1 port map( A1 => IR_IN(28), A2 => n131, ZN => n54);
   U59 : NOR4_X1 port map( A1 => n123, A2 => n49, A3 => IR_IN(28), A4 => 
                           IR_IN(30), ZN => n39);
   U60 : NOR3_X1 port map( A1 => n105, A2 => IR_IN(29), A3 => n132, ZN => n31);
   U61 : NOR2_X1 port map( A1 => IR_IN(26), A2 => IR_IN(27), ZN => n44);
   U62 : NOR4_X1 port map( A1 => IR_IN(28), A2 => IR_IN(29), A3 => IR_IN(30), 
                           A4 => IR_IN(31), ZN => n77);
   U63 : INV_X1 port map( A => IR_IN(29), ZN => n130);
   U64 : OAI221_X1 port map( B1 => n64, B2 => n35, C1 => n65, C2 => n132, A => 
                           n66, ZN => n50);
   U65 : AND3_X1 port map( A1 => n55, A2 => n71, A3 => n72, ZN => n64);
   U66 : AOI221_X1 port map( B1 => IR_IN(30), B2 => n67, C1 => IR_IN(27), C2 =>
                           n68, A => n69, ZN => n66);
   U67 : OAI21_X1 port map( B1 => n73, B2 => n115, A => n114, ZN => n72);
   U68 : OAI22_X1 port map( A1 => n121, A2 => n49, B1 => IR_IN(29), B2 => n54, 
                           ZN => n68);
   U69 : NOR4_X1 port map( A1 => IR_IN(6), A2 => IR_IN(4), A3 => IR_IN(10), A4 
                           => n94, ZN => n55);
   U70 : OR3_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), ZN =>
                           n94);
   U71 : NOR4_X1 port map( A1 => n91, A2 => n92, A3 => IR_IN(14), A4 => 
                           IR_IN(13), ZN => n90);
   U72 : OR3_X1 port map( A1 => IR_IN(17), A2 => IR_IN(16), A3 => IR_IN(15), ZN
                           => n92);
   U73 : NOR3_X1 port map( A1 => IR_IN(0), A2 => IR_IN(12), A3 => IR_IN(11), ZN
                           => n93);
   U74 : AND4_X1 port map( A1 => n87, A2 => n88, A3 => n89, A4 => n90, ZN => 
                           n34);
   U75 : NOR2_X1 port map( A1 => IR_IN(19), A2 => IR_IN(18), ZN => n87);
   U76 : NOR3_X1 port map( A1 => IR_IN(1), A2 => IR_IN(21), A3 => IR_IN(20), ZN
                           => n88);
   U77 : NOR4_X1 port map( A1 => n95, A2 => IR_IN(24), A3 => IR_IN(5), A4 => 
                           IR_IN(25), ZN => n89);
   U78 : NOR3_X1 port map( A1 => n70, A2 => IR_IN(30), A3 => IR_IN(28), ZN => 
                           n69);
   U79 : NOR2_X1 port map( A1 => n115, A2 => IR_IN(1), ZN => n59);
   U80 : OAI21_X1 port map( B1 => IR_IN(3), B2 => IR_IN(0), A => n113, ZN => 
                           n71);
   U81 : INV_X1 port map( A => IR_IN(5), ZN => n115);
   U82 : OAI222_X1 port map( A1 => IR_IN(29), A2 => n121, B1 => IR_IN(28), B2 
                           => IR_IN(26), C1 => n127, C2 => n130, ZN => n67);
   U83 : NAND4_X1 port map( A1 => n45, A2 => n28, A3 => n111, A4 => n46, ZN => 
                           aluOpcode_i_3_port);
   U84 : NOR3_X1 port map( A1 => n42, A2 => n47, A3 => n48, ZN => n46);
   U85 : INV_X1 port map( A => n50, ZN => n111);
   U86 : NOR3_X1 port map( A1 => IR_IN(29), A2 => IR_IN(31), A3 => n105, ZN => 
                           n47);
   U87 : NAND2_X1 port map( A1 => n37, A2 => n78, ZN => aluOpcode_i_0_port);
   U88 : NAND2_X1 port map( A1 => IR_IN(1), A2 => n82, ZN => n81);
   U89 : INV_X1 port map( A => IR_IN(2), ZN => n114);
   U90 : NOR2_X1 port map( A1 => IR_IN(3), A2 => IR_IN(2), ZN => n80);
   U91 : AOI211_X1 port map( C1 => IR_IN(2), C2 => n112, A => n115, B => n35, 
                           ZN => n63);
   U92 : INV_X1 port map( A => IR_IN(1), ZN => n112);
   U93 : OR2_X1 port map( A1 => IR_IN(23), A2 => IR_IN(22), ZN => n95);
   U94 : NAND2_X1 port map( A1 => IR_IN(3), A2 => n114, ZN => n58);
   U95 : AOI21_X1 port map( B1 => IR_IN(5), B2 => n109, A => n59, ZN => n57);
   U110 : INV_X1 port map( A => IR_IN(0), ZN => n109);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity dlx is

   port( Clk_port, Rst_port : in std_logic;  DATA_IRAM_port, DATAread_DRAM_port
         : in std_logic_vector (31 downto 0);  WE_DRAM_port : out std_logic;  
         ADDRESS_DRAM_port, DATAwrite_DRAM_port, ADDRESS_IRAM_port : out 
         std_logic_vector (31 downto 0));

end dlx;

architecture SYN_STRUCTURAL of dlx is

   component datapath_nbits32
      port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 
            downto 0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN, RegA_LATCH_EN, 
            RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE, MUXA_SEL, MUXB_SEL, 
            ALU_OUTREG_EN, EQ_COND : in std_logic;  ALU_OPCODE : in 
            std_logic_vector (0 to 3);  DRAM_DATA : in std_logic_vector (31 
            downto 0);  LMD_LATCH_EN, JUMP_EN, WB_MUX_SEL : in std_logic;  B, 
            ALU_OUT, ADDRESS_IRAM, IR_OUT : out std_logic_vector (31 downto 0)
            );
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
            std_logic;  ALU_OPCODE : out std_logic_vector (0 to 3);  DRAM_WE, 
            LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, WB_MUX_SEL, RF_WE : out 
            std_logic);
   end component;
   
   signal IR_OUT_signal_31_port, IR_OUT_signal_30_port, IR_OUT_signal_29_port, 
      IR_OUT_signal_28_port, IR_OUT_signal_27_port, IR_OUT_signal_26_port, 
      IR_OUT_signal_25_port, IR_OUT_signal_24_port, IR_OUT_signal_23_port, 
      IR_OUT_signal_22_port, IR_OUT_signal_21_port, IR_OUT_signal_20_port, 
      IR_OUT_signal_19_port, IR_OUT_signal_18_port, IR_OUT_signal_17_port, 
      IR_OUT_signal_16_port, IR_OUT_signal_15_port, IR_OUT_signal_14_port, 
      IR_OUT_signal_13_port, IR_OUT_signal_12_port, IR_OUT_signal_11_port, 
      IR_OUT_signal_10_port, IR_OUT_signal_9_port, IR_OUT_signal_8_port, 
      IR_OUT_signal_7_port, IR_OUT_signal_6_port, IR_OUT_signal_5_port, 
      IR_OUT_signal_4_port, IR_OUT_signal_3_port, IR_OUT_signal_2_port, 
      IR_OUT_signal_1_port, IR_OUT_signal_0_port, IR_LATCH_EN_signal, 
      NPC_LATCH_EN_signal, RegA_LATCH_EN_signal, RegB_LATCH_EN_signal, 
      RegIMM_LATCH_EN_signal, MUXA_SEL_signal, MUXB_SEL_signal, 
      ALU_OUTREG_EN_signal, EQ_COND_signal, ALU_OPCODE_signal_0_port, 
      ALU_OPCODE_signal_1_port, ALU_OPCODE_signal_2_port, 
      ALU_OPCODE_signal_3_port, LMD_LATCH_EN_signal, JUMP_EN_signal, 
      PC_LATCH_EN_signal, WB_MUX_SEL_signal, RF_WE_signal, n_1776, n_1777, 
      n_1778 : std_logic;

begin
   
   PC_LATCH_EN_signal <= '1';
   NPC_LATCH_EN_signal <= '1';
   IR_LATCH_EN_signal <= '1';
   CONTROL_UNIT : 
                           dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 
                           port map( Clk => Clk_port, Rst => Rst_port, 
                           IR_IN(31) => IR_OUT_signal_31_port, IR_IN(30) => 
                           IR_OUT_signal_30_port, IR_IN(29) => 
                           IR_OUT_signal_29_port, IR_IN(28) => 
                           IR_OUT_signal_28_port, IR_IN(27) => 
                           IR_OUT_signal_27_port, IR_IN(26) => 
                           IR_OUT_signal_26_port, IR_IN(25) => 
                           IR_OUT_signal_25_port, IR_IN(24) => 
                           IR_OUT_signal_24_port, IR_IN(23) => 
                           IR_OUT_signal_23_port, IR_IN(22) => 
                           IR_OUT_signal_22_port, IR_IN(21) => 
                           IR_OUT_signal_21_port, IR_IN(20) => 
                           IR_OUT_signal_20_port, IR_IN(19) => 
                           IR_OUT_signal_19_port, IR_IN(18) => 
                           IR_OUT_signal_18_port, IR_IN(17) => 
                           IR_OUT_signal_17_port, IR_IN(16) => 
                           IR_OUT_signal_16_port, IR_IN(15) => 
                           IR_OUT_signal_15_port, IR_IN(14) => 
                           IR_OUT_signal_14_port, IR_IN(13) => 
                           IR_OUT_signal_13_port, IR_IN(12) => 
                           IR_OUT_signal_12_port, IR_IN(11) => 
                           IR_OUT_signal_11_port, IR_IN(10) => 
                           IR_OUT_signal_10_port, IR_IN(9) => 
                           IR_OUT_signal_9_port, IR_IN(8) => 
                           IR_OUT_signal_8_port, IR_IN(7) => 
                           IR_OUT_signal_7_port, IR_IN(6) => 
                           IR_OUT_signal_6_port, IR_IN(5) => 
                           IR_OUT_signal_5_port, IR_IN(4) => 
                           IR_OUT_signal_4_port, IR_IN(3) => 
                           IR_OUT_signal_3_port, IR_IN(2) => 
                           IR_OUT_signal_2_port, IR_IN(1) => 
                           IR_OUT_signal_1_port, IR_IN(0) => 
                           IR_OUT_signal_0_port, IR_LATCH_EN => n_1776, 
                           NPC_LATCH_EN => n_1777, RegA_LATCH_EN => 
                           RegA_LATCH_EN_signal, RegB_LATCH_EN => 
                           RegB_LATCH_EN_signal, RegIMM_LATCH_EN => 
                           RegIMM_LATCH_EN_signal, MUXA_SEL => MUXA_SEL_signal,
                           MUXB_SEL => MUXB_SEL_signal, ALU_OUTREG_EN => 
                           ALU_OUTREG_EN_signal, EQ_COND => EQ_COND_signal, 
                           ALU_OPCODE(0) => ALU_OPCODE_signal_0_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_signal_1_port, 
                           ALU_OPCODE(2) => ALU_OPCODE_signal_2_port, 
                           ALU_OPCODE(3) => ALU_OPCODE_signal_3_port, DRAM_WE 
                           => WE_DRAM_port, LMD_LATCH_EN => LMD_LATCH_EN_signal
                           , JUMP_EN => JUMP_EN_signal, PC_LATCH_EN => n_1778, 
                           WB_MUX_SEL => WB_MUX_SEL_signal, RF_WE => 
                           RF_WE_signal);
   DATA_PATH : datapath_nbits32 port map( clk => Clk_port, rst => Rst_port, 
                           DATA_IRAM(31) => DATA_IRAM_port(31), DATA_IRAM(30) 
                           => DATA_IRAM_port(30), DATA_IRAM(29) => 
                           DATA_IRAM_port(29), DATA_IRAM(28) => 
                           DATA_IRAM_port(28), DATA_IRAM(27) => 
                           DATA_IRAM_port(27), DATA_IRAM(26) => 
                           DATA_IRAM_port(26), DATA_IRAM(25) => 
                           DATA_IRAM_port(25), DATA_IRAM(24) => 
                           DATA_IRAM_port(24), DATA_IRAM(23) => 
                           DATA_IRAM_port(23), DATA_IRAM(22) => 
                           DATA_IRAM_port(22), DATA_IRAM(21) => 
                           DATA_IRAM_port(21), DATA_IRAM(20) => 
                           DATA_IRAM_port(20), DATA_IRAM(19) => 
                           DATA_IRAM_port(19), DATA_IRAM(18) => 
                           DATA_IRAM_port(18), DATA_IRAM(17) => 
                           DATA_IRAM_port(17), DATA_IRAM(16) => 
                           DATA_IRAM_port(16), DATA_IRAM(15) => 
                           DATA_IRAM_port(15), DATA_IRAM(14) => 
                           DATA_IRAM_port(14), DATA_IRAM(13) => 
                           DATA_IRAM_port(13), DATA_IRAM(12) => 
                           DATA_IRAM_port(12), DATA_IRAM(11) => 
                           DATA_IRAM_port(11), DATA_IRAM(10) => 
                           DATA_IRAM_port(10), DATA_IRAM(9) => 
                           DATA_IRAM_port(9), DATA_IRAM(8) => DATA_IRAM_port(8)
                           , DATA_IRAM(7) => DATA_IRAM_port(7), DATA_IRAM(6) =>
                           DATA_IRAM_port(6), DATA_IRAM(5) => DATA_IRAM_port(5)
                           , DATA_IRAM(4) => DATA_IRAM_port(4), DATA_IRAM(3) =>
                           DATA_IRAM_port(3), DATA_IRAM(2) => DATA_IRAM_port(2)
                           , DATA_IRAM(1) => DATA_IRAM_port(1), DATA_IRAM(0) =>
                           DATA_IRAM_port(0), IR_LATCH_EN => IR_LATCH_EN_signal
                           , NPC_LATCH_EN => NPC_LATCH_EN_signal, PC_LATCH_EN 
                           => PC_LATCH_EN_signal, RegA_LATCH_EN => 
                           RegA_LATCH_EN_signal, RegB_LATCH_EN => 
                           RegB_LATCH_EN_signal, RegIMM_LATCH_EN => 
                           RegIMM_LATCH_EN_signal, RF_WE => RF_WE_signal, 
                           MUXA_SEL => MUXA_SEL_signal, MUXB_SEL => 
                           MUXB_SEL_signal, ALU_OUTREG_EN => 
                           ALU_OUTREG_EN_signal, EQ_COND => EQ_COND_signal, 
                           ALU_OPCODE(0) => ALU_OPCODE_signal_0_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_signal_1_port, 
                           ALU_OPCODE(2) => ALU_OPCODE_signal_2_port, 
                           ALU_OPCODE(3) => ALU_OPCODE_signal_3_port, 
                           DRAM_DATA(31) => DATAread_DRAM_port(31), 
                           DRAM_DATA(30) => DATAread_DRAM_port(30), 
                           DRAM_DATA(29) => DATAread_DRAM_port(29), 
                           DRAM_DATA(28) => DATAread_DRAM_port(28), 
                           DRAM_DATA(27) => DATAread_DRAM_port(27), 
                           DRAM_DATA(26) => DATAread_DRAM_port(26), 
                           DRAM_DATA(25) => DATAread_DRAM_port(25), 
                           DRAM_DATA(24) => DATAread_DRAM_port(24), 
                           DRAM_DATA(23) => DATAread_DRAM_port(23), 
                           DRAM_DATA(22) => DATAread_DRAM_port(22), 
                           DRAM_DATA(21) => DATAread_DRAM_port(21), 
                           DRAM_DATA(20) => DATAread_DRAM_port(20), 
                           DRAM_DATA(19) => DATAread_DRAM_port(19), 
                           DRAM_DATA(18) => DATAread_DRAM_port(18), 
                           DRAM_DATA(17) => DATAread_DRAM_port(17), 
                           DRAM_DATA(16) => DATAread_DRAM_port(16), 
                           DRAM_DATA(15) => DATAread_DRAM_port(15), 
                           DRAM_DATA(14) => DATAread_DRAM_port(14), 
                           DRAM_DATA(13) => DATAread_DRAM_port(13), 
                           DRAM_DATA(12) => DATAread_DRAM_port(12), 
                           DRAM_DATA(11) => DATAread_DRAM_port(11), 
                           DRAM_DATA(10) => DATAread_DRAM_port(10), 
                           DRAM_DATA(9) => DATAread_DRAM_port(9), DRAM_DATA(8) 
                           => DATAread_DRAM_port(8), DRAM_DATA(7) => 
                           DATAread_DRAM_port(7), DRAM_DATA(6) => 
                           DATAread_DRAM_port(6), DRAM_DATA(5) => 
                           DATAread_DRAM_port(5), DRAM_DATA(4) => 
                           DATAread_DRAM_port(4), DRAM_DATA(3) => 
                           DATAread_DRAM_port(3), DRAM_DATA(2) => 
                           DATAread_DRAM_port(2), DRAM_DATA(1) => 
                           DATAread_DRAM_port(1), DRAM_DATA(0) => 
                           DATAread_DRAM_port(0), LMD_LATCH_EN => 
                           LMD_LATCH_EN_signal, JUMP_EN => JUMP_EN_signal, 
                           WB_MUX_SEL => WB_MUX_SEL_signal, B(31) => 
                           DATAwrite_DRAM_port(31), B(30) => 
                           DATAwrite_DRAM_port(30), B(29) => 
                           DATAwrite_DRAM_port(29), B(28) => 
                           DATAwrite_DRAM_port(28), B(27) => 
                           DATAwrite_DRAM_port(27), B(26) => 
                           DATAwrite_DRAM_port(26), B(25) => 
                           DATAwrite_DRAM_port(25), B(24) => 
                           DATAwrite_DRAM_port(24), B(23) => 
                           DATAwrite_DRAM_port(23), B(22) => 
                           DATAwrite_DRAM_port(22), B(21) => 
                           DATAwrite_DRAM_port(21), B(20) => 
                           DATAwrite_DRAM_port(20), B(19) => 
                           DATAwrite_DRAM_port(19), B(18) => 
                           DATAwrite_DRAM_port(18), B(17) => 
                           DATAwrite_DRAM_port(17), B(16) => 
                           DATAwrite_DRAM_port(16), B(15) => 
                           DATAwrite_DRAM_port(15), B(14) => 
                           DATAwrite_DRAM_port(14), B(13) => 
                           DATAwrite_DRAM_port(13), B(12) => 
                           DATAwrite_DRAM_port(12), B(11) => 
                           DATAwrite_DRAM_port(11), B(10) => 
                           DATAwrite_DRAM_port(10), B(9) => 
                           DATAwrite_DRAM_port(9), B(8) => 
                           DATAwrite_DRAM_port(8), B(7) => 
                           DATAwrite_DRAM_port(7), B(6) => 
                           DATAwrite_DRAM_port(6), B(5) => 
                           DATAwrite_DRAM_port(5), B(4) => 
                           DATAwrite_DRAM_port(4), B(3) => 
                           DATAwrite_DRAM_port(3), B(2) => 
                           DATAwrite_DRAM_port(2), B(1) => 
                           DATAwrite_DRAM_port(1), B(0) => 
                           DATAwrite_DRAM_port(0), ALU_OUT(31) => 
                           ADDRESS_DRAM_port(31), ALU_OUT(30) => 
                           ADDRESS_DRAM_port(30), ALU_OUT(29) => 
                           ADDRESS_DRAM_port(29), ALU_OUT(28) => 
                           ADDRESS_DRAM_port(28), ALU_OUT(27) => 
                           ADDRESS_DRAM_port(27), ALU_OUT(26) => 
                           ADDRESS_DRAM_port(26), ALU_OUT(25) => 
                           ADDRESS_DRAM_port(25), ALU_OUT(24) => 
                           ADDRESS_DRAM_port(24), ALU_OUT(23) => 
                           ADDRESS_DRAM_port(23), ALU_OUT(22) => 
                           ADDRESS_DRAM_port(22), ALU_OUT(21) => 
                           ADDRESS_DRAM_port(21), ALU_OUT(20) => 
                           ADDRESS_DRAM_port(20), ALU_OUT(19) => 
                           ADDRESS_DRAM_port(19), ALU_OUT(18) => 
                           ADDRESS_DRAM_port(18), ALU_OUT(17) => 
                           ADDRESS_DRAM_port(17), ALU_OUT(16) => 
                           ADDRESS_DRAM_port(16), ALU_OUT(15) => 
                           ADDRESS_DRAM_port(15), ALU_OUT(14) => 
                           ADDRESS_DRAM_port(14), ALU_OUT(13) => 
                           ADDRESS_DRAM_port(13), ALU_OUT(12) => 
                           ADDRESS_DRAM_port(12), ALU_OUT(11) => 
                           ADDRESS_DRAM_port(11), ALU_OUT(10) => 
                           ADDRESS_DRAM_port(10), ALU_OUT(9) => 
                           ADDRESS_DRAM_port(9), ALU_OUT(8) => 
                           ADDRESS_DRAM_port(8), ALU_OUT(7) => 
                           ADDRESS_DRAM_port(7), ALU_OUT(6) => 
                           ADDRESS_DRAM_port(6), ALU_OUT(5) => 
                           ADDRESS_DRAM_port(5), ALU_OUT(4) => 
                           ADDRESS_DRAM_port(4), ALU_OUT(3) => 
                           ADDRESS_DRAM_port(3), ALU_OUT(2) => 
                           ADDRESS_DRAM_port(2), ALU_OUT(1) => 
                           ADDRESS_DRAM_port(1), ALU_OUT(0) => 
                           ADDRESS_DRAM_port(0), ADDRESS_IRAM(31) => 
                           ADDRESS_IRAM_port(31), ADDRESS_IRAM(30) => 
                           ADDRESS_IRAM_port(30), ADDRESS_IRAM(29) => 
                           ADDRESS_IRAM_port(29), ADDRESS_IRAM(28) => 
                           ADDRESS_IRAM_port(28), ADDRESS_IRAM(27) => 
                           ADDRESS_IRAM_port(27), ADDRESS_IRAM(26) => 
                           ADDRESS_IRAM_port(26), ADDRESS_IRAM(25) => 
                           ADDRESS_IRAM_port(25), ADDRESS_IRAM(24) => 
                           ADDRESS_IRAM_port(24), ADDRESS_IRAM(23) => 
                           ADDRESS_IRAM_port(23), ADDRESS_IRAM(22) => 
                           ADDRESS_IRAM_port(22), ADDRESS_IRAM(21) => 
                           ADDRESS_IRAM_port(21), ADDRESS_IRAM(20) => 
                           ADDRESS_IRAM_port(20), ADDRESS_IRAM(19) => 
                           ADDRESS_IRAM_port(19), ADDRESS_IRAM(18) => 
                           ADDRESS_IRAM_port(18), ADDRESS_IRAM(17) => 
                           ADDRESS_IRAM_port(17), ADDRESS_IRAM(16) => 
                           ADDRESS_IRAM_port(16), ADDRESS_IRAM(15) => 
                           ADDRESS_IRAM_port(15), ADDRESS_IRAM(14) => 
                           ADDRESS_IRAM_port(14), ADDRESS_IRAM(13) => 
                           ADDRESS_IRAM_port(13), ADDRESS_IRAM(12) => 
                           ADDRESS_IRAM_port(12), ADDRESS_IRAM(11) => 
                           ADDRESS_IRAM_port(11), ADDRESS_IRAM(10) => 
                           ADDRESS_IRAM_port(10), ADDRESS_IRAM(9) => 
                           ADDRESS_IRAM_port(9), ADDRESS_IRAM(8) => 
                           ADDRESS_IRAM_port(8), ADDRESS_IRAM(7) => 
                           ADDRESS_IRAM_port(7), ADDRESS_IRAM(6) => 
                           ADDRESS_IRAM_port(6), ADDRESS_IRAM(5) => 
                           ADDRESS_IRAM_port(5), ADDRESS_IRAM(4) => 
                           ADDRESS_IRAM_port(4), ADDRESS_IRAM(3) => 
                           ADDRESS_IRAM_port(3), ADDRESS_IRAM(2) => 
                           ADDRESS_IRAM_port(2), ADDRESS_IRAM(1) => 
                           ADDRESS_IRAM_port(1), ADDRESS_IRAM(0) => 
                           ADDRESS_IRAM_port(0), IR_OUT(31) => 
                           IR_OUT_signal_31_port, IR_OUT(30) => 
                           IR_OUT_signal_30_port, IR_OUT(29) => 
                           IR_OUT_signal_29_port, IR_OUT(28) => 
                           IR_OUT_signal_28_port, IR_OUT(27) => 
                           IR_OUT_signal_27_port, IR_OUT(26) => 
                           IR_OUT_signal_26_port, IR_OUT(25) => 
                           IR_OUT_signal_25_port, IR_OUT(24) => 
                           IR_OUT_signal_24_port, IR_OUT(23) => 
                           IR_OUT_signal_23_port, IR_OUT(22) => 
                           IR_OUT_signal_22_port, IR_OUT(21) => 
                           IR_OUT_signal_21_port, IR_OUT(20) => 
                           IR_OUT_signal_20_port, IR_OUT(19) => 
                           IR_OUT_signal_19_port, IR_OUT(18) => 
                           IR_OUT_signal_18_port, IR_OUT(17) => 
                           IR_OUT_signal_17_port, IR_OUT(16) => 
                           IR_OUT_signal_16_port, IR_OUT(15) => 
                           IR_OUT_signal_15_port, IR_OUT(14) => 
                           IR_OUT_signal_14_port, IR_OUT(13) => 
                           IR_OUT_signal_13_port, IR_OUT(12) => 
                           IR_OUT_signal_12_port, IR_OUT(11) => 
                           IR_OUT_signal_11_port, IR_OUT(10) => 
                           IR_OUT_signal_10_port, IR_OUT(9) => 
                           IR_OUT_signal_9_port, IR_OUT(8) => 
                           IR_OUT_signal_8_port, IR_OUT(7) => 
                           IR_OUT_signal_7_port, IR_OUT(6) => 
                           IR_OUT_signal_6_port, IR_OUT(5) => 
                           IR_OUT_signal_5_port, IR_OUT(4) => 
                           IR_OUT_signal_4_port, IR_OUT(3) => 
                           IR_OUT_signal_3_port, IR_OUT(2) => 
                           IR_OUT_signal_2_port, IR_OUT(1) => 
                           IR_OUT_signal_1_port, IR_OUT(0) => 
                           IR_OUT_signal_0_port);

end SYN_STRUCTURAL;
