
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_dlx is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (LLS, LRS, ADDS, SUBS, ANDS, ORS, XORS, SNES, SLES, SGES, NOP);
attribute ENUM_ENCODING of aluOp : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";

end CONV_PACK_dlx;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity logic_and_shift_N32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end logic_and_shift_N32_DW01_ash_0;

architecture SYN_mx2 of logic_and_shift_N32_DW01_ash_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal temp_int_SH_4_port, temp_int_SH_3_port, temp_int_SH_2_port, 
      temp_int_SH_1_port, temp_int_SH_0_port, SHMAG_5_port, ML_int_1_31_port, 
      ML_int_1_30_port, ML_int_1_29_port, ML_int_1_28_port, ML_int_1_27_port, 
      ML_int_1_26_port, ML_int_1_25_port, ML_int_1_24_port, ML_int_1_23_port, 
      ML_int_1_22_port, ML_int_1_21_port, ML_int_1_20_port, ML_int_1_19_port, 
      ML_int_1_18_port, ML_int_1_17_port, ML_int_1_16_port, ML_int_1_15_port, 
      ML_int_1_14_port, ML_int_1_13_port, ML_int_1_12_port, ML_int_1_11_port, 
      ML_int_1_10_port, ML_int_1_9_port, ML_int_1_8_port, ML_int_1_7_port, 
      ML_int_1_6_port, ML_int_1_5_port, ML_int_1_4_port, ML_int_1_3_port, 
      ML_int_1_2_port, ML_int_1_1_port, ML_int_1_0_port, ML_int_2_31_port, 
      ML_int_2_30_port, ML_int_2_29_port, ML_int_2_28_port, ML_int_2_27_port, 
      ML_int_2_26_port, ML_int_2_25_port, ML_int_2_24_port, ML_int_2_23_port, 
      ML_int_2_22_port, ML_int_2_21_port, ML_int_2_20_port, ML_int_2_19_port, 
      ML_int_2_18_port, ML_int_2_17_port, ML_int_2_16_port, ML_int_2_15_port, 
      ML_int_2_14_port, ML_int_2_13_port, ML_int_2_12_port, ML_int_2_11_port, 
      ML_int_2_10_port, ML_int_2_9_port, ML_int_2_8_port, ML_int_2_7_port, 
      ML_int_2_6_port, ML_int_2_5_port, ML_int_2_4_port, ML_int_2_3_port, 
      ML_int_2_2_port, ML_int_2_1_port, ML_int_2_0_port, ML_int_3_31_port, 
      ML_int_3_30_port, ML_int_3_29_port, ML_int_3_28_port, ML_int_3_27_port, 
      ML_int_3_26_port, ML_int_3_25_port, ML_int_3_24_port, ML_int_3_23_port, 
      ML_int_3_22_port, ML_int_3_21_port, ML_int_3_20_port, ML_int_3_19_port, 
      ML_int_3_18_port, ML_int_3_17_port, ML_int_3_16_port, ML_int_3_15_port, 
      ML_int_3_14_port, ML_int_3_13_port, ML_int_3_12_port, ML_int_3_11_port, 
      ML_int_3_10_port, ML_int_3_9_port, ML_int_3_8_port, ML_int_3_7_port, 
      ML_int_3_6_port, ML_int_3_5_port, ML_int_3_4_port, ML_int_3_3_port, 
      ML_int_3_2_port, ML_int_3_1_port, ML_int_3_0_port, ML_int_4_31_port, 
      ML_int_4_30_port, ML_int_4_29_port, ML_int_4_28_port, ML_int_4_27_port, 
      ML_int_4_26_port, ML_int_4_25_port, ML_int_4_24_port, ML_int_4_23_port, 
      ML_int_4_22_port, ML_int_4_21_port, ML_int_4_20_port, ML_int_4_19_port, 
      ML_int_4_18_port, ML_int_4_17_port, ML_int_4_16_port, ML_int_4_15_port, 
      ML_int_4_14_port, ML_int_4_13_port, ML_int_4_12_port, ML_int_4_11_port, 
      ML_int_4_10_port, ML_int_4_9_port, ML_int_4_8_port, ML_int_5_31_port, 
      ML_int_5_30_port, ML_int_5_29_port, ML_int_5_28_port, ML_int_5_27_port, 
      ML_int_5_26_port, ML_int_5_25_port, ML_int_5_24_port, ML_int_5_23_port, 
      ML_int_5_22_port, ML_int_5_21_port, ML_int_5_20_port, ML_int_5_19_port, 
      ML_int_5_18_port, ML_int_5_17_port, ML_int_5_16_port, n1, n2, n3, n4, n5,
      n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, 
      n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63 : 
      std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_31_port);
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_30_port);
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_29_port);
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_28_port);
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_27_port);
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_26_port);
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_25_port);
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_24_port);
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => n8, S => 
                           temp_int_SH_4_port, Z => ML_int_5_23_port);
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => n4, S => 
                           temp_int_SH_4_port, Z => ML_int_5_22_port);
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => n6, S => 
                           temp_int_SH_4_port, Z => ML_int_5_21_port);
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => n2, S => 
                           temp_int_SH_4_port, Z => ML_int_5_20_port);
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => n7, S => 
                           temp_int_SH_4_port, Z => ML_int_5_19_port);
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => n3, S => 
                           temp_int_SH_4_port, Z => ML_int_5_18_port);
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => n5, S => 
                           temp_int_SH_4_port, Z => ML_int_5_17_port);
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => n1, S => 
                           temp_int_SH_4_port, Z => ML_int_5_16_port);
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           temp_int_SH_3_port, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           temp_int_SH_3_port, Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => temp_int_SH_0_port,
                           Z => ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => temp_int_SH_0_port,
                           Z => ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => temp_int_SH_0_port,
                           Z => ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => temp_int_SH_0_port,
                           Z => ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => temp_int_SH_0_port,
                           Z => ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => temp_int_SH_0_port,
                           Z => ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => temp_int_SH_0_port,
                           Z => ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => temp_int_SH_0_port,
                           Z => ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => temp_int_SH_0_port,
                           Z => ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => temp_int_SH_0_port,
                           Z => ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => temp_int_SH_0_port,
                           Z => ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => temp_int_SH_0_port,
                           Z => ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => temp_int_SH_0_port,
                           Z => ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => temp_int_SH_0_port,
                           Z => ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => temp_int_SH_0_port,
                           Z => ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => temp_int_SH_0_port,
                           Z => ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => temp_int_SH_0_port,
                           Z => ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => temp_int_SH_0_port,
                           Z => ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => temp_int_SH_0_port,
                           Z => ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => temp_int_SH_0_port,
                           Z => ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => temp_int_SH_0_port,
                           Z => ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => temp_int_SH_0_port, 
                           Z => ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => temp_int_SH_0_port, Z 
                           => ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => temp_int_SH_0_port, Z 
                           => ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => temp_int_SH_0_port, Z 
                           => ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => temp_int_SH_0_port, Z 
                           => ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => temp_int_SH_0_port, Z 
                           => ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => temp_int_SH_0_port, Z 
                           => ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => temp_int_SH_0_port, Z 
                           => ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => temp_int_SH_0_port, Z 
                           => ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => temp_int_SH_0_port, Z 
                           => ML_int_1_1_port);
   U3 : NAND2_X2 port map( A1 => n38, A2 => n44, ZN => temp_int_SH_1_port);
   U4 : NAND2_X2 port map( A1 => n38, A2 => n45, ZN => temp_int_SH_0_port);
   U5 : NAND2_X2 port map( A1 => n38, A2 => n42, ZN => temp_int_SH_3_port);
   U6 : NAND2_X2 port map( A1 => n38, A2 => n43, ZN => temp_int_SH_2_port);
   U7 : INV_X1 port map( A => n37, ZN => n1);
   U8 : INV_X1 port map( A => n36, ZN => n5);
   U9 : INV_X1 port map( A => n35, ZN => n3);
   U10 : INV_X1 port map( A => n33, ZN => n7);
   U11 : INV_X1 port map( A => n32, ZN => n2);
   U12 : INV_X1 port map( A => n31, ZN => n6);
   U13 : INV_X1 port map( A => n30, ZN => n4);
   U14 : INV_X1 port map( A => n29, ZN => n8);
   U15 : INV_X1 port map( A => n28, ZN => n13);
   U16 : INV_X1 port map( A => temp_int_SH_4_port, ZN => n14);
   U17 : INV_X1 port map( A => temp_int_SH_3_port, ZN => n12);
   U18 : INV_X1 port map( A => temp_int_SH_2_port, ZN => n11);
   U19 : INV_X1 port map( A => temp_int_SH_1_port, ZN => n10);
   U20 : INV_X1 port map( A => SH(25), ZN => n24);
   U21 : INV_X1 port map( A => SH(21), ZN => n23);
   U22 : INV_X1 port map( A => SH(27), ZN => n26);
   U23 : INV_X1 port map( A => SH(9), ZN => n17);
   U24 : INV_X1 port map( A => SH(13), ZN => n18);
   U25 : INV_X1 port map( A => SH(19), ZN => n21);
   U26 : INV_X1 port map( A => SH(15), ZN => n20);
   U27 : INV_X1 port map( A => SH(7), ZN => n15);
   U28 : INV_X1 port map( A => SH(26), ZN => n25);
   U29 : INV_X1 port map( A => SH(8), ZN => n16);
   U30 : INV_X1 port map( A => SH(14), ZN => n19);
   U31 : INV_X1 port map( A => SH(20), ZN => n22);
   U32 : INV_X1 port map( A => SH(30), ZN => n27);
   U33 : INV_X1 port map( A => temp_int_SH_0_port, ZN => n9);
   U34 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n13, ZN => B(9));
   U35 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n13, ZN => B(8));
   U36 : NOR2_X1 port map( A1 => n28, A2 => n29, ZN => B(7));
   U37 : NOR2_X1 port map( A1 => n28, A2 => n30, ZN => B(6));
   U38 : NOR2_X1 port map( A1 => n28, A2 => n31, ZN => B(5));
   U39 : NOR2_X1 port map( A1 => n28, A2 => n32, ZN => B(4));
   U40 : NOR2_X1 port map( A1 => n28, A2 => n33, ZN => B(3));
   U41 : AND2_X1 port map( A1 => ML_int_5_31_port, A2 => n34, ZN => B(31));
   U42 : AND2_X1 port map( A1 => ML_int_5_30_port, A2 => n34, ZN => B(30));
   U43 : NOR2_X1 port map( A1 => n28, A2 => n35, ZN => B(2));
   U44 : AND2_X1 port map( A1 => ML_int_5_29_port, A2 => n34, ZN => B(29));
   U45 : AND2_X1 port map( A1 => ML_int_5_28_port, A2 => n34, ZN => B(28));
   U46 : AND2_X1 port map( A1 => ML_int_5_27_port, A2 => n34, ZN => B(27));
   U47 : AND2_X1 port map( A1 => ML_int_5_26_port, A2 => n34, ZN => B(26));
   U48 : AND2_X1 port map( A1 => ML_int_5_25_port, A2 => n34, ZN => B(25));
   U49 : AND2_X1 port map( A1 => ML_int_5_24_port, A2 => n34, ZN => B(24));
   U50 : AND2_X1 port map( A1 => ML_int_5_23_port, A2 => n34, ZN => B(23));
   U51 : AND2_X1 port map( A1 => ML_int_5_22_port, A2 => n34, ZN => B(22));
   U52 : AND2_X1 port map( A1 => ML_int_5_21_port, A2 => n34, ZN => B(21));
   U53 : AND2_X1 port map( A1 => ML_int_5_20_port, A2 => n34, ZN => B(20));
   U54 : NOR2_X1 port map( A1 => n28, A2 => n36, ZN => B(1));
   U55 : AND2_X1 port map( A1 => ML_int_5_19_port, A2 => n34, ZN => B(19));
   U56 : AND2_X1 port map( A1 => ML_int_5_18_port, A2 => n34, ZN => B(18));
   U57 : AND2_X1 port map( A1 => ML_int_5_17_port, A2 => n34, ZN => B(17));
   U58 : AND2_X1 port map( A1 => ML_int_5_16_port, A2 => n34, ZN => B(16));
   U59 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n13, ZN => B(15));
   U60 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n13, ZN => B(14));
   U61 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n13, ZN => B(13));
   U62 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n13, ZN => B(12));
   U63 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n13, ZN => B(11));
   U64 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n13, ZN => B(10));
   U65 : NOR2_X1 port map( A1 => n28, A2 => n37, ZN => B(0));
   U66 : NAND2_X1 port map( A1 => n34, A2 => n14, ZN => n28);
   U67 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => temp_int_SH_4_port);
   U68 : NAND2_X1 port map( A1 => SH(4), A2 => n40, ZN => n39);
   U69 : AND2_X1 port map( A1 => SHMAG_5_port, A2 => n27, ZN => n34);
   U70 : AND2_X1 port map( A1 => n38, A2 => n41, ZN => SHMAG_5_port);
   U71 : NAND2_X1 port map( A1 => SH(5), A2 => n40, ZN => n41);
   U72 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => n12, ZN => n29);
   U73 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => n12, ZN => n30);
   U74 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => n12, ZN => n31);
   U75 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => n12, ZN => n32);
   U76 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => n12, ZN => n33);
   U77 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => n12, ZN => n35);
   U78 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => n12, ZN => n36);
   U79 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => n12, ZN => n37);
   U80 : NAND2_X1 port map( A1 => SH(3), A2 => n40, ZN => n42);
   U81 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => n11, ZN => 
                           ML_int_3_3_port);
   U82 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => n11, ZN => 
                           ML_int_3_2_port);
   U83 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => n11, ZN => 
                           ML_int_3_1_port);
   U84 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => n11, ZN => 
                           ML_int_3_0_port);
   U85 : NAND2_X1 port map( A1 => SH(2), A2 => n40, ZN => n43);
   U86 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => n10, ZN => 
                           ML_int_2_1_port);
   U87 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => n10, ZN => 
                           ML_int_2_0_port);
   U88 : NAND2_X1 port map( A1 => SH(1), A2 => n40, ZN => n44);
   U89 : AND2_X1 port map( A1 => A(0), A2 => n9, ZN => ML_int_1_0_port);
   U90 : NAND2_X1 port map( A1 => SH(0), A2 => n40, ZN => n45);
   U91 : NAND2_X1 port map( A1 => SH(30), A2 => n46, ZN => n40);
   U92 : NAND4_X1 port map( A1 => n47, A2 => n48, A3 => n49, A4 => n50, ZN => 
                           n46);
   U93 : NOR4_X1 port map( A1 => n51, A2 => n20, A3 => n18, A4 => n19, ZN => 
                           n50);
   U94 : NAND3_X1 port map( A1 => SH(11), A2 => SH(10), A3 => SH(12), ZN => n51
                           );
   U95 : NOR4_X1 port map( A1 => n52, A2 => n23, A3 => n21, A4 => n22, ZN => 
                           n49);
   U96 : NAND3_X1 port map( A1 => SH(17), A2 => SH(16), A3 => SH(18), ZN => n52
                           );
   U97 : NOR4_X1 port map( A1 => n53, A2 => n26, A3 => n24, A4 => n25, ZN => 
                           n48);
   U98 : NAND3_X1 port map( A1 => SH(23), A2 => SH(22), A3 => SH(24), ZN => n53
                           );
   U99 : NOR4_X1 port map( A1 => n54, A2 => n17, A3 => n15, A4 => n16, ZN => 
                           n47);
   U100 : NAND3_X1 port map( A1 => SH(29), A2 => SH(28), A3 => SH(6), ZN => n54
                           );
   U101 : NAND2_X1 port map( A1 => n55, A2 => n27, ZN => n38);
   U102 : NAND4_X1 port map( A1 => n56, A2 => n57, A3 => n58, A4 => n59, ZN => 
                           n55);
   U103 : NOR4_X1 port map( A1 => n60, A2 => SH(28), A3 => SH(6), A4 => SH(29),
                           ZN => n59);
   U104 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => n15, ZN => n60);
   U105 : NOR4_X1 port map( A1 => n61, A2 => SH(22), A3 => SH(24), A4 => SH(23)
                           , ZN => n58);
   U106 : NAND3_X1 port map( A1 => n25, A2 => n26, A3 => n24, ZN => n61);
   U107 : NOR4_X1 port map( A1 => n62, A2 => SH(16), A3 => SH(18), A4 => SH(17)
                           , ZN => n57);
   U108 : NAND3_X1 port map( A1 => n22, A2 => n23, A3 => n21, ZN => n62);
   U109 : NOR4_X1 port map( A1 => n63, A2 => SH(10), A3 => SH(12), A4 => SH(11)
                           , ZN => n56);
   U110 : NAND3_X1 port map( A1 => n19, A2 => n20, A3 => n18, ZN => n63);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity logic_and_shift_N32_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end logic_and_shift_N32_DW_rash_0;

architecture SYN_mx2 of logic_and_shift_N32_DW_rash_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187 : std_logic;

begin
   
   U3 : NOR2_X2 port map( A1 => n52, A2 => SH(1), ZN => n116);
   U4 : NOR2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n117);
   U5 : INV_X1 port map( A => n117, ZN => n49);
   U6 : INV_X1 port map( A => n116, ZN => n51);
   U7 : INV_X1 port map( A => n100, ZN => n50);
   U8 : INV_X1 port map( A => n101, ZN => n53);
   U9 : INV_X1 port map( A => n163, ZN => n59);
   U10 : INV_X1 port map( A => n123, ZN => n56);
   U11 : INV_X1 port map( A => n122, ZN => n58);
   U12 : INV_X1 port map( A => n142, ZN => n54);
   U13 : INV_X1 port map( A => n118, ZN => n46);
   U14 : INV_X1 port map( A => n108, ZN => n47);
   U15 : INV_X1 port map( A => n105, ZN => n55);
   U16 : INV_X1 port map( A => n119, ZN => n44);
   U17 : INV_X1 port map( A => n129, ZN => n35);
   U18 : INV_X1 port map( A => n128, ZN => n37);
   U19 : INV_X1 port map( A => n139, ZN => n40);
   U20 : INV_X1 port map( A => n126, ZN => n32);
   U21 : INV_X1 port map( A => n93, ZN => n17);
   U22 : INV_X1 port map( A => n61, ZN => n10);
   U23 : INV_X1 port map( A => n71, ZN => n8);
   U24 : INV_X1 port map( A => n86, ZN => n12);
   U25 : INV_X1 port map( A => n80, ZN => n14);
   U26 : INV_X1 port map( A => n79, ZN => n21);
   U27 : INV_X1 port map( A => n68, ZN => n19);
   U28 : INV_X1 port map( A => n85, ZN => n20);
   U29 : INV_X1 port map( A => n124, ZN => n33);
   U30 : INV_X1 port map( A => n107, ZN => n48);
   U31 : INV_X1 port map( A => n103, ZN => n6);
   U32 : INV_X1 port map( A => n181, ZN => n45);
   U33 : INV_X1 port map( A => A(26), ZN => n39);
   U34 : INV_X1 port map( A => n165, ZN => n41);
   U35 : INV_X1 port map( A => A(11), ZN => n16);
   U36 : INV_X1 port map( A => n185, ZN => n18);
   U37 : INV_X1 port map( A => n157, ZN => n15);
   U38 : INV_X1 port map( A => n154, ZN => n43);
   U39 : INV_X1 port map( A => A(19), ZN => n28);
   U40 : INV_X1 port map( A => n120, ZN => n42);
   U41 : INV_X1 port map( A => n96, ZN => n60);
   U42 : INV_X1 port map( A => A(2), ZN => n1);
   U43 : INV_X1 port map( A => A(5), ZN => n4);
   U44 : INV_X1 port map( A => A(24), ZN => n36);
   U45 : INV_X1 port map( A => A(4), ZN => n3);
   U46 : INV_X1 port map( A => A(16), ZN => n24);
   U47 : INV_X1 port map( A => SH(2), ZN => n57);
   U48 : INV_X1 port map( A => A(6), ZN => n5);
   U49 : INV_X1 port map( A => A(25), ZN => n38);
   U50 : INV_X1 port map( A => A(23), ZN => n34);
   U51 : INV_X1 port map( A => A(3), ZN => n2);
   U52 : INV_X1 port map( A => A(20), ZN => n29);
   U53 : INV_X1 port map( A => A(21), ZN => n30);
   U54 : INV_X1 port map( A => A(22), ZN => n31);
   U55 : INV_X1 port map( A => A(17), ZN => n26);
   U56 : INV_X1 port map( A => A(15), ZN => n22);
   U57 : INV_X1 port map( A => A(7), ZN => n7);
   U58 : INV_X1 port map( A => A(8), ZN => n9);
   U59 : INV_X1 port map( A => A(9), ZN => n11);
   U60 : INV_X1 port map( A => A(10), ZN => n13);
   U61 : INV_X1 port map( A => SH(0), ZN => n52);
   U62 : INV_X1 port map( A => n141, ZN => n23);
   U63 : INV_X1 port map( A => n134, ZN => n25);
   U64 : INV_X1 port map( A => n113, ZN => n27);
   U65 : OAI221_X1 port map( B1 => n61, B2 => n62, C1 => n63, C2 => n64, A => 
                           n65, ZN => B(9));
   U66 : AOI222_X1 port map( A1 => n54, A2 => n66, B1 => n67, B2 => n68, C1 => 
                           n69, C2 => n70, ZN => n65);
   U67 : OAI221_X1 port map( B1 => n71, B2 => n62, C1 => n72, C2 => n64, A => 
                           n73, ZN => B(8));
   U68 : AOI222_X1 port map( A1 => n54, A2 => n74, B1 => n67, B2 => n17, C1 => 
                           n69, C2 => n75, ZN => n73);
   U69 : OAI221_X1 port map( B1 => n76, B2 => n62, C1 => n33, C2 => n64, A => 
                           n77, ZN => B(7));
   U70 : AOI222_X1 port map( A1 => n54, A2 => n78, B1 => n67, B2 => n14, C1 => 
                           n69, C2 => n79, ZN => n77);
   U71 : OAI221_X1 port map( B1 => n81, B2 => n62, C1 => n82, C2 => n64, A => 
                           n83, ZN => B(6));
   U72 : AOI222_X1 port map( A1 => n54, A2 => n84, B1 => n67, B2 => n12, C1 => 
                           n69, C2 => n85, ZN => n83);
   U73 : OAI221_X1 port map( B1 => n87, B2 => n62, C1 => n88, C2 => n64, A => 
                           n89, ZN => B(5));
   U74 : AOI222_X1 port map( A1 => n54, A2 => n70, B1 => n67, B2 => n10, C1 => 
                           n69, C2 => n68, ZN => n89);
   U75 : OAI221_X1 port map( B1 => n90, B2 => n62, C1 => n91, C2 => n64, A => 
                           n92, ZN => B(4));
   U76 : AOI222_X1 port map( A1 => n54, A2 => n75, B1 => n67, B2 => n8, C1 => 
                           n69, C2 => n17, ZN => n92);
   U77 : AOI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => B(3));
   U78 : OAI21_X1 port map( B1 => n97, B2 => n98, A => n99, ZN => n95);
   U79 : OAI22_X1 port map( A1 => n49, A2 => n2, B1 => n51, B2 => n3, ZN => n98
                           );
   U80 : OAI22_X1 port map( A1 => n100, A2 => n4, B1 => n101, B2 => n5, ZN => 
                           n97);
   U81 : MUX2_X1 port map( A => n6, B => n102, S => SH(4), Z => n94);
   U82 : OAI222_X1 port map( A1 => n56, A2 => n76, B1 => n104, B2 => n21, C1 =>
                           n105, C2 => n80, ZN => n103);
   U83 : AOI221_X1 port map( B1 => n53, B2 => A(10), C1 => n50, C2 => A(9), A 
                           => n106, ZN => n76);
   U84 : OAI22_X1 port map( A1 => n9, A2 => n51, B1 => n7, B2 => n49, ZN => 
                           n106);
   U85 : NOR2_X1 port map( A1 => n62, A2 => n107, ZN => B(31));
   U86 : NOR2_X1 port map( A1 => n108, A2 => n62, ZN => B(30));
   U87 : NOR2_X1 port map( A1 => n109, A2 => n96, ZN => B(2));
   U88 : AOI21_X1 port map( B1 => n99, B2 => n110, A => n111, ZN => n109);
   U89 : MUX2_X1 port map( A => n112, B => n27, S => SH(4), Z => n111);
   U90 : OAI222_X1 port map( A1 => n86, A2 => n105, B1 => n20, B2 => n104, C1 
                           => n81, C2 => n56, ZN => n112);
   U91 : AOI221_X1 port map( B1 => n53, B2 => A(9), C1 => n50, C2 => A(8), A =>
                           n114, ZN => n81);
   U92 : OAI22_X1 port map( A1 => n7, A2 => n51, B1 => n5, B2 => n49, ZN => 
                           n114);
   U93 : OAI221_X1 port map( B1 => n101, B2 => n4, C1 => n100, C2 => n3, A => 
                           n115, ZN => n110);
   U94 : AOI22_X1 port map( A1 => A(3), A2 => n116, B1 => A(2), B2 => n117, ZN 
                           => n115);
   U95 : NOR2_X1 port map( A1 => n118, A2 => n62, ZN => B(29));
   U96 : NOR2_X1 port map( A1 => n119, A2 => n62, ZN => B(28));
   U97 : NOR3_X1 port map( A1 => n59, A2 => SH(3), A3 => n120, ZN => B(27));
   U98 : NOR2_X1 port map( A1 => n121, A2 => n59, ZN => B(26));
   U99 : NOR2_X1 port map( A1 => n63, A2 => n59, ZN => B(25));
   U100 : AOI22_X1 port map( A1 => n37, A2 => n122, B1 => n46, B2 => n123, ZN 
                           => n63);
   U101 : NOR2_X1 port map( A1 => n72, A2 => n59, ZN => B(24));
   U102 : AOI22_X1 port map( A1 => n35, A2 => n122, B1 => n44, B2 => n123, ZN 
                           => n72);
   U103 : NOR2_X1 port map( A1 => n33, A2 => n59, ZN => B(23));
   U104 : OAI222_X1 port map( A1 => n125, A2 => n56, B1 => n107, B2 => n105, C1
                           => n126, C2 => n58, ZN => n124);
   U105 : NOR2_X1 port map( A1 => n82, A2 => n59, ZN => B(22));
   U106 : AOI222_X1 port map( A1 => n40, A2 => n123, B1 => n47, B2 => n55, C1 
                           => n127, C2 => n122, ZN => n82);
   U107 : NOR2_X1 port map( A1 => n88, A2 => n59, ZN => B(21));
   U108 : AOI222_X1 port map( A1 => n37, A2 => n123, B1 => n46, B2 => n55, C1 
                           => n66, C2 => n122, ZN => n88);
   U109 : NOR2_X1 port map( A1 => n91, A2 => n59, ZN => B(20));
   U110 : AOI222_X1 port map( A1 => n35, A2 => n123, B1 => n44, B2 => n55, C1 
                           => n74, C2 => n122, ZN => n91);
   U111 : NOR2_X1 port map( A1 => n130, A2 => n96, ZN => B(1));
   U112 : AOI21_X1 port map( B1 => n99, B2 => n131, A => n132, ZN => n130);
   U113 : MUX2_X1 port map( A => n133, B => n25, S => SH(4), Z => n132);
   U114 : OAI222_X1 port map( A1 => n61, A2 => n105, B1 => n19, B2 => n104, C1 
                           => n87, C2 => n56, ZN => n133);
   U115 : AOI221_X1 port map( B1 => n53, B2 => A(8), C1 => n50, C2 => A(7), A 
                           => n135, ZN => n87);
   U116 : OAI22_X1 port map( A1 => n5, A2 => n51, B1 => n4, B2 => n49, ZN => 
                           n135);
   U117 : AOI221_X1 port map( B1 => n53, B2 => A(12), C1 => n50, C2 => A(11), A
                           => n136, ZN => n61);
   U118 : OAI22_X1 port map( A1 => n13, A2 => n51, B1 => n11, B2 => n49, ZN => 
                           n136);
   U119 : OAI221_X1 port map( B1 => n101, B2 => n3, C1 => n100, C2 => n2, A => 
                           n137, ZN => n131);
   U120 : AOI22_X1 port map( A1 => A(2), A2 => n116, B1 => A(1), B2 => n117, ZN
                           => n137);
   U121 : NOR2_X1 port map( A1 => n102, A2 => n59, ZN => B(19));
   U122 : AOI222_X1 port map( A1 => n78, A2 => n122, B1 => n32, B2 => n123, C1 
                           => n42, C2 => SH(3), ZN => n102);
   U123 : NOR2_X1 port map( A1 => n113, A2 => n59, ZN => B(18));
   U124 : AOI221_X1 port map( B1 => n127, B2 => n123, C1 => n84, C2 => n122, A 
                           => n138, ZN => n113);
   U125 : OAI22_X1 port map( A1 => n104, A2 => n108, B1 => n105, B2 => n139, ZN
                           => n138);
   U126 : NOR2_X1 port map( A1 => n134, A2 => n59, ZN => B(17));
   U127 : AOI221_X1 port map( B1 => n66, B2 => n123, C1 => n70, C2 => n122, A 
                           => n140, ZN => n134);
   U128 : OAI22_X1 port map( A1 => n104, A2 => n118, B1 => n105, B2 => n128, ZN
                           => n140);
   U129 : NOR2_X1 port map( A1 => n141, A2 => n59, ZN => B(16));
   U130 : OAI221_X1 port map( B1 => n125, B2 => n142, C1 => n21, C2 => n62, A 
                           => n143, ZN => B(15));
   U131 : AOI222_X1 port map( A1 => n69, A2 => n32, B1 => n144, B2 => n48, C1 
                           => n67, C2 => n78, ZN => n143);
   U132 : OAI221_X1 port map( B1 => n139, B2 => n142, C1 => n20, C2 => n62, A 
                           => n145, ZN => B(14));
   U133 : AOI222_X1 port map( A1 => n69, A2 => n127, B1 => n144, B2 => n47, C1 
                           => n67, C2 => n84, ZN => n145);
   U134 : OAI221_X1 port map( B1 => n128, B2 => n142, C1 => n19, C2 => n62, A 
                           => n146, ZN => B(13));
   U135 : AOI222_X1 port map( A1 => n69, A2 => n66, B1 => n144, B2 => n46, C1 
                           => n67, C2 => n70, ZN => n146);
   U136 : OAI221_X1 port map( B1 => n101, B2 => n29, C1 => n100, C2 => n28, A 
                           => n147, ZN => n70);
   U137 : AOI22_X1 port map( A1 => A(18), A2 => n116, B1 => A(17), B2 => n117, 
                           ZN => n147);
   U138 : AOI222_X1 port map( A1 => n116, A2 => A(30), B1 => n50, B2 => A(31), 
                           C1 => n117, C2 => A(29), ZN => n118);
   U139 : OAI221_X1 port map( B1 => n101, B2 => n36, C1 => n100, C2 => n34, A 
                           => n148, ZN => n66);
   U140 : AOI22_X1 port map( A1 => A(22), A2 => n116, B1 => A(21), B2 => n117, 
                           ZN => n148);
   U141 : OAI221_X1 port map( B1 => n101, B2 => n24, C1 => n100, C2 => n22, A 
                           => n149, ZN => n68);
   U142 : AOI22_X1 port map( A1 => A(14), A2 => n116, B1 => A(13), B2 => n117, 
                           ZN => n149);
   U143 : AOI221_X1 port map( B1 => n53, B2 => A(28), C1 => n50, C2 => A(27), A
                           => n150, ZN => n128);
   U144 : OAI22_X1 port map( A1 => n39, A2 => n51, B1 => n38, B2 => n49, ZN => 
                           n150);
   U145 : OAI221_X1 port map( B1 => n129, B2 => n142, C1 => n93, C2 => n62, A 
                           => n151, ZN => B(12));
   U146 : AOI222_X1 port map( A1 => n69, A2 => n74, B1 => n144, B2 => n44, C1 
                           => n67, C2 => n75, ZN => n151);
   U147 : NOR2_X1 port map( A1 => n64, A2 => n58, ZN => n144);
   U148 : OAI221_X1 port map( B1 => n126, B2 => n142, C1 => n80, C2 => n62, A 
                           => n152, ZN => B(11));
   U149 : AOI221_X1 port map( B1 => n69, B2 => n78, C1 => n67, C2 => n79, A => 
                           n153, ZN => n152);
   U150 : NOR3_X1 port map( A1 => n64, A2 => SH(3), A3 => n120, ZN => n153);
   U151 : MUX2_X1 port map( A => n125, B => n107, S => SH(2), Z => n120);
   U152 : NAND2_X1 port map( A1 => A(31), A2 => n117, ZN => n107);
   U153 : AOI221_X1 port map( B1 => n53, B2 => A(30), C1 => n50, C2 => A(29), A
                           => n43, ZN => n125);
   U154 : AOI22_X1 port map( A1 => A(28), A2 => n116, B1 => A(27), B2 => n117, 
                           ZN => n154);
   U155 : OAI221_X1 port map( B1 => n24, B2 => n51, C1 => n22, C2 => n49, A => 
                           n155, ZN => n79);
   U156 : AOI22_X1 port map( A1 => A(18), A2 => n53, B1 => A(17), B2 => n50, ZN
                           => n155);
   U157 : OAI221_X1 port map( B1 => n101, B2 => n31, C1 => n100, C2 => n30, A 
                           => n156, ZN => n78);
   U158 : AOI22_X1 port map( A1 => A(20), A2 => n116, B1 => A(19), B2 => n117, 
                           ZN => n156);
   U159 : AOI221_X1 port map( B1 => n53, B2 => A(14), C1 => n50, C2 => A(13), A
                           => n15, ZN => n80);
   U160 : AOI22_X1 port map( A1 => A(12), A2 => n116, B1 => A(11), B2 => n117, 
                           ZN => n157);
   U161 : AOI221_X1 port map( B1 => n53, B2 => A(26), C1 => n50, C2 => A(25), A
                           => n158, ZN => n126);
   U162 : OAI22_X1 port map( A1 => n36, A2 => n51, B1 => n34, B2 => n49, ZN => 
                           n158);
   U163 : OAI221_X1 port map( B1 => n86, B2 => n62, C1 => n121, C2 => n64, A =>
                           n159, ZN => B(10));
   U164 : AOI222_X1 port map( A1 => n54, A2 => n127, B1 => n67, B2 => n85, C1 
                           => n69, C2 => n84, ZN => n159);
   U165 : OAI221_X1 port map( B1 => n101, B2 => n30, C1 => n100, C2 => n29, A 
                           => n160, ZN => n84);
   U166 : AOI22_X1 port map( A1 => A(19), A2 => n116, B1 => A(18), B2 => n117, 
                           ZN => n160);
   U167 : AND2_X1 port map( A1 => n161, A2 => n57, ZN => n69);
   U168 : OAI221_X1 port map( B1 => n101, B2 => n26, C1 => n24, C2 => n100, A 
                           => n162, ZN => n85);
   U169 : AOI22_X1 port map( A1 => n116, A2 => A(15), B1 => n117, B2 => A(14), 
                           ZN => n162);
   U170 : NOR2_X1 port map( A1 => n59, A2 => n56, ZN => n67);
   U171 : OAI221_X1 port map( B1 => n101, B2 => n38, C1 => n100, C2 => n36, A 
                           => n164, ZN => n127);
   U172 : AOI22_X1 port map( A1 => A(23), A2 => n116, B1 => A(22), B2 => n117, 
                           ZN => n164);
   U173 : NAND2_X1 port map( A1 => n161, A2 => SH(2), ZN => n142);
   U174 : AND2_X1 port map( A1 => SH(3), A2 => n163, ZN => n161);
   U175 : NAND2_X1 port map( A1 => SH(4), A2 => n60, ZN => n64);
   U176 : AOI22_X1 port map( A1 => n40, A2 => n122, B1 => n47, B2 => n123, ZN 
                           => n121);
   U177 : AOI22_X1 port map( A1 => n117, A2 => A(30), B1 => n116, B2 => A(31), 
                           ZN => n108);
   U178 : AOI221_X1 port map( B1 => n53, B2 => A(29), C1 => n50, C2 => A(28), A
                           => n41, ZN => n139);
   U179 : AOI22_X1 port map( A1 => A(27), A2 => n116, B1 => A(26), B2 => n117, 
                           ZN => n165);
   U180 : NAND2_X1 port map( A1 => n122, A2 => n163, ZN => n62);
   U181 : NOR2_X1 port map( A1 => n96, A2 => SH(4), ZN => n163);
   U182 : AOI221_X1 port map( B1 => n53, B2 => A(13), C1 => n50, C2 => A(12), A
                           => n166, ZN => n86);
   U183 : OAI22_X1 port map( A1 => n16, A2 => n51, B1 => n13, B2 => n49, ZN => 
                           n166);
   U184 : NOR2_X1 port map( A1 => n167, A2 => n96, ZN => B(0));
   U185 : NAND4_X1 port map( A1 => n168, A2 => n169, A3 => n170, A4 => n171, ZN
                           => n96);
   U186 : NOR4_X1 port map( A1 => n172, A2 => SH(29), A3 => SH(5), A4 => SH(30)
                           , ZN => n171);
   U187 : OR4_X1 port map( A1 => SH(7), A2 => SH(6), A3 => SH(9), A4 => SH(8), 
                           ZN => n172);
   U188 : NOR4_X1 port map( A1 => n173, A2 => SH(23), A3 => SH(25), A4 => 
                           SH(24), ZN => n170);
   U189 : OR3_X1 port map( A1 => SH(28), A2 => SH(27), A3 => SH(26), ZN => n173
                           );
   U190 : NOR4_X1 port map( A1 => n174, A2 => SH(16), A3 => SH(18), A4 => 
                           SH(17), ZN => n169);
   U191 : OR4_X1 port map( A1 => SH(20), A2 => SH(19), A3 => SH(22), A4 => 
                           SH(21), ZN => n174);
   U192 : NOR4_X1 port map( A1 => n175, A2 => SH(10), A3 => SH(12), A4 => 
                           SH(11), ZN => n168);
   U193 : OR3_X1 port map( A1 => SH(15), A2 => SH(14), A3 => SH(13), ZN => n175
                           );
   U194 : AOI21_X1 port map( B1 => n99, B2 => n176, A => n177, ZN => n167);
   U195 : MUX2_X1 port map( A => n178, B => n23, S => SH(4), Z => n177);
   U196 : AOI221_X1 port map( B1 => n74, B2 => n123, C1 => n75, C2 => n122, A 
                           => n179, ZN => n141);
   U197 : OAI22_X1 port map( A1 => n104, A2 => n119, B1 => n105, B2 => n129, ZN
                           => n179);
   U198 : AOI221_X1 port map( B1 => n53, B2 => A(27), C1 => n50, C2 => A(26), A
                           => n180, ZN => n129);
   U199 : OAI22_X1 port map( A1 => n38, A2 => n51, B1 => n36, B2 => n49, ZN => 
                           n180);
   U200 : AOI221_X1 port map( B1 => n53, B2 => A(31), C1 => n50, C2 => A(30), A
                           => n45, ZN => n119);
   U201 : AOI22_X1 port map( A1 => A(29), A2 => n116, B1 => A(28), B2 => n117, 
                           ZN => n181);
   U202 : OAI221_X1 port map( B1 => n51, B2 => n26, C1 => n24, C2 => n49, A => 
                           n182, ZN => n75);
   U203 : AOI22_X1 port map( A1 => A(19), A2 => n53, B1 => A(18), B2 => n50, ZN
                           => n182);
   U204 : OAI221_X1 port map( B1 => n101, B2 => n34, C1 => n100, C2 => n31, A 
                           => n183, ZN => n74);
   U205 : AOI22_X1 port map( A1 => A(21), A2 => n116, B1 => A(20), B2 => n117, 
                           ZN => n183);
   U206 : OAI222_X1 port map( A1 => n71, A2 => n105, B1 => n93, B2 => n104, C1 
                           => n90, C2 => n56, ZN => n178);
   U207 : NOR2_X1 port map( A1 => n57, A2 => SH(3), ZN => n123);
   U208 : AOI221_X1 port map( B1 => n53, B2 => A(7), C1 => n50, C2 => A(6), A 
                           => n184, ZN => n90);
   U209 : OAI22_X1 port map( A1 => n4, A2 => n51, B1 => n3, B2 => n49, ZN => 
                           n184);
   U210 : NAND2_X1 port map( A1 => SH(3), A2 => SH(2), ZN => n104);
   U211 : AOI221_X1 port map( B1 => n53, B2 => A(15), C1 => n50, C2 => A(14), A
                           => n18, ZN => n93);
   U212 : AOI22_X1 port map( A1 => A(13), A2 => n116, B1 => A(12), B2 => n117, 
                           ZN => n185);
   U213 : NAND2_X1 port map( A1 => SH(3), A2 => n57, ZN => n105);
   U214 : AOI221_X1 port map( B1 => n53, B2 => A(11), C1 => n50, C2 => A(10), A
                           => n186, ZN => n71);
   U215 : OAI22_X1 port map( A1 => n11, A2 => n51, B1 => n9, B2 => n49, ZN => 
                           n186);
   U216 : OAI221_X1 port map( B1 => n101, B2 => n2, C1 => n100, C2 => n1, A => 
                           n187, ZN => n176);
   U217 : AOI22_X1 port map( A1 => A(1), A2 => n116, B1 => A(0), B2 => n117, ZN
                           => n187);
   U218 : NAND2_X1 port map( A1 => SH(1), A2 => n52, ZN => n100);
   U219 : NAND2_X1 port map( A1 => SH(1), A2 => SH(0), ZN => n101);
   U220 : NOR2_X1 port map( A1 => n58, A2 => SH(4), ZN => n99);
   U221 : NOR2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n122);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_7;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U2 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_6;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U2 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_5;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U2 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_4;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U2 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_3;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U2 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_2;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U2 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_1;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U2 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_15;

architecture SYN_BEHAVIORAL of RCA_NBITS4_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_14;

architecture SYN_BEHAVIORAL of RCA_NBITS4_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_13;

architecture SYN_BEHAVIORAL of RCA_NBITS4_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_12;

architecture SYN_BEHAVIORAL of RCA_NBITS4_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_11;

architecture SYN_BEHAVIORAL of RCA_NBITS4_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_10;

architecture SYN_BEHAVIORAL of RCA_NBITS4_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_9;

architecture SYN_BEHAVIORAL of RCA_NBITS4_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_8;

architecture SYN_BEHAVIORAL of RCA_NBITS4_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_7;

architecture SYN_BEHAVIORAL of RCA_NBITS4_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_6;

architecture SYN_BEHAVIORAL of RCA_NBITS4_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_5;

architecture SYN_BEHAVIORAL of RCA_NBITS4_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_4;

architecture SYN_BEHAVIORAL of RCA_NBITS4_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_3;

architecture SYN_BEHAVIORAL of RCA_NBITS4_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_2;

architecture SYN_BEHAVIORAL of RCA_NBITS4_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_1;

architecture SYN_BEHAVIORAL of RCA_NBITS4_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_26 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_26;

architecture SYN_BEHAVIORAL of PG_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_25 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_25;

architecture SYN_BEHAVIORAL of PG_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_24 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_24;

architecture SYN_BEHAVIORAL of PG_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_23 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_23;

architecture SYN_BEHAVIORAL of PG_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_22 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_22;

architecture SYN_BEHAVIORAL of PG_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_21 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_21;

architecture SYN_BEHAVIORAL of PG_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_20 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_20;

architecture SYN_BEHAVIORAL of PG_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_19 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_19;

architecture SYN_BEHAVIORAL of PG_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_18 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_18;

architecture SYN_BEHAVIORAL of PG_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_17 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_17;

architecture SYN_BEHAVIORAL of PG_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_16 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_16;

architecture SYN_BEHAVIORAL of PG_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_15 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_15;

architecture SYN_BEHAVIORAL of PG_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_14 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_14;

architecture SYN_BEHAVIORAL of PG_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_13 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_13;

architecture SYN_BEHAVIORAL of PG_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_12 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_12;

architecture SYN_BEHAVIORAL of PG_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_11 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_11;

architecture SYN_BEHAVIORAL of PG_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_10 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_10;

architecture SYN_BEHAVIORAL of PG_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_9 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_9;

architecture SYN_BEHAVIORAL of PG_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_8 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_8;

architecture SYN_BEHAVIORAL of PG_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_7 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_7;

architecture SYN_BEHAVIORAL of PG_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_6 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_6;

architecture SYN_BEHAVIORAL of PG_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_5 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_5;

architecture SYN_BEHAVIORAL of PG_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_4 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_4;

architecture SYN_BEHAVIORAL of PG_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_3 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_3;

architecture SYN_BEHAVIORAL of PG_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_2 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_2;

architecture SYN_BEHAVIORAL of PG_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_1 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_1;

architecture SYN_BEHAVIORAL of PG_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_8 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_8;

architecture SYN_BEHAVIORAL of G_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_7 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_7;

architecture SYN_BEHAVIORAL of G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_6 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_6;

architecture SYN_BEHAVIORAL of G_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_5 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_5;

architecture SYN_BEHAVIORAL of G_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_4 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_4;

architecture SYN_BEHAVIORAL of G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_3 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_3;

architecture SYN_BEHAVIORAL of G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_2 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_2;

architecture SYN_BEHAVIORAL of G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_1 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_1;

architecture SYN_BEHAVIORAL of G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_31 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_31;

architecture SYN_BEHAVIORAL of pg_generator_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_30 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_30;

architecture SYN_BEHAVIORAL of pg_generator_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_29 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_29;

architecture SYN_BEHAVIORAL of pg_generator_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_28 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_28;

architecture SYN_BEHAVIORAL of pg_generator_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_27 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_27;

architecture SYN_BEHAVIORAL of pg_generator_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_26 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_26;

architecture SYN_BEHAVIORAL of pg_generator_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_25 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_25;

architecture SYN_BEHAVIORAL of pg_generator_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_24 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_24;

architecture SYN_BEHAVIORAL of pg_generator_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_23 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_23;

architecture SYN_BEHAVIORAL of pg_generator_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_22 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_22;

architecture SYN_BEHAVIORAL of pg_generator_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_21 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_21;

architecture SYN_BEHAVIORAL of pg_generator_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_20 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_20;

architecture SYN_BEHAVIORAL of pg_generator_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_19 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_19;

architecture SYN_BEHAVIORAL of pg_generator_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_18 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_18;

architecture SYN_BEHAVIORAL of pg_generator_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_17 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_17;

architecture SYN_BEHAVIORAL of pg_generator_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_16 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_16;

architecture SYN_BEHAVIORAL of pg_generator_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_15 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_15;

architecture SYN_BEHAVIORAL of pg_generator_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_14 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_14;

architecture SYN_BEHAVIORAL of pg_generator_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_13 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_13;

architecture SYN_BEHAVIORAL of pg_generator_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_12 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_12;

architecture SYN_BEHAVIORAL of pg_generator_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_11 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_11;

architecture SYN_BEHAVIORAL of pg_generator_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_10 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_10;

architecture SYN_BEHAVIORAL of pg_generator_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_9 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_9;

architecture SYN_BEHAVIORAL of pg_generator_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_8 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_8;

architecture SYN_BEHAVIORAL of pg_generator_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_7 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_7;

architecture SYN_BEHAVIORAL of pg_generator_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_6 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_6;

architecture SYN_BEHAVIORAL of pg_generator_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_5 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_5;

architecture SYN_BEHAVIORAL of pg_generator_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_4 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_4;

architecture SYN_BEHAVIORAL of pg_generator_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_3 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_3;

architecture SYN_BEHAVIORAL of pg_generator_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_2 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_2;

architecture SYN_BEHAVIORAL of pg_generator_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_1 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_1;

architecture SYN_BEHAVIORAL of pg_generator_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_7;

architecture SYN_STRUCTURAL of CarrySelect_7 is

   component MUX21_GENERIC_bits4_7
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1004, n_1005 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1004);
   RCA2 : RCA_NBITS4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1005);
   MUX21_GEN : MUX21_GENERIC_bits4_7 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_6;

architecture SYN_STRUCTURAL of CarrySelect_6 is

   component MUX21_GENERIC_bits4_6
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1006, n_1007 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1006);
   RCA2 : RCA_NBITS4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1007);
   MUX21_GEN : MUX21_GENERIC_bits4_6 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_5;

architecture SYN_STRUCTURAL of CarrySelect_5 is

   component MUX21_GENERIC_bits4_5
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1008, n_1009 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1008);
   RCA2 : RCA_NBITS4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1009);
   MUX21_GEN : MUX21_GENERIC_bits4_5 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_4;

architecture SYN_STRUCTURAL of CarrySelect_4 is

   component MUX21_GENERIC_bits4_4
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1010, n_1011 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1010);
   RCA2 : RCA_NBITS4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1011);
   MUX21_GEN : MUX21_GENERIC_bits4_4 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_3;

architecture SYN_STRUCTURAL of CarrySelect_3 is

   component MUX21_GENERIC_bits4_3
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1012, n_1013 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1012);
   RCA2 : RCA_NBITS4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1013);
   MUX21_GEN : MUX21_GENERIC_bits4_3 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_2;

architecture SYN_STRUCTURAL of CarrySelect_2 is

   component MUX21_GENERIC_bits4_2
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1014, n_1015 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1014);
   RCA2 : RCA_NBITS4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1015);
   MUX21_GEN : MUX21_GENERIC_bits4_2 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_1;

architecture SYN_STRUCTURAL of CarrySelect_1 is

   component MUX21_GENERIC_bits4_1
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1016, n_1017 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1016);
   RCA2 : RCA_NBITS4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1017);
   MUX21_GEN : MUX21_GENERIC_bits4_1 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_352 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_352;

architecture SYN_ASYNCH_FD of FD_352 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1018 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1018);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_351 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_351;

architecture SYN_ASYNCH_FD of FD_351 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1019 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1019);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_350 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_350;

architecture SYN_ASYNCH_FD of FD_350 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1020 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1020);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_349 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_349;

architecture SYN_ASYNCH_FD of FD_349 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1021 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1021);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_348 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_348;

architecture SYN_ASYNCH_FD of FD_348 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1022 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1022);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_347 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_347;

architecture SYN_ASYNCH_FD of FD_347 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1023 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1023);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_346 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_346;

architecture SYN_ASYNCH_FD of FD_346 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1024 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1024);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_345 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_345;

architecture SYN_ASYNCH_FD of FD_345 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1025 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1025);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_344 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_344;

architecture SYN_ASYNCH_FD of FD_344 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1026 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1026);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_343 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_343;

architecture SYN_ASYNCH_FD of FD_343 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1027 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1027);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_342 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_342;

architecture SYN_ASYNCH_FD of FD_342 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1028 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1028);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_341 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_341;

architecture SYN_ASYNCH_FD of FD_341 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1029 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1029);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_340 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_340;

architecture SYN_ASYNCH_FD of FD_340 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1030 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1030);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_339 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_339;

architecture SYN_ASYNCH_FD of FD_339 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1031 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1031);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_338 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_338;

architecture SYN_ASYNCH_FD of FD_338 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1032 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1032);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_337 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_337;

architecture SYN_ASYNCH_FD of FD_337 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1033 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1033);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_336 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_336;

architecture SYN_ASYNCH_FD of FD_336 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1034 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1034);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_335 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_335;

architecture SYN_ASYNCH_FD of FD_335 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1035 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1035);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_334 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_334;

architecture SYN_ASYNCH_FD of FD_334 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1036 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1036);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_333 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_333;

architecture SYN_ASYNCH_FD of FD_333 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1037 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1037);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_332 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_332;

architecture SYN_ASYNCH_FD of FD_332 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1038 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1038);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_331 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_331;

architecture SYN_ASYNCH_FD of FD_331 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1039 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1039);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_330 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_330;

architecture SYN_ASYNCH_FD of FD_330 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1040 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1040);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_329 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_329;

architecture SYN_ASYNCH_FD of FD_329 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1041 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1041);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_328 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_328;

architecture SYN_ASYNCH_FD of FD_328 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1042 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1042);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_327 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_327;

architecture SYN_ASYNCH_FD of FD_327 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1043 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1043);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_326 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_326;

architecture SYN_ASYNCH_FD of FD_326 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1044 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1044);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_325 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_325;

architecture SYN_ASYNCH_FD of FD_325 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1045 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1045);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_324 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_324;

architecture SYN_ASYNCH_FD of FD_324 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1046 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1046);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_323 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_323;

architecture SYN_ASYNCH_FD of FD_323 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1047 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1047);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_322 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_322;

architecture SYN_ASYNCH_FD of FD_322 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1048 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1048);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_321 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_321;

architecture SYN_ASYNCH_FD of FD_321 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1049 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1049);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_320 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_320;

architecture SYN_ASYNCH_FD of FD_320 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1050 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1050);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_319 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_319;

architecture SYN_ASYNCH_FD of FD_319 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1051 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1051);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_318 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_318;

architecture SYN_ASYNCH_FD of FD_318 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1052 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1052);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_317 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_317;

architecture SYN_ASYNCH_FD of FD_317 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1053 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1053);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_316 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_316;

architecture SYN_ASYNCH_FD of FD_316 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1054 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1054);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_315 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_315;

architecture SYN_ASYNCH_FD of FD_315 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1055 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1055);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_314 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_314;

architecture SYN_ASYNCH_FD of FD_314 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1056 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1056);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_313 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_313;

architecture SYN_ASYNCH_FD of FD_313 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1057 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1057);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_312 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_312;

architecture SYN_ASYNCH_FD of FD_312 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1058 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1058);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_311 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_311;

architecture SYN_ASYNCH_FD of FD_311 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1059 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1059);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_310 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_310;

architecture SYN_ASYNCH_FD of FD_310 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1060 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1060);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_309 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_309;

architecture SYN_ASYNCH_FD of FD_309 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1061 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1061);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_308 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_308;

architecture SYN_ASYNCH_FD of FD_308 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1062 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1062);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_307 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_307;

architecture SYN_ASYNCH_FD of FD_307 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1063 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1063);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_306 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_306;

architecture SYN_ASYNCH_FD of FD_306 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1064 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1064);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_305 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_305;

architecture SYN_ASYNCH_FD of FD_305 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1065 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1065);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_304 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_304;

architecture SYN_ASYNCH_FD of FD_304 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1066 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1066);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_303 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_303;

architecture SYN_ASYNCH_FD of FD_303 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1067 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1067);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_302 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_302;

architecture SYN_ASYNCH_FD of FD_302 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1068 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1068);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_301 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_301;

architecture SYN_ASYNCH_FD of FD_301 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1069 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1069);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_300 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_300;

architecture SYN_ASYNCH_FD of FD_300 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1070 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1070);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_299 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_299;

architecture SYN_ASYNCH_FD of FD_299 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1071 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1071);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_298 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_298;

architecture SYN_ASYNCH_FD of FD_298 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1072 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1072);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_297 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_297;

architecture SYN_ASYNCH_FD of FD_297 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1073 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1073);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_296 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_296;

architecture SYN_ASYNCH_FD of FD_296 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1074 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1074);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_295 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_295;

architecture SYN_ASYNCH_FD of FD_295 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1075 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1075);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_294 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_294;

architecture SYN_ASYNCH_FD of FD_294 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1076 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1076);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_293 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_293;

architecture SYN_ASYNCH_FD of FD_293 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1077 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1077);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_292 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_292;

architecture SYN_ASYNCH_FD of FD_292 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1078 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1078);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_291 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_291;

architecture SYN_ASYNCH_FD of FD_291 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1079 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1079);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_290 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_290;

architecture SYN_ASYNCH_FD of FD_290 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1080 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1080);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_289 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_289;

architecture SYN_ASYNCH_FD of FD_289 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1081 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1081);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_288 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_288;

architecture SYN_ASYNCH_FD of FD_288 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1082 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1082);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_287 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_287;

architecture SYN_ASYNCH_FD of FD_287 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1083 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1083);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_286 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_286;

architecture SYN_ASYNCH_FD of FD_286 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1084 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1084);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_285 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_285;

architecture SYN_ASYNCH_FD of FD_285 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1085 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1085);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_284 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_284;

architecture SYN_ASYNCH_FD of FD_284 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1086 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1086);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_283 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_283;

architecture SYN_ASYNCH_FD of FD_283 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1087 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1087);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_282 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_282;

architecture SYN_ASYNCH_FD of FD_282 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1088 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1088);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_281 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_281;

architecture SYN_ASYNCH_FD of FD_281 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1089 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1089);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_280 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_280;

architecture SYN_ASYNCH_FD of FD_280 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1090 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1090);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_279 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_279;

architecture SYN_ASYNCH_FD of FD_279 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1091 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1091);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_278 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_278;

architecture SYN_ASYNCH_FD of FD_278 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1092 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1092);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_277 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_277;

architecture SYN_ASYNCH_FD of FD_277 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1093 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1093);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_276 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_276;

architecture SYN_ASYNCH_FD of FD_276 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1094 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1094);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_275 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_275;

architecture SYN_ASYNCH_FD of FD_275 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1095 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1095);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_274 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_274;

architecture SYN_ASYNCH_FD of FD_274 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1096 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1096);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_273 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_273;

architecture SYN_ASYNCH_FD of FD_273 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1097 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1097);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_272 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_272;

architecture SYN_ASYNCH_FD of FD_272 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1098 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1098);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_271 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_271;

architecture SYN_ASYNCH_FD of FD_271 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1099 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1099);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_270 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_270;

architecture SYN_ASYNCH_FD of FD_270 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1100 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1100);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_269 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_269;

architecture SYN_ASYNCH_FD of FD_269 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1101 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1101);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_268 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_268;

architecture SYN_ASYNCH_FD of FD_268 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1102 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1102);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_267 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_267;

architecture SYN_ASYNCH_FD of FD_267 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1103 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1103);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_266 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_266;

architecture SYN_ASYNCH_FD of FD_266 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1104 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1104);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_265 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_265;

architecture SYN_ASYNCH_FD of FD_265 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1105 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1105);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_264 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_264;

architecture SYN_ASYNCH_FD of FD_264 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1106 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1106);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_263 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_263;

architecture SYN_ASYNCH_FD of FD_263 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1107 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1107);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_262 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_262;

architecture SYN_ASYNCH_FD of FD_262 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1108 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1108);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_261 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_261;

architecture SYN_ASYNCH_FD of FD_261 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1109 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1109);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_260 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_260;

architecture SYN_ASYNCH_FD of FD_260 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1110 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1110);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_259 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_259;

architecture SYN_ASYNCH_FD of FD_259 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1111 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1111);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_258 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_258;

architecture SYN_ASYNCH_FD of FD_258 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1112 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1112);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_257 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_257;

architecture SYN_ASYNCH_FD of FD_257 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1113 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1113);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_256 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_256;

architecture SYN_ASYNCH_FD of FD_256 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1114 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1114);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_255 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_255;

architecture SYN_ASYNCH_FD of FD_255 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1115 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1115);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_254 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_254;

architecture SYN_ASYNCH_FD of FD_254 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1116 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1116);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_253 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_253;

architecture SYN_ASYNCH_FD of FD_253 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1117 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1117);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_252 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_252;

architecture SYN_ASYNCH_FD of FD_252 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1118 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1118);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_251 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_251;

architecture SYN_ASYNCH_FD of FD_251 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1119 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1119);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_250 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_250;

architecture SYN_ASYNCH_FD of FD_250 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1120 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1120);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_249 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_249;

architecture SYN_ASYNCH_FD of FD_249 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1121 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1121);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_248 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_248;

architecture SYN_ASYNCH_FD of FD_248 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1122 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1122);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_247 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_247;

architecture SYN_ASYNCH_FD of FD_247 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1123 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1123);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_246 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_246;

architecture SYN_ASYNCH_FD of FD_246 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1124 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1124);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_245 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_245;

architecture SYN_ASYNCH_FD of FD_245 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1125 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1125);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_244 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_244;

architecture SYN_ASYNCH_FD of FD_244 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1126 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1126);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_243 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_243;

architecture SYN_ASYNCH_FD of FD_243 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1127 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1127);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_242 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_242;

architecture SYN_ASYNCH_FD of FD_242 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1128 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1128);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_241 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_241;

architecture SYN_ASYNCH_FD of FD_241 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1129 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1129);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_240 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_240;

architecture SYN_ASYNCH_FD of FD_240 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1130 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1130);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_239 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_239;

architecture SYN_ASYNCH_FD of FD_239 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1131 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1131);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_238 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_238;

architecture SYN_ASYNCH_FD of FD_238 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1132 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1132);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_237 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_237;

architecture SYN_ASYNCH_FD of FD_237 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1133 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1133);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_236 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_236;

architecture SYN_ASYNCH_FD of FD_236 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1134 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1134);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_235 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_235;

architecture SYN_ASYNCH_FD of FD_235 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1135 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1135);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_234 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_234;

architecture SYN_ASYNCH_FD of FD_234 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1136 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1136);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_233 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_233;

architecture SYN_ASYNCH_FD of FD_233 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1137 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1137);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_232 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_232;

architecture SYN_ASYNCH_FD of FD_232 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1138 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1138);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_231 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_231;

architecture SYN_ASYNCH_FD of FD_231 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1139 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1139);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_230 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_230;

architecture SYN_ASYNCH_FD of FD_230 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1140 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1140);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_229 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_229;

architecture SYN_ASYNCH_FD of FD_229 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1141 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1141);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_228 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_228;

architecture SYN_ASYNCH_FD of FD_228 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1142 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1142);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_227 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_227;

architecture SYN_ASYNCH_FD of FD_227 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1143 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1143);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_226 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_226;

architecture SYN_ASYNCH_FD of FD_226 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1144 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1144);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_225 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_225;

architecture SYN_ASYNCH_FD of FD_225 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1145 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1145);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_224 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_224;

architecture SYN_ASYNCH_FD of FD_224 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1146 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1146);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_223 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_223;

architecture SYN_ASYNCH_FD of FD_223 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1147 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1147);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_222 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_222;

architecture SYN_ASYNCH_FD of FD_222 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1148 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1148);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_221 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_221;

architecture SYN_ASYNCH_FD of FD_221 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1149 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1149);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_220 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_220;

architecture SYN_ASYNCH_FD of FD_220 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1150 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1150);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_219 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_219;

architecture SYN_ASYNCH_FD of FD_219 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1151 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1151);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_218 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_218;

architecture SYN_ASYNCH_FD of FD_218 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1152 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1152);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_217 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_217;

architecture SYN_ASYNCH_FD of FD_217 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1153 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1153);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_216 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_216;

architecture SYN_ASYNCH_FD of FD_216 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1154 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1154);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_215 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_215;

architecture SYN_ASYNCH_FD of FD_215 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1155 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1155);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_214 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_214;

architecture SYN_ASYNCH_FD of FD_214 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1156 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1156);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_213 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_213;

architecture SYN_ASYNCH_FD of FD_213 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1157 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1157);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_212 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_212;

architecture SYN_ASYNCH_FD of FD_212 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1158 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1158);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_211 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_211;

architecture SYN_ASYNCH_FD of FD_211 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1159 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1159);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_210 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_210;

architecture SYN_ASYNCH_FD of FD_210 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1160 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1160);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_209 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_209;

architecture SYN_ASYNCH_FD of FD_209 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1161 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1161);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_208 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_208;

architecture SYN_ASYNCH_FD of FD_208 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1162 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1162);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_207 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_207;

architecture SYN_ASYNCH_FD of FD_207 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1163 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1163);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_206 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_206;

architecture SYN_ASYNCH_FD of FD_206 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1164 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1164);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_205 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_205;

architecture SYN_ASYNCH_FD of FD_205 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1165 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1165);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_204 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_204;

architecture SYN_ASYNCH_FD of FD_204 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1166 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1166);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_203 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_203;

architecture SYN_ASYNCH_FD of FD_203 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1167 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1167);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_202 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_202;

architecture SYN_ASYNCH_FD of FD_202 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1168 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1168);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_201 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_201;

architecture SYN_ASYNCH_FD of FD_201 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1169 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1169);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_200 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_200;

architecture SYN_ASYNCH_FD of FD_200 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1170 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1170);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_199 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_199;

architecture SYN_ASYNCH_FD of FD_199 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1171 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1171);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_198 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_198;

architecture SYN_ASYNCH_FD of FD_198 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1172 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1172);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_197 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_197;

architecture SYN_ASYNCH_FD of FD_197 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1173 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1173);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_196 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_196;

architecture SYN_ASYNCH_FD of FD_196 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1174 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1174);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_195 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_195;

architecture SYN_ASYNCH_FD of FD_195 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1175 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1175);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_194 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_194;

architecture SYN_ASYNCH_FD of FD_194 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1176 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1176);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_193 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_193;

architecture SYN_ASYNCH_FD of FD_193 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1177 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1177);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_192 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_192;

architecture SYN_ASYNCH_FD of FD_192 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1178 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1178);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_191 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_191;

architecture SYN_ASYNCH_FD of FD_191 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1179 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1179);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_190 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_190;

architecture SYN_ASYNCH_FD of FD_190 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1180 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1180);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_189 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_189;

architecture SYN_ASYNCH_FD of FD_189 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1181 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1181);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_188 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_188;

architecture SYN_ASYNCH_FD of FD_188 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1182 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1182);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_187 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_187;

architecture SYN_ASYNCH_FD of FD_187 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1183 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1183);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_186 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_186;

architecture SYN_ASYNCH_FD of FD_186 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1184 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1184);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_185 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_185;

architecture SYN_ASYNCH_FD of FD_185 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1185 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1185);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_184 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_184;

architecture SYN_ASYNCH_FD of FD_184 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1186 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1186);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_183 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_183;

architecture SYN_ASYNCH_FD of FD_183 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1187 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1187);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_182 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_182;

architecture SYN_ASYNCH_FD of FD_182 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1188 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1188);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_181 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_181;

architecture SYN_ASYNCH_FD of FD_181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1189 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1189);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_180 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_180;

architecture SYN_ASYNCH_FD of FD_180 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1190 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1190);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_179 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_179;

architecture SYN_ASYNCH_FD of FD_179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1191 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1191);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_178 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_178;

architecture SYN_ASYNCH_FD of FD_178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1192 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1192);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_177 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_177;

architecture SYN_ASYNCH_FD of FD_177 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1193 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1193);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_176 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_176;

architecture SYN_ASYNCH_FD of FD_176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1194 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1194);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_175 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_175;

architecture SYN_ASYNCH_FD of FD_175 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1195 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1195);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_174 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_174;

architecture SYN_ASYNCH_FD of FD_174 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1196 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1196);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_173 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_173;

architecture SYN_ASYNCH_FD of FD_173 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1197 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1197);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_172 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_172;

architecture SYN_ASYNCH_FD of FD_172 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1198 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1198);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_171 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_171;

architecture SYN_ASYNCH_FD of FD_171 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1199 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1199);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_170 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_170;

architecture SYN_ASYNCH_FD of FD_170 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1200 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1200);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_169 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_169;

architecture SYN_ASYNCH_FD of FD_169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1201 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1201);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_168 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_168;

architecture SYN_ASYNCH_FD of FD_168 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1202 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1202);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_167 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_167;

architecture SYN_ASYNCH_FD of FD_167 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1203 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1203);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_166 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_166;

architecture SYN_ASYNCH_FD of FD_166 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1204 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1204);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_165 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_165;

architecture SYN_ASYNCH_FD of FD_165 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1205 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1205);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_164 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_164;

architecture SYN_ASYNCH_FD of FD_164 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1206 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1206);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_163 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_163;

architecture SYN_ASYNCH_FD of FD_163 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1207 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1207);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_162 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_162;

architecture SYN_ASYNCH_FD of FD_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1208 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1208);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_161 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_161;

architecture SYN_ASYNCH_FD of FD_161 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1209 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1209);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_160 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_160;

architecture SYN_ASYNCH_FD of FD_160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1210 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1210);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_159 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_159;

architecture SYN_ASYNCH_FD of FD_159 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1211 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1211);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_158 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_158;

architecture SYN_ASYNCH_FD of FD_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1212 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1212);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_157 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_157;

architecture SYN_ASYNCH_FD of FD_157 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1213 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1213);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_156 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_156;

architecture SYN_ASYNCH_FD of FD_156 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1214 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1214);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_155 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_155;

architecture SYN_ASYNCH_FD of FD_155 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1215 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1215);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_154 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_154;

architecture SYN_ASYNCH_FD of FD_154 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1216 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1216);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_153 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_153;

architecture SYN_ASYNCH_FD of FD_153 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1217 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1217);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_152 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_152;

architecture SYN_ASYNCH_FD of FD_152 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1218 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1218);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_151 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_151;

architecture SYN_ASYNCH_FD of FD_151 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1219 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1219);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_150 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_150;

architecture SYN_ASYNCH_FD of FD_150 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1220 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1220);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_149 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_149;

architecture SYN_ASYNCH_FD of FD_149 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1221 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1221);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_148 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_148;

architecture SYN_ASYNCH_FD of FD_148 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1222 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1222);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_147 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_147;

architecture SYN_ASYNCH_FD of FD_147 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1223 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1223);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_146 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_146;

architecture SYN_ASYNCH_FD of FD_146 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1224 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1224);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_145 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_145;

architecture SYN_ASYNCH_FD of FD_145 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1225 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1225);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_144 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_144;

architecture SYN_ASYNCH_FD of FD_144 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1226 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1226);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_143 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_143;

architecture SYN_ASYNCH_FD of FD_143 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1227 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1227);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_142 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_142;

architecture SYN_ASYNCH_FD of FD_142 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1228 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1228);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_141 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_141;

architecture SYN_ASYNCH_FD of FD_141 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1229 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1229);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_140 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_140;

architecture SYN_ASYNCH_FD of FD_140 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1230 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1230);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_139 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_139;

architecture SYN_ASYNCH_FD of FD_139 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1231 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1231);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_138 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_138;

architecture SYN_ASYNCH_FD of FD_138 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1232 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1232);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_137 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_137;

architecture SYN_ASYNCH_FD of FD_137 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1233 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1233);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_136 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_136;

architecture SYN_ASYNCH_FD of FD_136 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1234 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1234);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_135 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_135;

architecture SYN_ASYNCH_FD of FD_135 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1235 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1235);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_134 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_134;

architecture SYN_ASYNCH_FD of FD_134 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1236 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1236);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_133 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_133;

architecture SYN_ASYNCH_FD of FD_133 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1237 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1237);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_132 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_132;

architecture SYN_ASYNCH_FD of FD_132 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1238 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1238);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_131 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_131;

architecture SYN_ASYNCH_FD of FD_131 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1239 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1239);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_130 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_130;

architecture SYN_ASYNCH_FD of FD_130 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1240 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1240);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_129 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_129;

architecture SYN_ASYNCH_FD of FD_129 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1241 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1241);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_128 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_128;

architecture SYN_ASYNCH_FD of FD_128 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1242 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1242);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_127 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_127;

architecture SYN_ASYNCH_FD of FD_127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1243 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1243);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_126 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_126;

architecture SYN_ASYNCH_FD of FD_126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1244 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1244);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_125 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_125;

architecture SYN_ASYNCH_FD of FD_125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1245 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1245);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_124 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_124;

architecture SYN_ASYNCH_FD of FD_124 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1246 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1246);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_123 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_123;

architecture SYN_ASYNCH_FD of FD_123 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1247 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1247);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_122 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_122;

architecture SYN_ASYNCH_FD of FD_122 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1248 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1248);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_121 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_121;

architecture SYN_ASYNCH_FD of FD_121 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1249 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1249);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_120 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_120;

architecture SYN_ASYNCH_FD of FD_120 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1250 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1250);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_119 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_119;

architecture SYN_ASYNCH_FD of FD_119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1251 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1251);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_118 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_118;

architecture SYN_ASYNCH_FD of FD_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1252 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1252);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_117 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_117;

architecture SYN_ASYNCH_FD of FD_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1253 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1253);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_116 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_116;

architecture SYN_ASYNCH_FD of FD_116 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1254 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1254);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_115 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_115;

architecture SYN_ASYNCH_FD of FD_115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1255 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1255);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_114 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_114;

architecture SYN_ASYNCH_FD of FD_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1256 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1256);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_113 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_113;

architecture SYN_ASYNCH_FD of FD_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1257 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1257);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_112 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_112;

architecture SYN_ASYNCH_FD of FD_112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1258 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1258);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_111 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_111;

architecture SYN_ASYNCH_FD of FD_111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1259 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1259);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_110 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_110;

architecture SYN_ASYNCH_FD of FD_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1260 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1260);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_109 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_109;

architecture SYN_ASYNCH_FD of FD_109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1261 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1261);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_108 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_108;

architecture SYN_ASYNCH_FD of FD_108 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1262 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1262);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_107 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_107;

architecture SYN_ASYNCH_FD of FD_107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1263 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1263);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_106 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_106;

architecture SYN_ASYNCH_FD of FD_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1264 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1264);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_105 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_105;

architecture SYN_ASYNCH_FD of FD_105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1265 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1265);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_104 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_104;

architecture SYN_ASYNCH_FD of FD_104 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1266 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1266);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_103 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_103;

architecture SYN_ASYNCH_FD of FD_103 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1267 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1267);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_102 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_102;

architecture SYN_ASYNCH_FD of FD_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1268 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1268);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_101 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_101;

architecture SYN_ASYNCH_FD of FD_101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1269 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1269);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_100 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_100;

architecture SYN_ASYNCH_FD of FD_100 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1270 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1270);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_99 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_99;

architecture SYN_ASYNCH_FD of FD_99 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1271 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1271);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_98 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_98;

architecture SYN_ASYNCH_FD of FD_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1272 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1272);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_97 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_97;

architecture SYN_ASYNCH_FD of FD_97 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1273 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1273);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_96 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_96;

architecture SYN_ASYNCH_FD of FD_96 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1274 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1274);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_95 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_95;

architecture SYN_ASYNCH_FD of FD_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1275 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1275);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_94 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_94;

architecture SYN_ASYNCH_FD of FD_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1276 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1276);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_93 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_93;

architecture SYN_ASYNCH_FD of FD_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1277 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1277);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_92 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_92;

architecture SYN_ASYNCH_FD of FD_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1278 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1278);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_91 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_91;

architecture SYN_ASYNCH_FD of FD_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1279 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1279);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_90 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_90;

architecture SYN_ASYNCH_FD of FD_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1280 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1280);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_89 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_89;

architecture SYN_ASYNCH_FD of FD_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1281 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1281);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_88 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_88;

architecture SYN_ASYNCH_FD of FD_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1282 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1282);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_87 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_87;

architecture SYN_ASYNCH_FD of FD_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1283 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1283);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_86 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_86;

architecture SYN_ASYNCH_FD of FD_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1284 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1284);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_85 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_85;

architecture SYN_ASYNCH_FD of FD_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1285 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1285);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_84 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_84;

architecture SYN_ASYNCH_FD of FD_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1286 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1286);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_83 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_83;

architecture SYN_ASYNCH_FD of FD_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1287 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1287);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_82 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_82;

architecture SYN_ASYNCH_FD of FD_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1288 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1288);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_81 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_81;

architecture SYN_ASYNCH_FD of FD_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1289 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1289);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_80 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_80;

architecture SYN_ASYNCH_FD of FD_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1290 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1290);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_79 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_79;

architecture SYN_ASYNCH_FD of FD_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1291 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1291);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_78 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_78;

architecture SYN_ASYNCH_FD of FD_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1292 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1292);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_77 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_77;

architecture SYN_ASYNCH_FD of FD_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1293 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1293);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_76 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_76;

architecture SYN_ASYNCH_FD of FD_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1294 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1294);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_75 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_75;

architecture SYN_ASYNCH_FD of FD_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1295 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1295);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_74 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_74;

architecture SYN_ASYNCH_FD of FD_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1296 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1296);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_73 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_73;

architecture SYN_ASYNCH_FD of FD_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1297 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1297);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_72 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_72;

architecture SYN_ASYNCH_FD of FD_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1298 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1298);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_71 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_71;

architecture SYN_ASYNCH_FD of FD_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1299 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1299);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_70 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_70;

architecture SYN_ASYNCH_FD of FD_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1300 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1300);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_69 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_69;

architecture SYN_ASYNCH_FD of FD_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1301 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1301);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_68 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_68;

architecture SYN_ASYNCH_FD of FD_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1302 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1302);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_67 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_67;

architecture SYN_ASYNCH_FD of FD_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1303 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1303);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_66 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_66;

architecture SYN_ASYNCH_FD of FD_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1304 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1304);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_65 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_65;

architecture SYN_ASYNCH_FD of FD_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1305 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1305);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_64 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_64;

architecture SYN_ASYNCH_FD of FD_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1306 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1306);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_63 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_63;

architecture SYN_ASYNCH_FD of FD_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1307 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1307);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_62 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_62;

architecture SYN_ASYNCH_FD of FD_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1308 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1308);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_61 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_61;

architecture SYN_ASYNCH_FD of FD_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1309 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1309);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_60 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_60;

architecture SYN_ASYNCH_FD of FD_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1310 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1310);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_59 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_59;

architecture SYN_ASYNCH_FD of FD_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1311 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1311);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_58 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_58;

architecture SYN_ASYNCH_FD of FD_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1312 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1312);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_57 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_57;

architecture SYN_ASYNCH_FD of FD_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1313 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1313);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_56 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_56;

architecture SYN_ASYNCH_FD of FD_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1314 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1314);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_55 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_55;

architecture SYN_ASYNCH_FD of FD_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1315 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1315);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_54 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_54;

architecture SYN_ASYNCH_FD of FD_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1316 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1316);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_53 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_53;

architecture SYN_ASYNCH_FD of FD_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1317 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1317);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_52 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_52;

architecture SYN_ASYNCH_FD of FD_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1318 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1318);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_51 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_51;

architecture SYN_ASYNCH_FD of FD_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1319 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1319);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_50 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_50;

architecture SYN_ASYNCH_FD of FD_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1320 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1320);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_49 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_49;

architecture SYN_ASYNCH_FD of FD_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1321 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1321);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_48 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_48;

architecture SYN_ASYNCH_FD of FD_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1322 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1322);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_47 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_47;

architecture SYN_ASYNCH_FD of FD_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1323 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1323);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_46 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_46;

architecture SYN_ASYNCH_FD of FD_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1324 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1324);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_45 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_45;

architecture SYN_ASYNCH_FD of FD_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1325 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1325);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_44 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_44;

architecture SYN_ASYNCH_FD of FD_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1326 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1326);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_43 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_43;

architecture SYN_ASYNCH_FD of FD_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1327 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1327);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_42 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_42;

architecture SYN_ASYNCH_FD of FD_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1328 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1328);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_41 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_41;

architecture SYN_ASYNCH_FD of FD_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1329 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1329);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_40 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_40;

architecture SYN_ASYNCH_FD of FD_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1330 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1330);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_39 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_39;

architecture SYN_ASYNCH_FD of FD_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1331 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1331);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_38 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_38;

architecture SYN_ASYNCH_FD of FD_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1332 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1332);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_37 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_37;

architecture SYN_ASYNCH_FD of FD_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1333 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1333);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_36 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_36;

architecture SYN_ASYNCH_FD of FD_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1334 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1334);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_35 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_35;

architecture SYN_ASYNCH_FD of FD_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1335 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1335);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_34 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_34;

architecture SYN_ASYNCH_FD of FD_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1336 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1336);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_33 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_33;

architecture SYN_ASYNCH_FD of FD_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1337 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1337);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_32 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_32;

architecture SYN_ASYNCH_FD of FD_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1338 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1338);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_31 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_31;

architecture SYN_ASYNCH_FD of FD_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1339 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1339);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_30 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_30;

architecture SYN_ASYNCH_FD of FD_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1340 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1340);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_29 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_29;

architecture SYN_ASYNCH_FD of FD_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1341 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1341);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_28 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_28;

architecture SYN_ASYNCH_FD of FD_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1342 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1342);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_27 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_27;

architecture SYN_ASYNCH_FD of FD_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1343 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1343);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_26 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_26;

architecture SYN_ASYNCH_FD of FD_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1344 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1344);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_25 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_25;

architecture SYN_ASYNCH_FD of FD_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1345 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1345);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_24 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_24;

architecture SYN_ASYNCH_FD of FD_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1346 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1346);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_23 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_23;

architecture SYN_ASYNCH_FD of FD_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1347 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1347);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_22 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_22;

architecture SYN_ASYNCH_FD of FD_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1348 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1348);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_21 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_21;

architecture SYN_ASYNCH_FD of FD_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1349 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1349);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_20 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_20;

architecture SYN_ASYNCH_FD of FD_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1350 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1350);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_19 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_19;

architecture SYN_ASYNCH_FD of FD_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1351 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1351);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_18 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_18;

architecture SYN_ASYNCH_FD of FD_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1352 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1352);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_17 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_17;

architecture SYN_ASYNCH_FD of FD_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1353 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1353);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_16 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_16;

architecture SYN_ASYNCH_FD of FD_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1354 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1354);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_15 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_15;

architecture SYN_ASYNCH_FD of FD_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1355 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1355);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_14 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_14;

architecture SYN_ASYNCH_FD of FD_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1356 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1356);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_13 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_13;

architecture SYN_ASYNCH_FD of FD_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1357 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1357);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_12 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_12;

architecture SYN_ASYNCH_FD of FD_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1358 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1358);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_11 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_11;

architecture SYN_ASYNCH_FD of FD_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1359 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1359);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_10 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_10;

architecture SYN_ASYNCH_FD of FD_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1360 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1360);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_9 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_9;

architecture SYN_ASYNCH_FD of FD_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1361 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1361);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_8 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_8;

architecture SYN_ASYNCH_FD of FD_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1362 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1362);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_7 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_7;

architecture SYN_ASYNCH_FD of FD_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1363 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1363);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_6 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_6;

architecture SYN_ASYNCH_FD of FD_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1364 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1364);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_5 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_5;

architecture SYN_ASYNCH_FD of FD_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1365 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1365);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_4 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_4;

architecture SYN_ASYNCH_FD of FD_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1366 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1366);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_3 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_3;

architecture SYN_ASYNCH_FD of FD_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1367 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1367);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_2 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_2;

architecture SYN_ASYNCH_FD of FD_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1368 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1368);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_1 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_1;

architecture SYN_ASYNCH_FD of FD_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1369 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1369);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_3;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U5 : MUX2_X1 port map( A => B(4), B => A(4), S => S, Z => Y(4));
   U6 : MUX2_X1 port map( A => B(5), B => A(5), S => S, Z => Y(5));
   U7 : MUX2_X1 port map( A => B(6), B => A(6), S => S, Z => Y(6));
   U8 : MUX2_X1 port map( A => B(7), B => A(7), S => S, Z => Y(7));
   U9 : MUX2_X1 port map( A => B(8), B => A(8), S => S, Z => Y(8));
   U10 : MUX2_X1 port map( A => B(9), B => A(9), S => S, Z => Y(9));
   U11 : MUX2_X1 port map( A => B(10), B => A(10), S => S, Z => Y(10));
   U12 : MUX2_X1 port map( A => B(11), B => A(11), S => S, Z => Y(11));
   U13 : MUX2_X1 port map( A => B(12), B => A(12), S => S, Z => Y(12));
   U14 : MUX2_X1 port map( A => B(13), B => A(13), S => S, Z => Y(13));
   U15 : MUX2_X1 port map( A => B(14), B => A(14), S => S, Z => Y(14));
   U16 : MUX2_X1 port map( A => B(15), B => A(15), S => S, Z => Y(15));
   U17 : MUX2_X1 port map( A => B(16), B => A(16), S => S, Z => Y(16));
   U18 : MUX2_X1 port map( A => B(17), B => A(17), S => S, Z => Y(17));
   U19 : MUX2_X1 port map( A => B(18), B => A(18), S => S, Z => Y(18));
   U20 : MUX2_X1 port map( A => B(19), B => A(19), S => S, Z => Y(19));
   U21 : MUX2_X1 port map( A => B(20), B => A(20), S => S, Z => Y(20));
   U22 : MUX2_X1 port map( A => B(21), B => A(21), S => S, Z => Y(21));
   U23 : MUX2_X1 port map( A => B(22), B => A(22), S => S, Z => Y(22));
   U24 : MUX2_X1 port map( A => B(23), B => A(23), S => S, Z => Y(23));
   U25 : MUX2_X1 port map( A => B(24), B => A(24), S => S, Z => Y(24));
   U26 : MUX2_X1 port map( A => B(25), B => A(25), S => S, Z => Y(25));
   U27 : MUX2_X1 port map( A => B(26), B => A(26), S => S, Z => Y(26));
   U28 : MUX2_X1 port map( A => B(27), B => A(27), S => S, Z => Y(27));
   U29 : MUX2_X1 port map( A => B(28), B => A(28), S => S, Z => Y(28));
   U30 : MUX2_X1 port map( A => B(29), B => A(29), S => S, Z => Y(29));
   U31 : MUX2_X1 port map( A => B(30), B => A(30), S => S, Z => Y(30));
   U32 : MUX2_X1 port map( A => B(31), B => A(31), S => S, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_2;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(31), B => A(31), S => S, Z => Y(31));
   U2 : MUX2_X1 port map( A => B(30), B => A(30), S => S, Z => Y(30));
   U3 : MUX2_X1 port map( A => B(29), B => A(29), S => S, Z => Y(29));
   U4 : MUX2_X1 port map( A => B(28), B => A(28), S => S, Z => Y(28));
   U5 : MUX2_X1 port map( A => B(27), B => A(27), S => S, Z => Y(27));
   U6 : MUX2_X1 port map( A => B(26), B => A(26), S => S, Z => Y(26));
   U7 : MUX2_X1 port map( A => B(25), B => A(25), S => S, Z => Y(25));
   U8 : MUX2_X1 port map( A => B(24), B => A(24), S => S, Z => Y(24));
   U9 : MUX2_X1 port map( A => B(23), B => A(23), S => S, Z => Y(23));
   U10 : MUX2_X1 port map( A => B(22), B => A(22), S => S, Z => Y(22));
   U11 : MUX2_X1 port map( A => B(21), B => A(21), S => S, Z => Y(21));
   U12 : MUX2_X1 port map( A => B(20), B => A(20), S => S, Z => Y(20));
   U13 : MUX2_X1 port map( A => B(19), B => A(19), S => S, Z => Y(19));
   U14 : MUX2_X1 port map( A => B(18), B => A(18), S => S, Z => Y(18));
   U15 : MUX2_X1 port map( A => B(17), B => A(17), S => S, Z => Y(17));
   U16 : MUX2_X1 port map( A => B(16), B => A(16), S => S, Z => Y(16));
   U17 : MUX2_X1 port map( A => B(15), B => A(15), S => S, Z => Y(15));
   U18 : MUX2_X1 port map( A => B(14), B => A(14), S => S, Z => Y(14));
   U19 : MUX2_X1 port map( A => B(13), B => A(13), S => S, Z => Y(13));
   U20 : MUX2_X1 port map( A => B(12), B => A(12), S => S, Z => Y(12));
   U21 : MUX2_X1 port map( A => B(11), B => A(11), S => S, Z => Y(11));
   U22 : MUX2_X1 port map( A => B(10), B => A(10), S => S, Z => Y(10));
   U23 : MUX2_X1 port map( A => B(9), B => A(9), S => S, Z => Y(9));
   U24 : MUX2_X1 port map( A => B(8), B => A(8), S => S, Z => Y(8));
   U25 : MUX2_X1 port map( A => B(7), B => A(7), S => S, Z => Y(7));
   U26 : MUX2_X1 port map( A => B(6), B => A(6), S => S, Z => Y(6));
   U27 : MUX2_X1 port map( A => B(5), B => A(5), S => S, Z => Y(5));
   U28 : MUX2_X1 port map( A => B(4), B => A(4), S => S, Z => Y(4));
   U29 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U30 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U31 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U32 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_1;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U5 : MUX2_X1 port map( A => B(4), B => A(4), S => S, Z => Y(4));
   U6 : MUX2_X1 port map( A => B(5), B => A(5), S => S, Z => Y(5));
   U7 : MUX2_X1 port map( A => B(6), B => A(6), S => S, Z => Y(6));
   U8 : MUX2_X1 port map( A => B(7), B => A(7), S => S, Z => Y(7));
   U9 : MUX2_X1 port map( A => B(8), B => A(8), S => S, Z => Y(8));
   U10 : MUX2_X1 port map( A => B(9), B => A(9), S => S, Z => Y(9));
   U11 : MUX2_X1 port map( A => B(10), B => A(10), S => S, Z => Y(10));
   U12 : MUX2_X1 port map( A => B(11), B => A(11), S => S, Z => Y(11));
   U13 : MUX2_X1 port map( A => B(12), B => A(12), S => S, Z => Y(12));
   U14 : MUX2_X1 port map( A => B(13), B => A(13), S => S, Z => Y(13));
   U15 : MUX2_X1 port map( A => B(14), B => A(14), S => S, Z => Y(14));
   U16 : MUX2_X1 port map( A => B(15), B => A(15), S => S, Z => Y(15));
   U17 : MUX2_X1 port map( A => B(16), B => A(16), S => S, Z => Y(16));
   U18 : MUX2_X1 port map( A => B(17), B => A(17), S => S, Z => Y(17));
   U19 : MUX2_X1 port map( A => B(18), B => A(18), S => S, Z => Y(18));
   U20 : MUX2_X1 port map( A => B(19), B => A(19), S => S, Z => Y(19));
   U21 : MUX2_X1 port map( A => B(20), B => A(20), S => S, Z => Y(20));
   U22 : MUX2_X1 port map( A => B(21), B => A(21), S => S, Z => Y(21));
   U23 : MUX2_X1 port map( A => B(22), B => A(22), S => S, Z => Y(22));
   U24 : MUX2_X1 port map( A => B(23), B => A(23), S => S, Z => Y(23));
   U25 : MUX2_X1 port map( A => B(24), B => A(24), S => S, Z => Y(24));
   U26 : MUX2_X1 port map( A => B(25), B => A(25), S => S, Z => Y(25));
   U27 : MUX2_X1 port map( A => B(26), B => A(26), S => S, Z => Y(26));
   U28 : MUX2_X1 port map( A => B(27), B => A(27), S => S, Z => Y(27));
   U29 : MUX2_X1 port map( A => B(28), B => A(28), S => S, Z => Y(28));
   U30 : MUX2_X1 port map( A => B(29), B => A(29), S => S, Z => Y(29));
   U31 : MUX2_X1 port map( A => B(30), B => A(30), S => S, Z => Y(30));
   U32 : MUX2_X1 port map( A => B(31), B => A(31), S => S, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_10 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_10;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_10 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_289
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_290
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_291
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_292
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_293
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_294
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_295
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_296
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_297
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_298
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_299
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_300
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_301
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_302
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_303
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_304
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_305
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_306
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_307
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_308
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_309
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_310
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_311
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_312
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_313
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_314
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_315
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_316
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_317
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_318
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_319
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_320
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FF_0 : FD_320 port map( D => data_in(0), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_319 port map( D => data_in(1), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_318 port map( D => data_in(2), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_317 port map( D => data_in(3), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_316 port map( D => data_in(4), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_315 port map( D => data_in(5), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_314 port map( D => data_in(6), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_313 port map( D => data_in(7), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_312 port map( D => data_in(8), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_311 port map( D => data_in(9), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_310 port map( D => data_in(10), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_309 port map( D => data_in(11), CK => n6, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_308 port map( D => data_in(12), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_307 port map( D => data_in(13), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_306 port map( D => data_in(14), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_305 port map( D => data_in(15), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_304 port map( D => data_in(16), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_303 port map( D => data_in(17), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_302 port map( D => data_in(18), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_301 port map( D => data_in(19), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_300 port map( D => data_in(20), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_299 port map( D => data_in(21), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_298 port map( D => data_in(22), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_297 port map( D => data_in(23), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_296 port map( D => data_in(24), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_295 port map( D => data_in(25), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_294 port map( D => data_in(26), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_293 port map( D => data_in(27), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_292 port map( D => data_in(28), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_291 port map( D => data_in(29), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_290 port map( D => data_in(30), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_289 port map( D => data_in(31), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n4);
   U2 : BUF_X1 port map( A => CK, Z => n8);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_9 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_9;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_9 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_257
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_258
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_259
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_260
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_261
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_262
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_263
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_264
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_265
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_266
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_267
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_268
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_269
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_270
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_271
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_272
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_273
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_274
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_275
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_276
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_277
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_278
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_279
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_280
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_281
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_282
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_283
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_284
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_285
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_286
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_287
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_288
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FF_0 : FD_288 port map( D => data_in(0), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_287 port map( D => data_in(1), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_286 port map( D => data_in(2), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_285 port map( D => data_in(3), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_284 port map( D => data_in(4), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_283 port map( D => data_in(5), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_282 port map( D => data_in(6), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_281 port map( D => data_in(7), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_280 port map( D => data_in(8), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_279 port map( D => data_in(9), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_278 port map( D => data_in(10), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_277 port map( D => data_in(11), CK => n6, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_276 port map( D => data_in(12), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_275 port map( D => data_in(13), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_274 port map( D => data_in(14), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_273 port map( D => data_in(15), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_272 port map( D => data_in(16), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_271 port map( D => data_in(17), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_270 port map( D => data_in(18), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_269 port map( D => data_in(19), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_268 port map( D => data_in(20), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_267 port map( D => data_in(21), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_266 port map( D => data_in(22), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_265 port map( D => data_in(23), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_264 port map( D => data_in(24), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_263 port map( D => data_in(25), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_262 port map( D => data_in(26), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_261 port map( D => data_in(27), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_260 port map( D => data_in(28), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_259 port map( D => data_in(29), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_258 port map( D => data_in(30), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_257 port map( D => data_in(31), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n4);
   U2 : BUF_X1 port map( A => CK, Z => n8);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_8 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_8;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_8 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_225
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_226
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_227
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_228
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_229
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_230
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_231
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_232
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_233
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_234
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_235
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_236
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_237
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_238
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_239
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_240
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_241
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_242
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_243
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_244
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_245
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_246
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_247
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_248
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_249
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_250
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_251
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_252
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_253
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_254
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_255
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_256
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FF_0 : FD_256 port map( D => data_in(0), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_255 port map( D => data_in(1), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_254 port map( D => data_in(2), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_253 port map( D => data_in(3), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_252 port map( D => data_in(4), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_251 port map( D => data_in(5), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_250 port map( D => data_in(6), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_249 port map( D => data_in(7), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_248 port map( D => data_in(8), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_247 port map( D => data_in(9), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_246 port map( D => data_in(10), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_245 port map( D => data_in(11), CK => n6, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_244 port map( D => data_in(12), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_243 port map( D => data_in(13), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_242 port map( D => data_in(14), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_241 port map( D => data_in(15), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_240 port map( D => data_in(16), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_239 port map( D => data_in(17), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_238 port map( D => data_in(18), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_237 port map( D => data_in(19), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_236 port map( D => data_in(20), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_235 port map( D => data_in(21), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_234 port map( D => data_in(22), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_233 port map( D => data_in(23), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_232 port map( D => data_in(24), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_231 port map( D => data_in(25), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_230 port map( D => data_in(26), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_229 port map( D => data_in(27), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_228 port map( D => data_in(28), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_227 port map( D => data_in(29), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_226 port map( D => data_in(30), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_225 port map( D => data_in(31), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => CK, Z => n8);
   U2 : BUF_X1 port map( A => RESET, Z => n4);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_7 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_7;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_7 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_193
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_194
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_195
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_196
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_197
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_198
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_199
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_200
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_201
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_202
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_203
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_204
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_205
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_206
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_207
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_208
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_209
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_210
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_211
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_212
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_213
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_214
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_215
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_216
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_217
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_218
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_219
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_220
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_221
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_222
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_223
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_224
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FF_0 : FD_224 port map( D => data_in(0), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_223 port map( D => data_in(1), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_222 port map( D => data_in(2), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_221 port map( D => data_in(3), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_220 port map( D => data_in(4), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_219 port map( D => data_in(5), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_218 port map( D => data_in(6), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_217 port map( D => data_in(7), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_216 port map( D => data_in(8), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_215 port map( D => data_in(9), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_214 port map( D => data_in(10), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_213 port map( D => data_in(11), CK => n6, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_212 port map( D => data_in(12), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_211 port map( D => data_in(13), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_210 port map( D => data_in(14), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_209 port map( D => data_in(15), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_208 port map( D => data_in(16), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_207 port map( D => data_in(17), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_206 port map( D => data_in(18), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_205 port map( D => data_in(19), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_204 port map( D => data_in(20), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_203 port map( D => data_in(21), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_202 port map( D => data_in(22), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_201 port map( D => data_in(23), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_200 port map( D => data_in(24), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_199 port map( D => data_in(25), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_198 port map( D => data_in(26), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_197 port map( D => data_in(27), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_196 port map( D => data_in(28), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_195 port map( D => data_in(29), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_194 port map( D => data_in(30), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_193 port map( D => data_in(31), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => CK, Z => n8);
   U2 : BUF_X1 port map( A => RESET, Z => n4);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_6 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_6;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_161
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_162
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_163
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_164
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_165
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_166
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_167
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_168
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_169
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_170
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_171
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_172
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_173
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_174
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_175
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_176
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_177
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_178
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_179
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_180
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_181
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_182
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_183
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_184
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_185
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_186
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_187
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_188
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_189
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_190
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_191
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_192
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FF_0 : FD_192 port map( D => data_in(0), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_191 port map( D => data_in(1), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_190 port map( D => data_in(2), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_189 port map( D => data_in(3), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_188 port map( D => data_in(4), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_187 port map( D => data_in(5), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_186 port map( D => data_in(6), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_185 port map( D => data_in(7), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_184 port map( D => data_in(8), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_183 port map( D => data_in(9), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_182 port map( D => data_in(10), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_181 port map( D => data_in(11), CK => n6, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_180 port map( D => data_in(12), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_179 port map( D => data_in(13), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_178 port map( D => data_in(14), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_177 port map( D => data_in(15), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_176 port map( D => data_in(16), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_175 port map( D => data_in(17), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_174 port map( D => data_in(18), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_173 port map( D => data_in(19), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_172 port map( D => data_in(20), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_171 port map( D => data_in(21), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_170 port map( D => data_in(22), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_169 port map( D => data_in(23), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_168 port map( D => data_in(24), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_167 port map( D => data_in(25), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_166 port map( D => data_in(26), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_165 port map( D => data_in(27), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_164 port map( D => data_in(28), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_163 port map( D => data_in(29), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_162 port map( D => data_in(30), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_161 port map( D => data_in(31), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => CK, Z => n8);
   U2 : BUF_X1 port map( A => RESET, Z => n4);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_5 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_5;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_129
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_130
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_131
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_132
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_133
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_134
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_135
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_136
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_137
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_138
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_139
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_140
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_141
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_142
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_143
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_144
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_145
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_146
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_147
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_148
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_149
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_150
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_151
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_152
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_153
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_154
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_155
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_156
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_157
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_158
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_159
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_160
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FF_0 : FD_160 port map( D => data_in(0), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_159 port map( D => data_in(1), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_158 port map( D => data_in(2), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_157 port map( D => data_in(3), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_156 port map( D => data_in(4), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_155 port map( D => data_in(5), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_154 port map( D => data_in(6), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_153 port map( D => data_in(7), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_152 port map( D => data_in(8), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_151 port map( D => data_in(9), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_150 port map( D => data_in(10), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_149 port map( D => data_in(11), CK => n6, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_148 port map( D => data_in(12), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_147 port map( D => data_in(13), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_146 port map( D => data_in(14), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_145 port map( D => data_in(15), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_144 port map( D => data_in(16), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_143 port map( D => data_in(17), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_142 port map( D => data_in(18), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_141 port map( D => data_in(19), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_140 port map( D => data_in(20), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_139 port map( D => data_in(21), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_138 port map( D => data_in(22), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_137 port map( D => data_in(23), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_136 port map( D => data_in(24), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_135 port map( D => data_in(25), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_134 port map( D => data_in(26), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_133 port map( D => data_in(27), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_132 port map( D => data_in(28), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_131 port map( D => data_in(29), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_130 port map( D => data_in(30), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_129 port map( D => data_in(31), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n4);
   U2 : BUF_X1 port map( A => CK, Z => n8);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_4 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_4;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_97
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_98
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_99
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_100
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_101
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_102
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_103
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_104
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_105
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_106
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_107
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_108
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_109
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_110
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_111
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_112
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_113
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_114
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_115
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_116
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_117
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_118
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_119
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_120
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_121
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_122
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_123
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_124
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_125
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_126
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_127
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_128
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FF_0 : FD_128 port map( D => data_in(0), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_127 port map( D => data_in(1), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_126 port map( D => data_in(2), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_125 port map( D => data_in(3), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_124 port map( D => data_in(4), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_123 port map( D => data_in(5), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_122 port map( D => data_in(6), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_121 port map( D => data_in(7), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_120 port map( D => data_in(8), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_119 port map( D => data_in(9), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_118 port map( D => data_in(10), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_117 port map( D => data_in(11), CK => n6, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_116 port map( D => data_in(12), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_115 port map( D => data_in(13), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_114 port map( D => data_in(14), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_113 port map( D => data_in(15), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_112 port map( D => data_in(16), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_111 port map( D => data_in(17), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_110 port map( D => data_in(18), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_109 port map( D => data_in(19), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_108 port map( D => data_in(20), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_107 port map( D => data_in(21), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_106 port map( D => data_in(22), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_105 port map( D => data_in(23), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_104 port map( D => data_in(24), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_103 port map( D => data_in(25), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_102 port map( D => data_in(26), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_101 port map( D => data_in(27), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_100 port map( D => data_in(28), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_99 port map( D => data_in(29), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_98 port map( D => data_in(30), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_97 port map( D => data_in(31), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n4);
   U2 : BUF_X1 port map( A => CK, Z => n8);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_3 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_3;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_65
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_66
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_67
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_68
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_69
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_70
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_71
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_72
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_73
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_74
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_75
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_76
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_77
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_78
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_79
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_80
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_81
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_82
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_83
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_84
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_85
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_86
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_87
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_88
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_89
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_90
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_91
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_92
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_93
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_94
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_95
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_96
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FF_0 : FD_96 port map( D => data_in(0), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_95 port map( D => data_in(1), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_94 port map( D => data_in(2), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_93 port map( D => data_in(3), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_92 port map( D => data_in(4), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_91 port map( D => data_in(5), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_90 port map( D => data_in(6), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_89 port map( D => data_in(7), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_88 port map( D => data_in(8), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_87 port map( D => data_in(9), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_86 port map( D => data_in(10), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_85 port map( D => data_in(11), CK => n6, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_84 port map( D => data_in(12), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_83 port map( D => data_in(13), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_82 port map( D => data_in(14), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_81 port map( D => data_in(15), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_80 port map( D => data_in(16), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_79 port map( D => data_in(17), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_78 port map( D => data_in(18), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_77 port map( D => data_in(19), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_76 port map( D => data_in(20), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_75 port map( D => data_in(21), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_74 port map( D => data_in(22), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_73 port map( D => data_in(23), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_72 port map( D => data_in(24), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_71 port map( D => data_in(25), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_70 port map( D => data_in(26), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_69 port map( D => data_in(27), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_68 port map( D => data_in(28), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_67 port map( D => data_in(29), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_66 port map( D => data_in(30), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_65 port map( D => data_in(31), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n4);
   U2 : BUF_X1 port map( A => CK, Z => n8);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_2 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_2;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_33
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_34
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_35
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_36
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_37
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_38
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_39
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_40
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_41
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_42
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_43
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_44
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_45
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_46
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_47
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_48
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_49
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_50
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_51
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_52
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_53
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_54
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_55
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_56
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_57
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_58
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_59
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_60
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_61
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_62
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_63
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_64
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FF_0 : FD_64 port map( D => data_in(0), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_63 port map( D => data_in(1), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_62 port map( D => data_in(2), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_61 port map( D => data_in(3), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_60 port map( D => data_in(4), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_59 port map( D => data_in(5), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_58 port map( D => data_in(6), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_57 port map( D => data_in(7), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_56 port map( D => data_in(8), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_55 port map( D => data_in(9), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_54 port map( D => data_in(10), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_53 port map( D => data_in(11), CK => n6, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_52 port map( D => data_in(12), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_51 port map( D => data_in(13), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_50 port map( D => data_in(14), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_49 port map( D => data_in(15), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_48 port map( D => data_in(16), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_47 port map( D => data_in(17), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_46 port map( D => data_in(18), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_45 port map( D => data_in(19), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_44 port map( D => data_in(20), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_43 port map( D => data_in(21), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_42 port map( D => data_in(22), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_41 port map( D => data_in(23), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_40 port map( D => data_in(24), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_39 port map( D => data_in(25), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_38 port map( D => data_in(26), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_37 port map( D => data_in(27), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_36 port map( D => data_in(28), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_35 port map( D => data_in(29), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_34 port map( D => data_in(30), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_33 port map( D => data_in(31), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n4);
   U2 : BUF_X1 port map( A => CK, Z => n8);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_1 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_1;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_3
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_4
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_5
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_6
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_7
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_8
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_9
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_10
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_11
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_12
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_13
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_14
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_15
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_16
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_17
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_18
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_19
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_20
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_21
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_22
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_23
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_24
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_25
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_26
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_27
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_28
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_29
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_30
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_31
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_32
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FF_0 : FD_32 port map( D => data_in(0), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_31 port map( D => data_in(1), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_30 port map( D => data_in(2), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_29 port map( D => data_in(3), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_28 port map( D => data_in(4), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_27 port map( D => data_in(5), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_26 port map( D => data_in(6), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_25 port map( D => data_in(7), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_24 port map( D => data_in(8), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_23 port map( D => data_in(9), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_22 port map( D => data_in(10), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_21 port map( D => data_in(11), CK => n6, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_20 port map( D => data_in(12), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_19 port map( D => data_in(13), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_18 port map( D => data_in(14), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_17 port map( D => data_in(15), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_16 port map( D => data_in(16), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_15 port map( D => data_in(17), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_14 port map( D => data_in(18), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_13 port map( D => data_in(19), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_12 port map( D => data_in(20), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_11 port map( D => data_in(21), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_10 port map( D => data_in(22), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_9 port map( D => data_in(23), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_8 port map( D => data_in(24), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_7 port map( D => data_in(25), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_6 port map( D => data_in(26), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_5 port map( D => data_in(27), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_4 port map( D => data_in(28), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_3 port map( D => data_in(29), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_2 port map( D => data_in(30), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_1 port map( D => data_in(31), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n4);
   U2 : BUF_X1 port map( A => CK, Z => n8);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_0;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_0;

architecture SYN_BEHAVIORAL of RCA_NBITS4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(3));
   U3 : XOR2_X1 port map( A => n3, B => A(3), Z => n2);
   U4 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(2));
   U6 : XOR2_X1 port map( A => Ci, B => B(2), Z => n5);
   U7 : XOR2_X1 port map( A => A(2), B => n6, Z => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(1));
   U9 : XNOR2_X1 port map( A => n9, B => A(1), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n7);
   U11 : MUX2_X1 port map( A => n10, B => n11, S => Ci, Z => S(0));
   U12 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n12, ZN => n11);
   U13 : XOR2_X1 port map( A => B(0), B => A(0), Z => n10);
   U14 : OAI21_X1 port map( B1 => n13, B2 => n3, A => n14, ZN => Co);
   U15 : OAI21_X1 port map( B1 => n15, B2 => A(3), A => B(3), ZN => n14);
   U16 : INV_X1 port map( A => n3, ZN => n15);
   U17 : OAI21_X1 port map( B1 => A(2), B2 => n6, A => n16, ZN => n3);
   U18 : INV_X1 port map( A => n17, ZN => n16);
   U19 : AOI21_X1 port map( B1 => n6, B2 => A(2), A => B(2), ZN => n17);
   U20 : OAI21_X1 port map( B1 => n12, B2 => n18, A => n19, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n9, B2 => A(1), A => B(1), ZN => n19);
   U22 : INV_X1 port map( A => n12, ZN => n9);
   U23 : INV_X1 port map( A => A(1), ZN => n18);
   U24 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n12);
   U25 : INV_X1 port map( A => A(3), ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_0 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_0;

architecture SYN_BEHAVIORAL of PG_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_0 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_0;

architecture SYN_BEHAVIORAL of G_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_0 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_0;

architecture SYN_BEHAVIORAL of pg_generator_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_0;

architecture SYN_STRUCTURAL of CarrySelect_0 is

   component MUX21_GENERIC_bits4_0
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1370, n_1371 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1370);
   RCA2 : RCA_NBITS4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1371);
   MUX21_GEN : MUX21_GENERIC_bits4_0 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4 is

   port( A, B : in std_logic_vector (32 downto 1);  C0 : in std_logic;  COUT : 
         out std_logic_vector (8 downto 0));

end CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4;

architecture SYN_STRUCTURAL of CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_1
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_2
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_3
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_4
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_1
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_2
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_5
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_6
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_3
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_4
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_5
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_7
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_6
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_7
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_8
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_9
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_10
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_11
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_12
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_8
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_13
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_14
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_15
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_16
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_17
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_18
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_19
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_20
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_21
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_22
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_23
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_24
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_25
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_26
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_0
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_0
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component pg_generator_1
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_2
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_3
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_4
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_5
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_6
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_7
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_8
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_9
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_10
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_11
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_12
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_13
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_14
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_15
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_16
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_17
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_18
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_19
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_20
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_21
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_22
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_23
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_24
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_25
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_26
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_27
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_28
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_29
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_30
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_31
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_0
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   signal COUT_8_port, COUT_7_port, COUT_6_port, COUT_5_port, COUT_4_port, 
      COUT_3_port, COUT_2_port, COUT_1_port, gi_1_port, pi_1_port, 
      gSignal_16_16_port, gSignal_16_15_port, gSignal_16_13_port, 
      gSignal_16_9_port, gSignal_15_15_port, gSignal_14_14_port, 
      gSignal_14_13_port, gSignal_13_13_port, gSignal_12_12_port, 
      gSignal_12_11_port, gSignal_12_9_port, gSignal_11_11_port, 
      gSignal_10_10_port, gSignal_10_9_port, gSignal_9_9_port, gSignal_8_8_port
      , gSignal_8_7_port, gSignal_8_5_port, gSignal_7_7_port, gSignal_6_6_port,
      gSignal_6_5_port, gSignal_5_5_port, gSignal_4_4_port, gSignal_4_3_port, 
      gSignal_3_3_port, gSignal_2_2_port, gSignal_2_1_port, pSignal_16_16_port,
      pSignal_16_15_port, pSignal_16_13_port, pSignal_16_9_port, 
      pSignal_15_15_port, pSignal_14_14_port, pSignal_14_13_port, 
      pSignal_13_13_port, pSignal_12_12_port, pSignal_12_11_port, 
      pSignal_12_9_port, pSignal_11_11_port, pSignal_10_10_port, 
      pSignal_10_9_port, pSignal_9_9_port, pSignal_8_8_port, pSignal_8_7_port, 
      pSignal_8_5_port, pSignal_7_7_port, pSignal_6_6_port, pSignal_6_5_port, 
      pSignal_5_5_port, pSignal_4_4_port, pSignal_4_3_port, pSignal_3_3_port, 
      pSignal_2_2_port, pSignal_32_32_port, pSignal_32_31_port, 
      pSignal_32_29_port, pSignal_32_25_port, pSignal_32_17_port, 
      pSignal_31_31_port, pSignal_30_30_port, pSignal_30_29_port, 
      pSignal_29_29_port, pSignal_28_28_port, pSignal_28_27_port, 
      pSignal_28_25_port, pSignal_28_17_port, pSignal_27_27_port, 
      pSignal_26_26_port, pSignal_26_25_port, pSignal_25_25_port, 
      pSignal_24_24_port, pSignal_24_23_port, pSignal_24_21_port, 
      pSignal_24_17_port, pSignal_23_23_port, pSignal_22_22_port, 
      pSignal_22_21_port, pSignal_21_21_port, pSignal_20_20_port, 
      pSignal_20_19_port, pSignal_20_17_port, pSignal_19_19_port, 
      pSignal_18_18_port, pSignal_18_17_port, pSignal_17_17_port, 
      gSignal_32_32_port, gSignal_32_31_port, gSignal_32_29_port, 
      gSignal_32_25_port, gSignal_32_17_port, gSignal_31_31_port, 
      gSignal_30_30_port, gSignal_30_29_port, gSignal_29_29_port, 
      gSignal_28_28_port, gSignal_28_27_port, gSignal_28_25_port, 
      gSignal_28_17_port, gSignal_27_27_port, gSignal_26_26_port, 
      gSignal_26_25_port, gSignal_25_25_port, gSignal_24_24_port, 
      gSignal_24_23_port, gSignal_24_21_port, gSignal_24_17_port, 
      gSignal_23_23_port, gSignal_22_22_port, gSignal_22_21_port, 
      gSignal_21_21_port, gSignal_20_20_port, gSignal_20_19_port, 
      gSignal_20_17_port, gSignal_19_19_port, gSignal_18_18_port, 
      gSignal_18_17_port, gSignal_17_17_port, n1, n2 : std_logic;

begin
   COUT <= ( COUT_8_port, COUT_7_port, COUT_6_port, COUT_5_port, COUT_4_port, 
      COUT_3_port, COUT_2_port, COUT_1_port, C0 );
   
   pg_inst_1 : pg_generator_0 port map( A => A(1), B => B(1), P => pi_1_port, G
                           => gi_1_port);
   pg_inst_2 : pg_generator_31 port map( A => A(2), B => B(2), P => 
                           pSignal_2_2_port, G => gSignal_2_2_port);
   pg_inst_3 : pg_generator_30 port map( A => A(3), B => B(3), P => 
                           pSignal_3_3_port, G => gSignal_3_3_port);
   pg_inst_4 : pg_generator_29 port map( A => A(4), B => B(4), P => 
                           pSignal_4_4_port, G => gSignal_4_4_port);
   pg_inst_5 : pg_generator_28 port map( A => A(5), B => B(5), P => 
                           pSignal_5_5_port, G => gSignal_5_5_port);
   pg_inst_6 : pg_generator_27 port map( A => A(6), B => B(6), P => 
                           pSignal_6_6_port, G => gSignal_6_6_port);
   pg_inst_7 : pg_generator_26 port map( A => A(7), B => B(7), P => 
                           pSignal_7_7_port, G => gSignal_7_7_port);
   pg_inst_8 : pg_generator_25 port map( A => A(8), B => B(8), P => 
                           pSignal_8_8_port, G => gSignal_8_8_port);
   pg_inst_9 : pg_generator_24 port map( A => A(9), B => B(9), P => 
                           pSignal_9_9_port, G => gSignal_9_9_port);
   pg_inst_10 : pg_generator_23 port map( A => A(10), B => B(10), P => 
                           pSignal_10_10_port, G => gSignal_10_10_port);
   pg_inst_11 : pg_generator_22 port map( A => A(11), B => B(11), P => 
                           pSignal_11_11_port, G => gSignal_11_11_port);
   pg_inst_12 : pg_generator_21 port map( A => A(12), B => B(12), P => 
                           pSignal_12_12_port, G => gSignal_12_12_port);
   pg_inst_13 : pg_generator_20 port map( A => A(13), B => B(13), P => 
                           pSignal_13_13_port, G => gSignal_13_13_port);
   pg_inst_14 : pg_generator_19 port map( A => A(14), B => B(14), P => 
                           pSignal_14_14_port, G => gSignal_14_14_port);
   pg_inst_15 : pg_generator_18 port map( A => A(15), B => B(15), P => 
                           pSignal_15_15_port, G => gSignal_15_15_port);
   pg_inst_16 : pg_generator_17 port map( A => A(16), B => B(16), P => 
                           pSignal_16_16_port, G => gSignal_16_16_port);
   pg_inst_17 : pg_generator_16 port map( A => A(17), B => B(17), P => 
                           pSignal_17_17_port, G => gSignal_17_17_port);
   pg_inst_18 : pg_generator_15 port map( A => A(18), B => B(18), P => 
                           pSignal_18_18_port, G => gSignal_18_18_port);
   pg_inst_19 : pg_generator_14 port map( A => A(19), B => B(19), P => 
                           pSignal_19_19_port, G => gSignal_19_19_port);
   pg_inst_20 : pg_generator_13 port map( A => A(20), B => B(20), P => 
                           pSignal_20_20_port, G => gSignal_20_20_port);
   pg_inst_21 : pg_generator_12 port map( A => A(21), B => B(21), P => 
                           pSignal_21_21_port, G => gSignal_21_21_port);
   pg_inst_22 : pg_generator_11 port map( A => A(22), B => B(22), P => 
                           pSignal_22_22_port, G => gSignal_22_22_port);
   pg_inst_23 : pg_generator_10 port map( A => A(23), B => B(23), P => 
                           pSignal_23_23_port, G => gSignal_23_23_port);
   pg_inst_24 : pg_generator_9 port map( A => A(24), B => B(24), P => 
                           pSignal_24_24_port, G => gSignal_24_24_port);
   pg_inst_25 : pg_generator_8 port map( A => A(25), B => B(25), P => 
                           pSignal_25_25_port, G => gSignal_25_25_port);
   pg_inst_26 : pg_generator_7 port map( A => A(26), B => B(26), P => 
                           pSignal_26_26_port, G => gSignal_26_26_port);
   pg_inst_27 : pg_generator_6 port map( A => A(27), B => B(27), P => 
                           pSignal_27_27_port, G => gSignal_27_27_port);
   pg_inst_28 : pg_generator_5 port map( A => A(28), B => B(28), P => 
                           pSignal_28_28_port, G => gSignal_28_28_port);
   pg_inst_29 : pg_generator_4 port map( A => A(29), B => B(29), P => 
                           pSignal_29_29_port, G => gSignal_29_29_port);
   pg_inst_30 : pg_generator_3 port map( A => A(30), B => B(30), P => 
                           pSignal_30_30_port, G => gSignal_30_30_port);
   pg_inst_31 : pg_generator_2 port map( A => A(31), B => B(31), P => 
                           pSignal_31_31_port, G => gSignal_31_31_port);
   pg_inst_32 : pg_generator_1 port map( A => A(32), B => B(32), P => 
                           pSignal_32_32_port, G => gSignal_32_32_port);
   G1_1_2 : G_0 port map( p_ik => pSignal_2_2_port, g_ik => gSignal_2_2_port, 
                           g_k1j => n2, G_ij => gSignal_2_1_port);
   PG_inst1_1_4 : PG_0 port map( p_ik => pSignal_4_4_port, g_ik => 
                           gSignal_4_4_port, p_k1j => pSignal_3_3_port, g_k1j 
                           => gSignal_3_3_port, P_ij => pSignal_4_3_port, G_ij 
                           => gSignal_4_3_port);
   PG_inst1_1_6 : PG_26 port map( p_ik => pSignal_6_6_port, g_ik => 
                           gSignal_6_6_port, p_k1j => pSignal_5_5_port, g_k1j 
                           => gSignal_5_5_port, P_ij => pSignal_6_5_port, G_ij 
                           => gSignal_6_5_port);
   PG_inst1_1_8 : PG_25 port map( p_ik => pSignal_8_8_port, g_ik => 
                           gSignal_8_8_port, p_k1j => pSignal_7_7_port, g_k1j 
                           => gSignal_7_7_port, P_ij => pSignal_8_7_port, G_ij 
                           => gSignal_8_7_port);
   PG_inst1_1_10 : PG_24 port map( p_ik => pSignal_10_10_port, g_ik => 
                           gSignal_10_10_port, p_k1j => pSignal_9_9_port, g_k1j
                           => gSignal_9_9_port, P_ij => pSignal_10_9_port, G_ij
                           => gSignal_10_9_port);
   PG_inst1_1_12 : PG_23 port map( p_ik => pSignal_12_12_port, g_ik => 
                           gSignal_12_12_port, p_k1j => pSignal_11_11_port, 
                           g_k1j => gSignal_11_11_port, P_ij => 
                           pSignal_12_11_port, G_ij => gSignal_12_11_port);
   PG_inst1_1_14 : PG_22 port map( p_ik => pSignal_14_14_port, g_ik => 
                           gSignal_14_14_port, p_k1j => pSignal_13_13_port, 
                           g_k1j => gSignal_13_13_port, P_ij => 
                           pSignal_14_13_port, G_ij => gSignal_14_13_port);
   PG_inst1_1_16 : PG_21 port map( p_ik => pSignal_16_16_port, g_ik => 
                           gSignal_16_16_port, p_k1j => pSignal_15_15_port, 
                           g_k1j => gSignal_15_15_port, P_ij => 
                           pSignal_16_15_port, G_ij => gSignal_16_15_port);
   PG_inst1_1_18 : PG_20 port map( p_ik => pSignal_18_18_port, g_ik => 
                           gSignal_18_18_port, p_k1j => pSignal_17_17_port, 
                           g_k1j => gSignal_17_17_port, P_ij => 
                           pSignal_18_17_port, G_ij => gSignal_18_17_port);
   PG_inst1_1_20 : PG_19 port map( p_ik => pSignal_20_20_port, g_ik => 
                           gSignal_20_20_port, p_k1j => pSignal_19_19_port, 
                           g_k1j => gSignal_19_19_port, P_ij => 
                           pSignal_20_19_port, G_ij => gSignal_20_19_port);
   PG_inst1_1_22 : PG_18 port map( p_ik => pSignal_22_22_port, g_ik => 
                           gSignal_22_22_port, p_k1j => pSignal_21_21_port, 
                           g_k1j => gSignal_21_21_port, P_ij => 
                           pSignal_22_21_port, G_ij => gSignal_22_21_port);
   PG_inst1_1_24 : PG_17 port map( p_ik => pSignal_24_24_port, g_ik => 
                           gSignal_24_24_port, p_k1j => pSignal_23_23_port, 
                           g_k1j => gSignal_23_23_port, P_ij => 
                           pSignal_24_23_port, G_ij => gSignal_24_23_port);
   PG_inst1_1_26 : PG_16 port map( p_ik => pSignal_26_26_port, g_ik => 
                           gSignal_26_26_port, p_k1j => pSignal_25_25_port, 
                           g_k1j => gSignal_25_25_port, P_ij => 
                           pSignal_26_25_port, G_ij => gSignal_26_25_port);
   PG_inst1_1_28 : PG_15 port map( p_ik => pSignal_28_28_port, g_ik => 
                           gSignal_28_28_port, p_k1j => pSignal_27_27_port, 
                           g_k1j => gSignal_27_27_port, P_ij => 
                           pSignal_28_27_port, G_ij => gSignal_28_27_port);
   PG_inst1_1_30 : PG_14 port map( p_ik => pSignal_30_30_port, g_ik => 
                           gSignal_30_30_port, p_k1j => pSignal_29_29_port, 
                           g_k1j => gSignal_29_29_port, P_ij => 
                           pSignal_30_29_port, G_ij => gSignal_30_29_port);
   PG_inst1_1_32 : PG_13 port map( p_ik => pSignal_32_32_port, g_ik => 
                           gSignal_32_32_port, p_k1j => pSignal_31_31_port, 
                           g_k1j => gSignal_31_31_port, P_ij => 
                           pSignal_32_31_port, G_ij => gSignal_32_31_port);
   G1_2_4 : G_8 port map( p_ik => pSignal_4_3_port, g_ik => gSignal_4_3_port, 
                           g_k1j => gSignal_2_1_port, G_ij => COUT_1_port);
   PG_inst1_2_8 : PG_12 port map( p_ik => pSignal_8_7_port, g_ik => 
                           gSignal_8_7_port, p_k1j => pSignal_6_5_port, g_k1j 
                           => gSignal_6_5_port, P_ij => pSignal_8_5_port, G_ij 
                           => gSignal_8_5_port);
   PG_inst1_2_12 : PG_11 port map( p_ik => pSignal_12_11_port, g_ik => 
                           gSignal_12_11_port, p_k1j => pSignal_10_9_port, 
                           g_k1j => gSignal_10_9_port, P_ij => 
                           pSignal_12_9_port, G_ij => gSignal_12_9_port);
   PG_inst1_2_16 : PG_10 port map( p_ik => pSignal_16_15_port, g_ik => 
                           gSignal_16_15_port, p_k1j => pSignal_14_13_port, 
                           g_k1j => gSignal_14_13_port, P_ij => 
                           pSignal_16_13_port, G_ij => gSignal_16_13_port);
   PG_inst1_2_20 : PG_9 port map( p_ik => pSignal_20_19_port, g_ik => 
                           gSignal_20_19_port, p_k1j => pSignal_18_17_port, 
                           g_k1j => gSignal_18_17_port, P_ij => 
                           pSignal_20_17_port, G_ij => gSignal_20_17_port);
   PG_inst1_2_24 : PG_8 port map( p_ik => pSignal_24_23_port, g_ik => 
                           gSignal_24_23_port, p_k1j => pSignal_22_21_port, 
                           g_k1j => gSignal_22_21_port, P_ij => 
                           pSignal_24_21_port, G_ij => gSignal_24_21_port);
   PG_inst1_2_28 : PG_7 port map( p_ik => pSignal_28_27_port, g_ik => 
                           gSignal_28_27_port, p_k1j => pSignal_26_25_port, 
                           g_k1j => gSignal_26_25_port, P_ij => 
                           pSignal_28_25_port, G_ij => gSignal_28_25_port);
   PG_inst1_2_32 : PG_6 port map( p_ik => pSignal_32_31_port, g_ik => 
                           gSignal_32_31_port, p_k1j => pSignal_30_29_port, 
                           g_k1j => gSignal_30_29_port, P_ij => 
                           pSignal_32_29_port, G_ij => gSignal_32_29_port);
   G_INST2_0_4_8 : G_7 port map( p_ik => pSignal_8_5_port, g_ik => 
                           gSignal_8_5_port, g_k1j => COUT_1_port, G_ij => 
                           COUT_2_port);
   PG_INST2_0_12_16 : PG_5 port map( p_ik => pSignal_16_13_port, g_ik => 
                           gSignal_16_13_port, p_k1j => pSignal_12_9_port, 
                           g_k1j => gSignal_12_9_port, P_ij => 
                           pSignal_16_9_port, G_ij => gSignal_16_9_port);
   PG_INST2_0_20_24 : PG_4 port map( p_ik => pSignal_24_21_port, g_ik => 
                           gSignal_24_21_port, p_k1j => pSignal_20_17_port, 
                           g_k1j => gSignal_20_17_port, P_ij => 
                           pSignal_24_17_port, G_ij => gSignal_24_17_port);
   PG_INST2_0_28_32 : PG_3 port map( p_ik => pSignal_32_29_port, g_ik => 
                           gSignal_32_29_port, p_k1j => pSignal_28_25_port, 
                           g_k1j => gSignal_28_25_port, P_ij => 
                           pSignal_32_25_port, G_ij => gSignal_32_25_port);
   G_INST2_1_8_12 : G_6 port map( p_ik => pSignal_12_9_port, g_ik => 
                           gSignal_12_9_port, g_k1j => COUT_2_port, G_ij => 
                           COUT_3_port);
   G_INST2_1_8_16 : G_5 port map( p_ik => pSignal_16_9_port, g_ik => 
                           gSignal_16_9_port, g_k1j => COUT_2_port, G_ij => 
                           COUT_4_port);
   PG_INST2_1_24_28 : PG_2 port map( p_ik => pSignal_28_25_port, g_ik => 
                           gSignal_28_25_port, p_k1j => pSignal_24_17_port, 
                           g_k1j => gSignal_24_17_port, P_ij => 
                           pSignal_28_17_port, G_ij => gSignal_28_17_port);
   PG_INST2_1_24_32 : PG_1 port map( p_ik => pSignal_32_25_port, g_ik => 
                           gSignal_32_25_port, p_k1j => pSignal_24_17_port, 
                           g_k1j => gSignal_24_17_port, P_ij => 
                           pSignal_32_17_port, G_ij => gSignal_32_17_port);
   G_INST2_2_16_20 : G_4 port map( p_ik => pSignal_20_17_port, g_ik => 
                           gSignal_20_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_5_port);
   G_INST2_2_16_24 : G_3 port map( p_ik => pSignal_24_17_port, g_ik => 
                           gSignal_24_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_6_port);
   G_INST2_2_16_28 : G_2 port map( p_ik => pSignal_28_17_port, g_ik => 
                           gSignal_28_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_7_port);
   G_INST2_2_16_32 : G_1 port map( p_ik => pSignal_32_17_port, g_ik => 
                           gSignal_32_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_8_port);
   U1 : INV_X1 port map( A => n1, ZN => n2);
   U2 : AOI21_X1 port map( B1 => pi_1_port, B2 => C0, A => gi_1_port, ZN => n1)
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (8
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8;

architecture SYN_STRUCTURAL of 
   SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8 is

   component CarrySelect_1
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_2
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_3
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_4
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_5
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_6
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_7
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_0
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   carrySel_0 : CarrySelect_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Cin => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   carrySel_1 : CarrySelect_7 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Cin => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   carrySel_2 : CarrySelect_6 port map( A(3) => A(11), A(2) => A(10), A(1) => 
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Cin => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   carrySel_3 : CarrySelect_5 port map( A(3) => A(15), A(2) => A(14), A(1) => 
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Cin => Ci(3), S(3) => 
                           S(15), S(2) => S(14), S(1) => S(13), S(0) => S(12));
   carrySel_4 : CarrySelect_4 port map( A(3) => A(19), A(2) => A(18), A(1) => 
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Cin => Ci(4), S(3) => 
                           S(19), S(2) => S(18), S(1) => S(17), S(0) => S(16));
   carrySel_5 : CarrySelect_3 port map( A(3) => A(23), A(2) => A(22), A(1) => 
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Cin => Ci(5), S(3) => 
                           S(23), S(2) => S(22), S(1) => S(21), S(0) => S(20));
   carrySel_6 : CarrySelect_2 port map( A(3) => A(27), A(2) => A(26), A(1) => 
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Cin => Ci(6), S(3) => 
                           S(27), S(2) => S(26), S(1) => S(25), S(0) => S(24));
   carrySel_7 : CarrySelect_1 port map( A(3) => A(31), A(2) => A(30), A(1) => 
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Cin => Ci(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_logic_nbits32 is

   port( Cin : in std_logic;  B0 : in std_logic_vector (31 downto 0);  B : out 
         std_logic_vector (31 downto 0));

end xor_logic_nbits32;

architecture SYN_BEHAVIORAL of xor_logic_nbits32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => Cin, B => B0(9), Z => B(9));
   U2 : XOR2_X1 port map( A => Cin, B => B0(8), Z => B(8));
   U3 : XOR2_X1 port map( A => Cin, B => B0(7), Z => B(7));
   U4 : XOR2_X1 port map( A => Cin, B => B0(6), Z => B(6));
   U5 : XOR2_X1 port map( A => Cin, B => B0(5), Z => B(5));
   U6 : XOR2_X1 port map( A => Cin, B => B0(4), Z => B(4));
   U7 : XOR2_X1 port map( A => Cin, B => B0(3), Z => B(3));
   U8 : XOR2_X1 port map( A => Cin, B => B0(31), Z => B(31));
   U9 : XOR2_X1 port map( A => Cin, B => B0(30), Z => B(30));
   U10 : XOR2_X1 port map( A => Cin, B => B0(2), Z => B(2));
   U11 : XOR2_X1 port map( A => Cin, B => B0(29), Z => B(29));
   U12 : XOR2_X1 port map( A => Cin, B => B0(28), Z => B(28));
   U13 : XOR2_X1 port map( A => Cin, B => B0(27), Z => B(27));
   U14 : XOR2_X1 port map( A => Cin, B => B0(26), Z => B(26));
   U15 : XOR2_X1 port map( A => Cin, B => B0(25), Z => B(25));
   U16 : XOR2_X1 port map( A => Cin, B => B0(24), Z => B(24));
   U17 : XOR2_X1 port map( A => Cin, B => B0(23), Z => B(23));
   U18 : XOR2_X1 port map( A => Cin, B => B0(22), Z => B(22));
   U19 : XOR2_X1 port map( A => Cin, B => B0(21), Z => B(21));
   U20 : XOR2_X1 port map( A => Cin, B => B0(20), Z => B(20));
   U21 : XOR2_X1 port map( A => Cin, B => B0(1), Z => B(1));
   U22 : XOR2_X1 port map( A => Cin, B => B0(19), Z => B(19));
   U23 : XOR2_X1 port map( A => Cin, B => B0(18), Z => B(18));
   U24 : XOR2_X1 port map( A => Cin, B => B0(17), Z => B(17));
   U25 : XOR2_X1 port map( A => Cin, B => B0(16), Z => B(16));
   U26 : XOR2_X1 port map( A => Cin, B => B0(15), Z => B(15));
   U27 : XOR2_X1 port map( A => Cin, B => B0(14), Z => B(14));
   U28 : XOR2_X1 port map( A => Cin, B => B0(13), Z => B(13));
   U29 : XOR2_X1 port map( A => Cin, B => B0(12), Z => B(12));
   U30 : XOR2_X1 port map( A => Cin, B => B0(11), Z => B(11));
   U31 : XOR2_X1 port map( A => Cin, B => B0(10), Z => B(10));
   U32 : XOR2_X1 port map( A => Cin, B => B0(0), Z => B(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity logic_and_shift_N32 is

   port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
         downto 0));

end logic_and_shift_N32;

architecture SYN_BEHAVIOR of logic_and_shift_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component logic_and_shift_N32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component logic_and_shift_N32_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,
      N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57
      , N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, 
      N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86
      , N87, N88, N89, N90, N91, N92, N190, N191, N192, N193, N194, N195, N196,
      N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, 
      N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, 
      N221, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29_port
      , n30_port, n31_port, n32_port, n33_port, n34_port, n35_port, n36_port, 
      n37_port, n38_port, n39_port, n40_port, n41_port, n42_port, n43_port, 
      n44_port, n45_port, n46_port, n47_port, n48_port, n49_port, n50_port, 
      n51_port, n52_port, n53_port, n54_port, n55_port, n56_port, n57_port, 
      n58_port, n59_port, n60_port, n61_port, n62_port, n63_port, n64_port, 
      n65_port, n66_port, n67_port, n68_port, n69_port, n70_port, n71_port, 
      n72_port, n73_port, n74_port, n75_port, n76_port, n77_port, n78_port, 
      n79_port, n80_port, n81_port, n82_port, n83_port, n84_port, n85_port, 
      n86_port, n87_port, n88_port, n89_port, n90_port, n91_port, n92_port, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190_port, n191_port, n192_port, n193_port, n194_port, n195_port, 
      n196_port, n197_port, n198_port, n199_port, n200_port, n201_port, 
      n202_port, n203_port, n204_port, n205_port, n206_port : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   OUTALU_reg_31_inst : DLH_X1 port map( G => n4, D => N221, Q => OUTALU(31));
   OUTALU_reg_30_inst : DLH_X1 port map( G => n4, D => N220, Q => OUTALU(30));
   OUTALU_reg_29_inst : DLH_X1 port map( G => n4, D => N219, Q => OUTALU(29));
   OUTALU_reg_28_inst : DLH_X1 port map( G => n4, D => N218, Q => OUTALU(28));
   OUTALU_reg_27_inst : DLH_X1 port map( G => n4, D => N217, Q => OUTALU(27));
   OUTALU_reg_26_inst : DLH_X1 port map( G => n4, D => N216, Q => OUTALU(26));
   OUTALU_reg_25_inst : DLH_X1 port map( G => n4, D => N215, Q => OUTALU(25));
   OUTALU_reg_24_inst : DLH_X1 port map( G => n4, D => N214, Q => OUTALU(24));
   OUTALU_reg_23_inst : DLH_X1 port map( G => n4, D => N213, Q => OUTALU(23));
   OUTALU_reg_22_inst : DLH_X1 port map( G => n4, D => N212, Q => OUTALU(22));
   OUTALU_reg_21_inst : DLH_X1 port map( G => n4, D => N211, Q => OUTALU(21));
   OUTALU_reg_20_inst : DLH_X1 port map( G => n4, D => N210, Q => OUTALU(20));
   OUTALU_reg_19_inst : DLH_X1 port map( G => n4, D => N209, Q => OUTALU(19));
   OUTALU_reg_18_inst : DLH_X1 port map( G => n4, D => N208, Q => OUTALU(18));
   OUTALU_reg_17_inst : DLH_X1 port map( G => n4, D => N207, Q => OUTALU(17));
   OUTALU_reg_16_inst : DLH_X1 port map( G => n4, D => N206, Q => OUTALU(16));
   OUTALU_reg_15_inst : DLH_X1 port map( G => n4, D => N205, Q => OUTALU(15));
   OUTALU_reg_14_inst : DLH_X1 port map( G => n4, D => N204, Q => OUTALU(14));
   OUTALU_reg_13_inst : DLH_X1 port map( G => n4, D => N203, Q => OUTALU(13));
   OUTALU_reg_12_inst : DLH_X1 port map( G => n4, D => N202, Q => OUTALU(12));
   OUTALU_reg_11_inst : DLH_X1 port map( G => n4, D => N201, Q => OUTALU(11));
   OUTALU_reg_10_inst : DLH_X1 port map( G => n4, D => N200, Q => OUTALU(10));
   OUTALU_reg_9_inst : DLH_X1 port map( G => n4, D => N199, Q => OUTALU(9));
   OUTALU_reg_8_inst : DLH_X1 port map( G => n4, D => N198, Q => OUTALU(8));
   OUTALU_reg_7_inst : DLH_X1 port map( G => n4, D => N197, Q => OUTALU(7));
   OUTALU_reg_6_inst : DLH_X1 port map( G => n4, D => N196, Q => OUTALU(6));
   OUTALU_reg_5_inst : DLH_X1 port map( G => n4, D => N195, Q => OUTALU(5));
   OUTALU_reg_4_inst : DLH_X1 port map( G => n4, D => N194, Q => OUTALU(4));
   OUTALU_reg_3_inst : DLH_X1 port map( G => n4, D => N193, Q => OUTALU(3));
   OUTALU_reg_2_inst : DLH_X1 port map( G => n4, D => N192, Q => OUTALU(2));
   OUTALU_reg_1_inst : DLH_X1 port map( G => n4, D => N191, Q => OUTALU(1));
   OUTALU_reg_0_inst : DLH_X1 port map( G => n4, D => N190, Q => OUTALU(0));
   srl_39 : logic_and_shift_N32_DW_rash_0 port map( A(31) => DATA1(31), A(30) 
                           => DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28)
                           , A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), DATA_TC => n1,
                           SH(30) => DATA2(30), SH(29) => DATA2(29), SH(28) => 
                           DATA2(28), SH(27) => DATA2(27), SH(26) => DATA2(26),
                           SH(25) => DATA2(25), SH(24) => DATA2(24), SH(23) => 
                           DATA2(23), SH(22) => DATA2(22), SH(21) => DATA2(21),
                           SH(20) => DATA2(20), SH(19) => DATA2(19), SH(18) => 
                           DATA2(18), SH(17) => DATA2(17), SH(16) => DATA2(16),
                           SH(15) => DATA2(15), SH(14) => DATA2(14), SH(13) => 
                           DATA2(13), SH(12) => DATA2(12), SH(11) => DATA2(11),
                           SH(10) => DATA2(10), SH(9) => DATA2(9), SH(8) => 
                           DATA2(8), SH(7) => DATA2(7), SH(6) => DATA2(6), 
                           SH(5) => DATA2(5), SH(4) => DATA2(4), SH(3) => 
                           DATA2(3), SH(2) => DATA2(2), SH(1) => DATA2(1), 
                           SH(0) => DATA2(0), SH_TC => n1, B(31) => N92, B(30) 
                           => N91, B(29) => N90, B(28) => N89, B(27) => N88, 
                           B(26) => N87, B(25) => N86, B(24) => N85, B(23) => 
                           N84, B(22) => N83, B(21) => N82, B(20) => N81, B(19)
                           => N80, B(18) => N79, B(17) => N78, B(16) => N77, 
                           B(15) => N76, B(14) => N75, B(13) => N74, B(12) => 
                           N73, B(11) => N72, B(10) => N71, B(9) => N70, B(8) 
                           => N69, B(7) => N68, B(6) => N67, B(5) => N66, B(4) 
                           => N65, B(3) => N64, B(2) => N63, B(1) => N62, B(0) 
                           => N61);
   sll_37 : logic_and_shift_N32_DW01_ash_0 port map( A(31) => DATA1(31), A(30) 
                           => DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28)
                           , A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), DATA_TC => n2,
                           SH(30) => DATA2(30), SH(29) => DATA2(29), SH(28) => 
                           DATA2(28), SH(27) => DATA2(27), SH(26) => DATA2(26),
                           SH(25) => DATA2(25), SH(24) => DATA2(24), SH(23) => 
                           DATA2(23), SH(22) => DATA2(22), SH(21) => DATA2(21),
                           SH(20) => DATA2(20), SH(19) => DATA2(19), SH(18) => 
                           DATA2(18), SH(17) => DATA2(17), SH(16) => DATA2(16),
                           SH(15) => DATA2(15), SH(14) => DATA2(14), SH(13) => 
                           DATA2(13), SH(12) => DATA2(12), SH(11) => DATA2(11),
                           SH(10) => DATA2(10), SH(9) => DATA2(9), SH(8) => 
                           DATA2(8), SH(7) => DATA2(7), SH(6) => DATA2(6), 
                           SH(5) => DATA2(5), SH(4) => DATA2(4), SH(3) => 
                           DATA2(3), SH(2) => DATA2(2), SH(1) => DATA2(1), 
                           SH(0) => DATA2(0), SH_TC => n2, B(31) => N60, B(30) 
                           => N59, B(29) => N58, B(28) => N57, B(27) => N56, 
                           B(26) => N55, B(25) => N54, B(24) => N53, B(23) => 
                           N52, B(22) => N51, B(21) => N50, B(20) => N49, B(19)
                           => N48, B(18) => N47, B(17) => N46, B(16) => N45, 
                           B(15) => N44, B(14) => N43, B(13) => N42, B(12) => 
                           N41, B(11) => N40, B(10) => N39, B(9) => N38, B(8) 
                           => N37, B(7) => N36, B(6) => N35, B(5) => N34, B(4) 
                           => N33, B(3) => N32, B(2) => N31, B(1) => N30, B(0) 
                           => N29);
   U3 : OR2_X1 port map( A1 => FUNC(0), A2 => n7, ZN => n3);
   U4 : INV_X1 port map( A => n3, ZN => n4);
   U7 : AND3_X4 port map( A1 => FUNC(2), A2 => n203_port, A3 => FUNC(1), ZN => 
                           n8);
   U8 : AND2_X4 port map( A1 => n9, A2 => FUNC(3), ZN => n16);
   U9 : NOR2_X4 port map( A1 => n206_port, A2 => FUNC(2), ZN => n9);
   U10 : OR3_X1 port map( A1 => FUNC(2), A2 => FUNC(1), A3 => n203_port, ZN => 
                           n10);
   U11 : INV_X2 port map( A => n10, ZN => n5);
   U12 : OR3_X1 port map( A1 => FUNC(2), A2 => FUNC(1), A3 => FUNC(3), ZN => 
                           n11);
   U13 : INV_X2 port map( A => n11, ZN => n6);
   U14 : NOR4_X1 port map( A1 => n8, A2 => n9, A3 => n5, A4 => n6, ZN => n7);
   U15 : OAI211_X1 port map( C1 => n12, C2 => n13, A => n14, B => n15, ZN => 
                           N221);
   U16 : AOI22_X1 port map( A1 => N60, A2 => n6, B1 => N92, B2 => n5, ZN => n15
                           );
   U17 : OAI21_X1 port map( B1 => n16, B2 => n17, A => DATA2(31), ZN => n14);
   U18 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(31), Z => n17);
   U19 : INV_X1 port map( A => DATA1(31), ZN => n13);
   U20 : AOI21_X1 port map( B1 => n8, B2 => n18, A => n16, ZN => n12);
   U21 : INV_X1 port map( A => DATA2(31), ZN => n18);
   U22 : OAI211_X1 port map( C1 => n19, C2 => n20, A => n21, B => n22, ZN => 
                           N220);
   U23 : AOI22_X1 port map( A1 => N59, A2 => n6, B1 => N91, B2 => n5, ZN => n22
                           );
   U24 : OAI21_X1 port map( B1 => n16, B2 => n23, A => DATA2(30), ZN => n21);
   U25 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(30), Z => n23);
   U26 : INV_X1 port map( A => DATA1(30), ZN => n20);
   U27 : AOI21_X1 port map( B1 => n8, B2 => n24, A => n16, ZN => n19);
   U28 : INV_X1 port map( A => DATA2(30), ZN => n24);
   U29 : OAI211_X1 port map( C1 => n25, C2 => n26, A => n27, B => n28, ZN => 
                           N219);
   U30 : AOI22_X1 port map( A1 => N58, A2 => n6, B1 => N90, B2 => n5, ZN => n28
                           );
   U31 : OAI21_X1 port map( B1 => n16, B2 => n29_port, A => DATA2(29), ZN => 
                           n27);
   U32 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(29), Z => n29_port);
   U33 : INV_X1 port map( A => DATA1(29), ZN => n26);
   U34 : AOI21_X1 port map( B1 => n8, B2 => n30_port, A => n16, ZN => n25);
   U35 : INV_X1 port map( A => DATA2(29), ZN => n30_port);
   U36 : OAI211_X1 port map( C1 => n31_port, C2 => n32_port, A => n33_port, B 
                           => n34_port, ZN => N218);
   U37 : AOI22_X1 port map( A1 => N57, A2 => n6, B1 => N89, B2 => n5, ZN => 
                           n34_port);
   U38 : OAI21_X1 port map( B1 => n16, B2 => n35_port, A => DATA2(28), ZN => 
                           n33_port);
   U39 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(28), Z => n35_port);
   U40 : INV_X1 port map( A => DATA1(28), ZN => n32_port);
   U41 : AOI21_X1 port map( B1 => n8, B2 => n36_port, A => n16, ZN => n31_port)
                           ;
   U42 : INV_X1 port map( A => DATA2(28), ZN => n36_port);
   U43 : OAI211_X1 port map( C1 => n37_port, C2 => n38_port, A => n39_port, B 
                           => n40_port, ZN => N217);
   U44 : AOI22_X1 port map( A1 => N56, A2 => n6, B1 => N88, B2 => n5, ZN => 
                           n40_port);
   U45 : OAI21_X1 port map( B1 => n16, B2 => n41_port, A => DATA2(27), ZN => 
                           n39_port);
   U46 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(27), Z => n41_port);
   U47 : INV_X1 port map( A => DATA1(27), ZN => n38_port);
   U48 : AOI21_X1 port map( B1 => n8, B2 => n42_port, A => n16, ZN => n37_port)
                           ;
   U49 : INV_X1 port map( A => DATA2(27), ZN => n42_port);
   U50 : OAI211_X1 port map( C1 => n43_port, C2 => n44_port, A => n45_port, B 
                           => n46_port, ZN => N216);
   U51 : AOI22_X1 port map( A1 => N55, A2 => n6, B1 => N87, B2 => n5, ZN => 
                           n46_port);
   U52 : OAI21_X1 port map( B1 => n16, B2 => n47_port, A => DATA2(26), ZN => 
                           n45_port);
   U53 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(26), Z => n47_port);
   U54 : INV_X1 port map( A => DATA1(26), ZN => n44_port);
   U55 : AOI21_X1 port map( B1 => n8, B2 => n48_port, A => n16, ZN => n43_port)
                           ;
   U56 : INV_X1 port map( A => DATA2(26), ZN => n48_port);
   U57 : OAI211_X1 port map( C1 => n49_port, C2 => n50_port, A => n51_port, B 
                           => n52_port, ZN => N215);
   U58 : AOI22_X1 port map( A1 => N54, A2 => n6, B1 => N86, B2 => n5, ZN => 
                           n52_port);
   U59 : OAI21_X1 port map( B1 => n16, B2 => n53_port, A => DATA2(25), ZN => 
                           n51_port);
   U60 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(25), Z => n53_port);
   U61 : INV_X1 port map( A => DATA1(25), ZN => n50_port);
   U62 : AOI21_X1 port map( B1 => n8, B2 => n54_port, A => n16, ZN => n49_port)
                           ;
   U63 : INV_X1 port map( A => DATA2(25), ZN => n54_port);
   U64 : OAI211_X1 port map( C1 => n55_port, C2 => n56_port, A => n57_port, B 
                           => n58_port, ZN => N214);
   U65 : AOI22_X1 port map( A1 => N53, A2 => n6, B1 => N85, B2 => n5, ZN => 
                           n58_port);
   U66 : OAI21_X1 port map( B1 => n16, B2 => n59_port, A => DATA2(24), ZN => 
                           n57_port);
   U67 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(24), Z => n59_port);
   U68 : INV_X1 port map( A => DATA1(24), ZN => n56_port);
   U69 : AOI21_X1 port map( B1 => n8, B2 => n60_port, A => n16, ZN => n55_port)
                           ;
   U70 : INV_X1 port map( A => DATA2(24), ZN => n60_port);
   U71 : OAI211_X1 port map( C1 => n61_port, C2 => n62_port, A => n63_port, B 
                           => n64_port, ZN => N213);
   U72 : AOI22_X1 port map( A1 => N52, A2 => n6, B1 => N84, B2 => n5, ZN => 
                           n64_port);
   U73 : OAI21_X1 port map( B1 => n16, B2 => n65_port, A => DATA2(23), ZN => 
                           n63_port);
   U74 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(23), Z => n65_port);
   U75 : INV_X1 port map( A => DATA1(23), ZN => n62_port);
   U76 : AOI21_X1 port map( B1 => n8, B2 => n66_port, A => n16, ZN => n61_port)
                           ;
   U77 : INV_X1 port map( A => DATA2(23), ZN => n66_port);
   U78 : OAI211_X1 port map( C1 => n67_port, C2 => n68_port, A => n69_port, B 
                           => n70_port, ZN => N212);
   U79 : AOI22_X1 port map( A1 => N51, A2 => n6, B1 => N83, B2 => n5, ZN => 
                           n70_port);
   U80 : OAI21_X1 port map( B1 => n16, B2 => n71_port, A => DATA2(22), ZN => 
                           n69_port);
   U81 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(22), Z => n71_port);
   U82 : INV_X1 port map( A => DATA1(22), ZN => n68_port);
   U83 : AOI21_X1 port map( B1 => n8, B2 => n72_port, A => n16, ZN => n67_port)
                           ;
   U84 : INV_X1 port map( A => DATA2(22), ZN => n72_port);
   U85 : OAI211_X1 port map( C1 => n73_port, C2 => n74_port, A => n75_port, B 
                           => n76_port, ZN => N211);
   U86 : AOI22_X1 port map( A1 => N50, A2 => n6, B1 => N82, B2 => n5, ZN => 
                           n76_port);
   U87 : OAI21_X1 port map( B1 => n16, B2 => n77_port, A => DATA2(21), ZN => 
                           n75_port);
   U88 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(21), Z => n77_port);
   U89 : INV_X1 port map( A => DATA1(21), ZN => n74_port);
   U90 : AOI21_X1 port map( B1 => n8, B2 => n78_port, A => n16, ZN => n73_port)
                           ;
   U91 : INV_X1 port map( A => DATA2(21), ZN => n78_port);
   U92 : OAI211_X1 port map( C1 => n79_port, C2 => n80_port, A => n81_port, B 
                           => n82_port, ZN => N210);
   U93 : AOI22_X1 port map( A1 => N49, A2 => n6, B1 => N81, B2 => n5, ZN => 
                           n82_port);
   U94 : OAI21_X1 port map( B1 => n16, B2 => n83_port, A => DATA2(20), ZN => 
                           n81_port);
   U95 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(20), Z => n83_port);
   U96 : INV_X1 port map( A => DATA1(20), ZN => n80_port);
   U97 : AOI21_X1 port map( B1 => n8, B2 => n84_port, A => n16, ZN => n79_port)
                           ;
   U98 : INV_X1 port map( A => DATA2(20), ZN => n84_port);
   U99 : OAI211_X1 port map( C1 => n85_port, C2 => n86_port, A => n87_port, B 
                           => n88_port, ZN => N209);
   U100 : AOI22_X1 port map( A1 => N48, A2 => n6, B1 => N80, B2 => n5, ZN => 
                           n88_port);
   U101 : OAI21_X1 port map( B1 => n16, B2 => n89_port, A => DATA2(19), ZN => 
                           n87_port);
   U102 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(19), Z => n89_port);
   U103 : INV_X1 port map( A => DATA1(19), ZN => n86_port);
   U104 : AOI21_X1 port map( B1 => n8, B2 => n90_port, A => n16, ZN => n85_port
                           );
   U105 : INV_X1 port map( A => DATA2(19), ZN => n90_port);
   U106 : OAI211_X1 port map( C1 => n91_port, C2 => n92_port, A => n93, B => 
                           n94, ZN => N208);
   U107 : AOI22_X1 port map( A1 => N47, A2 => n6, B1 => N79, B2 => n5, ZN => 
                           n94);
   U108 : OAI21_X1 port map( B1 => n16, B2 => n95, A => DATA2(18), ZN => n93);
   U109 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(18), Z => n95);
   U110 : INV_X1 port map( A => DATA1(18), ZN => n92_port);
   U111 : AOI21_X1 port map( B1 => n8, B2 => n96, A => n16, ZN => n91_port);
   U112 : INV_X1 port map( A => DATA2(18), ZN => n96);
   U113 : OAI211_X1 port map( C1 => n97, C2 => n98, A => n99, B => n100, ZN => 
                           N207);
   U114 : AOI22_X1 port map( A1 => N46, A2 => n6, B1 => N78, B2 => n5, ZN => 
                           n100);
   U115 : OAI21_X1 port map( B1 => n16, B2 => n101, A => DATA2(17), ZN => n99);
   U116 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(17), Z => n101);
   U117 : INV_X1 port map( A => DATA1(17), ZN => n98);
   U118 : AOI21_X1 port map( B1 => n8, B2 => n102, A => n16, ZN => n97);
   U119 : INV_X1 port map( A => DATA2(17), ZN => n102);
   U120 : OAI211_X1 port map( C1 => n103, C2 => n104, A => n105, B => n106, ZN 
                           => N206);
   U121 : AOI22_X1 port map( A1 => N45, A2 => n6, B1 => N77, B2 => n5, ZN => 
                           n106);
   U122 : OAI21_X1 port map( B1 => n16, B2 => n107, A => DATA2(16), ZN => n105)
                           ;
   U123 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(16), Z => n107);
   U124 : INV_X1 port map( A => DATA1(16), ZN => n104);
   U125 : AOI21_X1 port map( B1 => n8, B2 => n108, A => n16, ZN => n103);
   U126 : INV_X1 port map( A => DATA2(16), ZN => n108);
   U127 : OAI211_X1 port map( C1 => n109, C2 => n110, A => n111, B => n112, ZN 
                           => N205);
   U128 : AOI22_X1 port map( A1 => N44, A2 => n6, B1 => N76, B2 => n5, ZN => 
                           n112);
   U129 : OAI21_X1 port map( B1 => n16, B2 => n113, A => DATA2(15), ZN => n111)
                           ;
   U130 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(15), Z => n113);
   U131 : INV_X1 port map( A => DATA1(15), ZN => n110);
   U132 : AOI21_X1 port map( B1 => n8, B2 => n114, A => n16, ZN => n109);
   U133 : INV_X1 port map( A => DATA2(15), ZN => n114);
   U134 : OAI211_X1 port map( C1 => n115, C2 => n116, A => n117, B => n118, ZN 
                           => N204);
   U135 : AOI22_X1 port map( A1 => N43, A2 => n6, B1 => N75, B2 => n5, ZN => 
                           n118);
   U136 : OAI21_X1 port map( B1 => n16, B2 => n119, A => DATA2(14), ZN => n117)
                           ;
   U137 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(14), Z => n119);
   U138 : INV_X1 port map( A => DATA1(14), ZN => n116);
   U139 : AOI21_X1 port map( B1 => n8, B2 => n120, A => n16, ZN => n115);
   U140 : INV_X1 port map( A => DATA2(14), ZN => n120);
   U141 : OAI211_X1 port map( C1 => n121, C2 => n122, A => n123, B => n124, ZN 
                           => N203);
   U142 : AOI22_X1 port map( A1 => N42, A2 => n6, B1 => N74, B2 => n5, ZN => 
                           n124);
   U143 : OAI21_X1 port map( B1 => n16, B2 => n125, A => DATA2(13), ZN => n123)
                           ;
   U144 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(13), Z => n125);
   U145 : INV_X1 port map( A => DATA1(13), ZN => n122);
   U146 : AOI21_X1 port map( B1 => n8, B2 => n126, A => n16, ZN => n121);
   U147 : INV_X1 port map( A => DATA2(13), ZN => n126);
   U148 : OAI211_X1 port map( C1 => n127, C2 => n128, A => n129, B => n130, ZN 
                           => N202);
   U149 : AOI22_X1 port map( A1 => N41, A2 => n6, B1 => N73, B2 => n5, ZN => 
                           n130);
   U150 : OAI21_X1 port map( B1 => n16, B2 => n131, A => DATA2(12), ZN => n129)
                           ;
   U151 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(12), Z => n131);
   U152 : INV_X1 port map( A => DATA1(12), ZN => n128);
   U153 : AOI21_X1 port map( B1 => n8, B2 => n132, A => n16, ZN => n127);
   U154 : INV_X1 port map( A => DATA2(12), ZN => n132);
   U155 : OAI211_X1 port map( C1 => n133, C2 => n134, A => n135, B => n136, ZN 
                           => N201);
   U156 : AOI22_X1 port map( A1 => N40, A2 => n6, B1 => N72, B2 => n5, ZN => 
                           n136);
   U157 : OAI21_X1 port map( B1 => n16, B2 => n137, A => DATA2(11), ZN => n135)
                           ;
   U158 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(11), Z => n137);
   U159 : INV_X1 port map( A => DATA1(11), ZN => n134);
   U160 : AOI21_X1 port map( B1 => n8, B2 => n138, A => n16, ZN => n133);
   U161 : INV_X1 port map( A => DATA2(11), ZN => n138);
   U162 : OAI211_X1 port map( C1 => n139, C2 => n140, A => n141, B => n142, ZN 
                           => N200);
   U163 : AOI22_X1 port map( A1 => N39, A2 => n6, B1 => N71, B2 => n5, ZN => 
                           n142);
   U164 : OAI21_X1 port map( B1 => n16, B2 => n143, A => DATA2(10), ZN => n141)
                           ;
   U165 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(10), Z => n143);
   U166 : INV_X1 port map( A => DATA1(10), ZN => n140);
   U167 : AOI21_X1 port map( B1 => n8, B2 => n144, A => n16, ZN => n139);
   U168 : INV_X1 port map( A => DATA2(10), ZN => n144);
   U169 : OAI211_X1 port map( C1 => n145, C2 => n146, A => n147, B => n148, ZN 
                           => N199);
   U170 : AOI22_X1 port map( A1 => N38, A2 => n6, B1 => N70, B2 => n5, ZN => 
                           n148);
   U171 : OAI21_X1 port map( B1 => n16, B2 => n149, A => DATA2(9), ZN => n147);
   U172 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(9), Z => n149);
   U173 : INV_X1 port map( A => DATA1(9), ZN => n146);
   U174 : AOI21_X1 port map( B1 => n8, B2 => n150, A => n16, ZN => n145);
   U175 : INV_X1 port map( A => DATA2(9), ZN => n150);
   U176 : OAI211_X1 port map( C1 => n151, C2 => n152, A => n153, B => n154, ZN 
                           => N198);
   U177 : AOI22_X1 port map( A1 => N37, A2 => n6, B1 => N69, B2 => n5, ZN => 
                           n154);
   U178 : OAI21_X1 port map( B1 => n16, B2 => n155, A => DATA2(8), ZN => n153);
   U179 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(8), Z => n155);
   U180 : INV_X1 port map( A => DATA1(8), ZN => n152);
   U181 : AOI21_X1 port map( B1 => n8, B2 => n156, A => n16, ZN => n151);
   U182 : INV_X1 port map( A => DATA2(8), ZN => n156);
   U183 : OAI211_X1 port map( C1 => n157, C2 => n158, A => n159, B => n160, ZN 
                           => N197);
   U184 : AOI22_X1 port map( A1 => N36, A2 => n6, B1 => N68, B2 => n5, ZN => 
                           n160);
   U185 : OAI21_X1 port map( B1 => n16, B2 => n161, A => DATA2(7), ZN => n159);
   U186 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(7), Z => n161);
   U187 : INV_X1 port map( A => DATA1(7), ZN => n158);
   U188 : AOI21_X1 port map( B1 => n8, B2 => n162, A => n16, ZN => n157);
   U189 : INV_X1 port map( A => DATA2(7), ZN => n162);
   U190 : OAI211_X1 port map( C1 => n163, C2 => n164, A => n165, B => n166, ZN 
                           => N196);
   U191 : AOI22_X1 port map( A1 => N35, A2 => n6, B1 => N67, B2 => n5, ZN => 
                           n166);
   U192 : OAI21_X1 port map( B1 => n16, B2 => n167, A => DATA2(6), ZN => n165);
   U193 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(6), Z => n167);
   U194 : INV_X1 port map( A => DATA1(6), ZN => n164);
   U195 : AOI21_X1 port map( B1 => n8, B2 => n168, A => n16, ZN => n163);
   U196 : INV_X1 port map( A => DATA2(6), ZN => n168);
   U197 : OAI211_X1 port map( C1 => n169, C2 => n170, A => n171, B => n172, ZN 
                           => N195);
   U198 : AOI22_X1 port map( A1 => N34, A2 => n6, B1 => N66, B2 => n5, ZN => 
                           n172);
   U199 : OAI21_X1 port map( B1 => n16, B2 => n173, A => DATA2(5), ZN => n171);
   U200 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(5), Z => n173);
   U201 : INV_X1 port map( A => DATA1(5), ZN => n170);
   U202 : AOI21_X1 port map( B1 => n8, B2 => n174, A => n16, ZN => n169);
   U203 : INV_X1 port map( A => DATA2(5), ZN => n174);
   U204 : OAI211_X1 port map( C1 => n175, C2 => n176, A => n177, B => n178, ZN 
                           => N194);
   U205 : AOI22_X1 port map( A1 => N33, A2 => n6, B1 => N65, B2 => n5, ZN => 
                           n178);
   U206 : OAI21_X1 port map( B1 => n16, B2 => n179, A => DATA2(4), ZN => n177);
   U207 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(4), Z => n179);
   U208 : INV_X1 port map( A => DATA1(4), ZN => n176);
   U209 : AOI21_X1 port map( B1 => n8, B2 => n180, A => n16, ZN => n175);
   U210 : INV_X1 port map( A => DATA2(4), ZN => n180);
   U211 : OAI211_X1 port map( C1 => n181, C2 => n182, A => n183, B => n184, ZN 
                           => N193);
   U212 : AOI22_X1 port map( A1 => N32, A2 => n6, B1 => N64, B2 => n5, ZN => 
                           n184);
   U213 : OAI21_X1 port map( B1 => n16, B2 => n185, A => DATA2(3), ZN => n183);
   U214 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(3), Z => n185);
   U215 : INV_X1 port map( A => DATA1(3), ZN => n182);
   U216 : AOI21_X1 port map( B1 => n8, B2 => n186, A => n16, ZN => n181);
   U217 : INV_X1 port map( A => DATA2(3), ZN => n186);
   U218 : OAI211_X1 port map( C1 => n187, C2 => n188, A => n189, B => n190_port
                           , ZN => N192);
   U219 : AOI22_X1 port map( A1 => N31, A2 => n6, B1 => N63, B2 => n5, ZN => 
                           n190_port);
   U220 : OAI21_X1 port map( B1 => n16, B2 => n191_port, A => DATA2(2), ZN => 
                           n189);
   U221 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(2), Z => n191_port);
   U222 : INV_X1 port map( A => DATA1(2), ZN => n188);
   U223 : AOI21_X1 port map( B1 => n8, B2 => n192_port, A => n16, ZN => n187);
   U224 : INV_X1 port map( A => DATA2(2), ZN => n192_port);
   U225 : OAI211_X1 port map( C1 => n193_port, C2 => n194_port, A => n195_port,
                           B => n196_port, ZN => N191);
   U226 : AOI22_X1 port map( A1 => N30, A2 => n6, B1 => N62, B2 => n5, ZN => 
                           n196_port);
   U227 : OAI21_X1 port map( B1 => n16, B2 => n197_port, A => DATA2(1), ZN => 
                           n195_port);
   U228 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(1), Z => n197_port);
   U229 : INV_X1 port map( A => DATA1(1), ZN => n194_port);
   U230 : AOI21_X1 port map( B1 => n8, B2 => n198_port, A => n16, ZN => 
                           n193_port);
   U231 : INV_X1 port map( A => DATA2(1), ZN => n198_port);
   U232 : OAI211_X1 port map( C1 => n199_port, C2 => n200_port, A => n201_port,
                           B => n202_port, ZN => N190);
   U233 : AOI22_X1 port map( A1 => N29, A2 => n6, B1 => N61, B2 => n5, ZN => 
                           n202_port);
   U234 : OAI21_X1 port map( B1 => n16, B2 => n204_port, A => DATA2(0), ZN => 
                           n201_port);
   U235 : MUX2_X1 port map( A => n8, B => n9, S => DATA1(0), Z => n204_port);
   U236 : INV_X1 port map( A => DATA1(0), ZN => n200_port);
   U237 : AOI21_X1 port map( B1 => n8, B2 => n205_port, A => n16, ZN => 
                           n199_port);
   U238 : INV_X1 port map( A => FUNC(1), ZN => n206_port);
   U239 : INV_X1 port map( A => DATA2(0), ZN => n205_port);
   U240 : INV_X1 port map( A => FUNC(3), ZN => n203_port);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity P4_ADDER_NBITS32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end P4_ADDER_NBITS32;

architecture SYN_STRUCTURAL of P4_ADDER_NBITS32 is

   component CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4
      port( A, B : in std_logic_vector (32 downto 1);  C0 : in std_logic;  COUT
            : out std_logic_vector (8 downto 0));
   end component;
   
   component SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (8 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component xor_logic_nbits32
      port( Cin : in std_logic;  B0 : in std_logic_vector (31 downto 0);  B : 
            out std_logic_vector (31 downto 0));
   end component;
   
   signal Co_port, B_diff_31_port, B_diff_30_port, B_diff_29_port, 
      B_diff_28_port, B_diff_27_port, B_diff_26_port, B_diff_25_port, 
      B_diff_24_port, B_diff_23_port, B_diff_22_port, B_diff_21_port, 
      B_diff_20_port, B_diff_19_port, B_diff_18_port, B_diff_17_port, 
      B_diff_16_port, B_diff_15_port, B_diff_14_port, B_diff_13_port, 
      B_diff_12_port, B_diff_11_port, B_diff_10_port, B_diff_9_port, 
      B_diff_8_port, B_diff_7_port, B_diff_6_port, B_diff_5_port, B_diff_4_port
      , B_diff_3_port, B_diff_2_port, B_diff_1_port, B_diff_0_port, 
      fromCarry_to_adder_7_port, fromCarry_to_adder_6_port, 
      fromCarry_to_adder_5_port, fromCarry_to_adder_4_port, 
      fromCarry_to_adder_3_port, fromCarry_to_adder_2_port, 
      fromCarry_to_adder_1_port, fromCarry_to_adder_0_port : std_logic;

begin
   Co <= Co_port;
   
   xor_gate : xor_logic_nbits32 port map( Cin => Ci, B0(31) => B(31), B0(30) =>
                           B(30), B0(29) => B(29), B0(28) => B(28), B0(27) => 
                           B(27), B0(26) => B(26), B0(25) => B(25), B0(24) => 
                           B(24), B0(23) => B(23), B0(22) => B(22), B0(21) => 
                           B(21), B0(20) => B(20), B0(19) => B(19), B0(18) => 
                           B(18), B0(17) => B(17), B0(16) => B(16), B0(15) => 
                           B(15), B0(14) => B(14), B0(13) => B(13), B0(12) => 
                           B(12), B0(11) => B(11), B0(10) => B(10), B0(9) => 
                           B(9), B0(8) => B(8), B0(7) => B(7), B0(6) => B(6), 
                           B0(5) => B(5), B0(4) => B(4), B0(3) => B(3), B0(2) 
                           => B(2), B0(1) => B(1), B0(0) => B(0), B(31) => 
                           B_diff_31_port, B(30) => B_diff_30_port, B(29) => 
                           B_diff_29_port, B(28) => B_diff_28_port, B(27) => 
                           B_diff_27_port, B(26) => B_diff_26_port, B(25) => 
                           B_diff_25_port, B(24) => B_diff_24_port, B(23) => 
                           B_diff_23_port, B(22) => B_diff_22_port, B(21) => 
                           B_diff_21_port, B(20) => B_diff_20_port, B(19) => 
                           B_diff_19_port, B(18) => B_diff_18_port, B(17) => 
                           B_diff_17_port, B(16) => B_diff_16_port, B(15) => 
                           B_diff_15_port, B(14) => B_diff_14_port, B(13) => 
                           B_diff_13_port, B(12) => B_diff_12_port, B(11) => 
                           B_diff_11_port, B(10) => B_diff_10_port, B(9) => 
                           B_diff_9_port, B(8) => B_diff_8_port, B(7) => 
                           B_diff_7_port, B(6) => B_diff_6_port, B(5) => 
                           B_diff_5_port, B(4) => B_diff_4_port, B(3) => 
                           B_diff_3_port, B(2) => B_diff_2_port, B(1) => 
                           B_diff_1_port, B(0) => B_diff_0_port);
   SUM_GEN : SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8 port map( A(31)
                           => A(31), A(30) => A(30), A(29) => A(29), A(28) => 
                           A(28), A(27) => A(27), A(26) => A(26), A(25) => 
                           A(25), A(24) => A(24), A(23) => A(23), A(22) => 
                           A(22), A(21) => A(21), A(20) => A(20), A(19) => 
                           A(19), A(18) => A(18), A(17) => A(17), A(16) => 
                           A(16), A(15) => A(15), A(14) => A(14), A(13) => 
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => B_diff_31_port, B(30) => B_diff_30_port, 
                           B(29) => B_diff_29_port, B(28) => B_diff_28_port, 
                           B(27) => B_diff_27_port, B(26) => B_diff_26_port, 
                           B(25) => B_diff_25_port, B(24) => B_diff_24_port, 
                           B(23) => B_diff_23_port, B(22) => B_diff_22_port, 
                           B(21) => B_diff_21_port, B(20) => B_diff_20_port, 
                           B(19) => B_diff_19_port, B(18) => B_diff_18_port, 
                           B(17) => B_diff_17_port, B(16) => B_diff_16_port, 
                           B(15) => B_diff_15_port, B(14) => B_diff_14_port, 
                           B(13) => B_diff_13_port, B(12) => B_diff_12_port, 
                           B(11) => B_diff_11_port, B(10) => B_diff_10_port, 
                           B(9) => B_diff_9_port, B(8) => B_diff_8_port, B(7) 
                           => B_diff_7_port, B(6) => B_diff_6_port, B(5) => 
                           B_diff_5_port, B(4) => B_diff_4_port, B(3) => 
                           B_diff_3_port, B(2) => B_diff_2_port, B(1) => 
                           B_diff_1_port, B(0) => B_diff_0_port, Ci(8) => 
                           Co_port, Ci(7) => fromCarry_to_adder_7_port, Ci(6) 
                           => fromCarry_to_adder_6_port, Ci(5) => 
                           fromCarry_to_adder_5_port, Ci(4) => 
                           fromCarry_to_adder_4_port, Ci(3) => 
                           fromCarry_to_adder_3_port, Ci(2) => 
                           fromCarry_to_adder_2_port, Ci(1) => 
                           fromCarry_to_adder_1_port, Ci(0) => 
                           fromCarry_to_adder_0_port, S(31) => S(31), S(30) => 
                           S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));
   CLA : CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4 port map( A(32) => A(31), A(31)
                           => A(30), A(30) => A(29), A(29) => A(28), A(28) => 
                           A(27), A(27) => A(26), A(26) => A(25), A(25) => 
                           A(24), A(24) => A(23), A(23) => A(22), A(22) => 
                           A(21), A(21) => A(20), A(20) => A(19), A(19) => 
                           A(18), A(18) => A(17), A(17) => A(16), A(16) => 
                           A(15), A(15) => A(14), A(14) => A(13), A(13) => 
                           A(12), A(12) => A(11), A(11) => A(10), A(10) => A(9)
                           , A(9) => A(8), A(8) => A(7), A(7) => A(6), A(6) => 
                           A(5), A(5) => A(4), A(4) => A(3), A(3) => A(2), A(2)
                           => A(1), A(1) => A(0), B(32) => B_diff_31_port, 
                           B(31) => B_diff_30_port, B(30) => B_diff_29_port, 
                           B(29) => B_diff_28_port, B(28) => B_diff_27_port, 
                           B(27) => B_diff_26_port, B(26) => B_diff_25_port, 
                           B(25) => B_diff_24_port, B(24) => B_diff_23_port, 
                           B(23) => B_diff_22_port, B(22) => B_diff_21_port, 
                           B(21) => B_diff_20_port, B(20) => B_diff_19_port, 
                           B(19) => B_diff_18_port, B(18) => B_diff_17_port, 
                           B(17) => B_diff_16_port, B(16) => B_diff_15_port, 
                           B(15) => B_diff_14_port, B(14) => B_diff_13_port, 
                           B(13) => B_diff_12_port, B(12) => B_diff_11_port, 
                           B(11) => B_diff_10_port, B(10) => B_diff_9_port, 
                           B(9) => B_diff_8_port, B(8) => B_diff_7_port, B(7) 
                           => B_diff_6_port, B(6) => B_diff_5_port, B(5) => 
                           B_diff_4_port, B(4) => B_diff_3_port, B(3) => 
                           B_diff_2_port, B(2) => B_diff_1_port, B(1) => 
                           B_diff_0_port, C0 => Ci, COUT(8) => Co_port, COUT(7)
                           => fromCarry_to_adder_7_port, COUT(6) => 
                           fromCarry_to_adder_6_port, COUT(5) => 
                           fromCarry_to_adder_5_port, COUT(4) => 
                           fromCarry_to_adder_4_port, COUT(3) => 
                           fromCarry_to_adder_3_port, COUT(2) => 
                           fromCarry_to_adder_2_port, COUT(1) => 
                           fromCarry_to_adder_1_port, COUT(0) => 
                           fromCarry_to_adder_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ctrl_alu_NBITS32 is

   port( A, B : in std_logic_vector (31 downto 0);  FUNC : in std_logic_vector 
         (0 to 3);  Ap4, Bp4 : out std_logic_vector (31 downto 0);  Cin : out 
         std_logic;  Als, Bls : out std_logic_vector (31 downto 0);  enableComp
         : out std_logic);

end ctrl_alu_NBITS32;

architecture SYN_BEHAVIORAL of ctrl_alu_NBITS32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76 : std_logic;

begin
   
   U3 : OAI21_X1 port map( B1 => n2, B2 => n3, A => n4, ZN => n76);
   U4 : AND2_X4 port map( A1 => n4, A2 => n2, ZN => n5);
   U5 : NAND2_X4 port map( A1 => n72, A2 => n75, ZN => n38);
   U6 : CLKBUF_X2 port map( A => n76, Z => Cin);
   U7 : INV_X1 port map( A => FUNC(3), ZN => n3);
   U8 : INV_X1 port map( A => n4, ZN => enableComp);
   U9 : NOR2_X1 port map( A1 => n5, A2 => n6, ZN => Bp4(9));
   U10 : NOR2_X1 port map( A1 => n5, A2 => n7, ZN => Bp4(8));
   U11 : NOR2_X1 port map( A1 => n5, A2 => n8, ZN => Bp4(7));
   U12 : NOR2_X1 port map( A1 => n5, A2 => n9, ZN => Bp4(6));
   U13 : NOR2_X1 port map( A1 => n5, A2 => n10, ZN => Bp4(5));
   U14 : NOR2_X1 port map( A1 => n5, A2 => n11, ZN => Bp4(4));
   U15 : NOR2_X1 port map( A1 => n5, A2 => n12, ZN => Bp4(3));
   U16 : NOR2_X1 port map( A1 => n5, A2 => n13, ZN => Bp4(31));
   U17 : NOR2_X1 port map( A1 => n5, A2 => n14, ZN => Bp4(30));
   U18 : NOR2_X1 port map( A1 => n5, A2 => n15, ZN => Bp4(2));
   U19 : NOR2_X1 port map( A1 => n5, A2 => n16, ZN => Bp4(29));
   U20 : NOR2_X1 port map( A1 => n5, A2 => n17, ZN => Bp4(28));
   U21 : NOR2_X1 port map( A1 => n5, A2 => n18, ZN => Bp4(27));
   U22 : NOR2_X1 port map( A1 => n5, A2 => n19, ZN => Bp4(26));
   U23 : NOR2_X1 port map( A1 => n5, A2 => n20, ZN => Bp4(25));
   U24 : NOR2_X1 port map( A1 => n5, A2 => n21, ZN => Bp4(24));
   U25 : NOR2_X1 port map( A1 => n5, A2 => n22, ZN => Bp4(23));
   U26 : NOR2_X1 port map( A1 => n5, A2 => n23, ZN => Bp4(22));
   U27 : NOR2_X1 port map( A1 => n5, A2 => n24, ZN => Bp4(21));
   U28 : NOR2_X1 port map( A1 => n5, A2 => n25, ZN => Bp4(20));
   U29 : NOR2_X1 port map( A1 => n5, A2 => n26, ZN => Bp4(1));
   U30 : NOR2_X1 port map( A1 => n5, A2 => n27, ZN => Bp4(19));
   U31 : NOR2_X1 port map( A1 => n5, A2 => n28, ZN => Bp4(18));
   U32 : NOR2_X1 port map( A1 => n5, A2 => n29, ZN => Bp4(17));
   U33 : NOR2_X1 port map( A1 => n5, A2 => n30, ZN => Bp4(16));
   U34 : NOR2_X1 port map( A1 => n5, A2 => n31, ZN => Bp4(15));
   U35 : NOR2_X1 port map( A1 => n5, A2 => n32, ZN => Bp4(14));
   U36 : NOR2_X1 port map( A1 => n5, A2 => n33, ZN => Bp4(13));
   U37 : NOR2_X1 port map( A1 => n5, A2 => n34, ZN => Bp4(12));
   U38 : NOR2_X1 port map( A1 => n5, A2 => n35, ZN => Bp4(11));
   U39 : NOR2_X1 port map( A1 => n5, A2 => n36, ZN => Bp4(10));
   U40 : NOR2_X1 port map( A1 => n5, A2 => n37, ZN => Bp4(0));
   U41 : NOR2_X1 port map( A1 => n6, A2 => n38, ZN => Bls(9));
   U42 : INV_X1 port map( A => B(9), ZN => n6);
   U43 : NOR2_X1 port map( A1 => n7, A2 => n38, ZN => Bls(8));
   U44 : INV_X1 port map( A => B(8), ZN => n7);
   U45 : NOR2_X1 port map( A1 => n8, A2 => n38, ZN => Bls(7));
   U46 : INV_X1 port map( A => B(7), ZN => n8);
   U47 : NOR2_X1 port map( A1 => n9, A2 => n38, ZN => Bls(6));
   U48 : INV_X1 port map( A => B(6), ZN => n9);
   U49 : NOR2_X1 port map( A1 => n10, A2 => n38, ZN => Bls(5));
   U50 : INV_X1 port map( A => B(5), ZN => n10);
   U51 : NOR2_X1 port map( A1 => n11, A2 => n38, ZN => Bls(4));
   U52 : INV_X1 port map( A => B(4), ZN => n11);
   U53 : NOR2_X1 port map( A1 => n12, A2 => n38, ZN => Bls(3));
   U54 : INV_X1 port map( A => B(3), ZN => n12);
   U55 : NOR2_X1 port map( A1 => n13, A2 => n38, ZN => Bls(31));
   U56 : INV_X1 port map( A => B(31), ZN => n13);
   U57 : NOR2_X1 port map( A1 => n14, A2 => n38, ZN => Bls(30));
   U58 : INV_X1 port map( A => B(30), ZN => n14);
   U59 : NOR2_X1 port map( A1 => n15, A2 => n38, ZN => Bls(2));
   U60 : INV_X1 port map( A => B(2), ZN => n15);
   U61 : NOR2_X1 port map( A1 => n16, A2 => n38, ZN => Bls(29));
   U62 : INV_X1 port map( A => B(29), ZN => n16);
   U63 : NOR2_X1 port map( A1 => n17, A2 => n38, ZN => Bls(28));
   U64 : INV_X1 port map( A => B(28), ZN => n17);
   U65 : NOR2_X1 port map( A1 => n18, A2 => n38, ZN => Bls(27));
   U66 : INV_X1 port map( A => B(27), ZN => n18);
   U67 : NOR2_X1 port map( A1 => n19, A2 => n38, ZN => Bls(26));
   U68 : INV_X1 port map( A => B(26), ZN => n19);
   U69 : NOR2_X1 port map( A1 => n20, A2 => n38, ZN => Bls(25));
   U70 : INV_X1 port map( A => B(25), ZN => n20);
   U71 : NOR2_X1 port map( A1 => n21, A2 => n38, ZN => Bls(24));
   U72 : INV_X1 port map( A => B(24), ZN => n21);
   U73 : NOR2_X1 port map( A1 => n22, A2 => n38, ZN => Bls(23));
   U74 : INV_X1 port map( A => B(23), ZN => n22);
   U75 : NOR2_X1 port map( A1 => n23, A2 => n38, ZN => Bls(22));
   U76 : INV_X1 port map( A => B(22), ZN => n23);
   U77 : NOR2_X1 port map( A1 => n24, A2 => n38, ZN => Bls(21));
   U78 : INV_X1 port map( A => B(21), ZN => n24);
   U79 : NOR2_X1 port map( A1 => n25, A2 => n38, ZN => Bls(20));
   U80 : INV_X1 port map( A => B(20), ZN => n25);
   U81 : NOR2_X1 port map( A1 => n26, A2 => n38, ZN => Bls(1));
   U82 : INV_X1 port map( A => B(1), ZN => n26);
   U83 : NOR2_X1 port map( A1 => n27, A2 => n38, ZN => Bls(19));
   U84 : INV_X1 port map( A => B(19), ZN => n27);
   U85 : NOR2_X1 port map( A1 => n28, A2 => n38, ZN => Bls(18));
   U86 : INV_X1 port map( A => B(18), ZN => n28);
   U87 : NOR2_X1 port map( A1 => n29, A2 => n38, ZN => Bls(17));
   U88 : INV_X1 port map( A => B(17), ZN => n29);
   U89 : NOR2_X1 port map( A1 => n30, A2 => n38, ZN => Bls(16));
   U90 : INV_X1 port map( A => B(16), ZN => n30);
   U91 : NOR2_X1 port map( A1 => n31, A2 => n38, ZN => Bls(15));
   U92 : INV_X1 port map( A => B(15), ZN => n31);
   U93 : NOR2_X1 port map( A1 => n32, A2 => n38, ZN => Bls(14));
   U94 : INV_X1 port map( A => B(14), ZN => n32);
   U95 : NOR2_X1 port map( A1 => n33, A2 => n38, ZN => Bls(13));
   U96 : INV_X1 port map( A => B(13), ZN => n33);
   U97 : NOR2_X1 port map( A1 => n34, A2 => n38, ZN => Bls(12));
   U98 : INV_X1 port map( A => B(12), ZN => n34);
   U99 : NOR2_X1 port map( A1 => n35, A2 => n38, ZN => Bls(11));
   U100 : INV_X1 port map( A => B(11), ZN => n35);
   U101 : NOR2_X1 port map( A1 => n36, A2 => n38, ZN => Bls(10));
   U102 : INV_X1 port map( A => B(10), ZN => n36);
   U103 : NOR2_X1 port map( A1 => n37, A2 => n38, ZN => Bls(0));
   U104 : INV_X1 port map( A => B(0), ZN => n37);
   U105 : NOR2_X1 port map( A1 => n5, A2 => n39, ZN => Ap4(9));
   U106 : NOR2_X1 port map( A1 => n5, A2 => n40, ZN => Ap4(8));
   U107 : NOR2_X1 port map( A1 => n5, A2 => n41, ZN => Ap4(7));
   U108 : NOR2_X1 port map( A1 => n5, A2 => n42, ZN => Ap4(6));
   U109 : NOR2_X1 port map( A1 => n5, A2 => n43, ZN => Ap4(5));
   U110 : NOR2_X1 port map( A1 => n5, A2 => n44, ZN => Ap4(4));
   U111 : NOR2_X1 port map( A1 => n5, A2 => n45, ZN => Ap4(3));
   U112 : NOR2_X1 port map( A1 => n5, A2 => n46, ZN => Ap4(31));
   U113 : NOR2_X1 port map( A1 => n5, A2 => n47, ZN => Ap4(30));
   U114 : NOR2_X1 port map( A1 => n5, A2 => n48, ZN => Ap4(2));
   U115 : NOR2_X1 port map( A1 => n5, A2 => n49, ZN => Ap4(29));
   U116 : NOR2_X1 port map( A1 => n5, A2 => n50, ZN => Ap4(28));
   U117 : NOR2_X1 port map( A1 => n5, A2 => n51, ZN => Ap4(27));
   U118 : NOR2_X1 port map( A1 => n5, A2 => n52, ZN => Ap4(26));
   U119 : NOR2_X1 port map( A1 => n5, A2 => n53, ZN => Ap4(25));
   U120 : NOR2_X1 port map( A1 => n5, A2 => n54, ZN => Ap4(24));
   U121 : NOR2_X1 port map( A1 => n5, A2 => n55, ZN => Ap4(23));
   U122 : NOR2_X1 port map( A1 => n5, A2 => n56, ZN => Ap4(22));
   U123 : NOR2_X1 port map( A1 => n5, A2 => n57, ZN => Ap4(21));
   U124 : NOR2_X1 port map( A1 => n5, A2 => n58, ZN => Ap4(20));
   U125 : NOR2_X1 port map( A1 => n5, A2 => n59, ZN => Ap4(1));
   U126 : NOR2_X1 port map( A1 => n5, A2 => n60, ZN => Ap4(19));
   U127 : NOR2_X1 port map( A1 => n5, A2 => n61, ZN => Ap4(18));
   U128 : NOR2_X1 port map( A1 => n5, A2 => n62, ZN => Ap4(17));
   U129 : NOR2_X1 port map( A1 => n5, A2 => n63, ZN => Ap4(16));
   U130 : NOR2_X1 port map( A1 => n5, A2 => n64, ZN => Ap4(15));
   U131 : NOR2_X1 port map( A1 => n5, A2 => n65, ZN => Ap4(14));
   U132 : NOR2_X1 port map( A1 => n5, A2 => n66, ZN => Ap4(13));
   U133 : NOR2_X1 port map( A1 => n5, A2 => n67, ZN => Ap4(12));
   U134 : NOR2_X1 port map( A1 => n5, A2 => n68, ZN => Ap4(11));
   U135 : NOR2_X1 port map( A1 => n5, A2 => n69, ZN => Ap4(10));
   U136 : NOR2_X1 port map( A1 => n5, A2 => n70, ZN => Ap4(0));
   U137 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => FUNC(2), ZN => n2);
   U138 : MUX2_X1 port map( A => n73, B => n74, S => n71, Z => n4);
   U139 : OR2_X1 port map( A1 => n72, A2 => FUNC(2), ZN => n74);
   U140 : NAND3_X1 port map( A1 => FUNC(2), A2 => n72, A3 => FUNC(3), ZN => n73
                           );
   U141 : NOR2_X1 port map( A1 => n38, A2 => n39, ZN => Als(9));
   U142 : INV_X1 port map( A => A(9), ZN => n39);
   U143 : NOR2_X1 port map( A1 => n38, A2 => n40, ZN => Als(8));
   U144 : INV_X1 port map( A => A(8), ZN => n40);
   U145 : NOR2_X1 port map( A1 => n38, A2 => n41, ZN => Als(7));
   U146 : INV_X1 port map( A => A(7), ZN => n41);
   U147 : NOR2_X1 port map( A1 => n38, A2 => n42, ZN => Als(6));
   U148 : INV_X1 port map( A => A(6), ZN => n42);
   U149 : NOR2_X1 port map( A1 => n38, A2 => n43, ZN => Als(5));
   U150 : INV_X1 port map( A => A(5), ZN => n43);
   U151 : NOR2_X1 port map( A1 => n38, A2 => n44, ZN => Als(4));
   U152 : INV_X1 port map( A => A(4), ZN => n44);
   U153 : NOR2_X1 port map( A1 => n38, A2 => n45, ZN => Als(3));
   U154 : INV_X1 port map( A => A(3), ZN => n45);
   U155 : NOR2_X1 port map( A1 => n38, A2 => n46, ZN => Als(31));
   U156 : INV_X1 port map( A => A(31), ZN => n46);
   U157 : NOR2_X1 port map( A1 => n38, A2 => n47, ZN => Als(30));
   U158 : INV_X1 port map( A => A(30), ZN => n47);
   U159 : NOR2_X1 port map( A1 => n38, A2 => n48, ZN => Als(2));
   U160 : INV_X1 port map( A => A(2), ZN => n48);
   U161 : NOR2_X1 port map( A1 => n38, A2 => n49, ZN => Als(29));
   U162 : INV_X1 port map( A => A(29), ZN => n49);
   U163 : NOR2_X1 port map( A1 => n38, A2 => n50, ZN => Als(28));
   U164 : INV_X1 port map( A => A(28), ZN => n50);
   U165 : NOR2_X1 port map( A1 => n38, A2 => n51, ZN => Als(27));
   U166 : INV_X1 port map( A => A(27), ZN => n51);
   U167 : NOR2_X1 port map( A1 => n38, A2 => n52, ZN => Als(26));
   U168 : INV_X1 port map( A => A(26), ZN => n52);
   U169 : NOR2_X1 port map( A1 => n38, A2 => n53, ZN => Als(25));
   U170 : INV_X1 port map( A => A(25), ZN => n53);
   U171 : NOR2_X1 port map( A1 => n38, A2 => n54, ZN => Als(24));
   U172 : INV_X1 port map( A => A(24), ZN => n54);
   U173 : NOR2_X1 port map( A1 => n38, A2 => n55, ZN => Als(23));
   U174 : INV_X1 port map( A => A(23), ZN => n55);
   U175 : NOR2_X1 port map( A1 => n38, A2 => n56, ZN => Als(22));
   U176 : INV_X1 port map( A => A(22), ZN => n56);
   U177 : NOR2_X1 port map( A1 => n38, A2 => n57, ZN => Als(21));
   U178 : INV_X1 port map( A => A(21), ZN => n57);
   U179 : NOR2_X1 port map( A1 => n38, A2 => n58, ZN => Als(20));
   U180 : INV_X1 port map( A => A(20), ZN => n58);
   U181 : NOR2_X1 port map( A1 => n38, A2 => n59, ZN => Als(1));
   U182 : INV_X1 port map( A => A(1), ZN => n59);
   U183 : NOR2_X1 port map( A1 => n38, A2 => n60, ZN => Als(19));
   U184 : INV_X1 port map( A => A(19), ZN => n60);
   U185 : NOR2_X1 port map( A1 => n38, A2 => n61, ZN => Als(18));
   U186 : INV_X1 port map( A => A(18), ZN => n61);
   U187 : NOR2_X1 port map( A1 => n38, A2 => n62, ZN => Als(17));
   U188 : INV_X1 port map( A => A(17), ZN => n62);
   U189 : NOR2_X1 port map( A1 => n38, A2 => n63, ZN => Als(16));
   U190 : INV_X1 port map( A => A(16), ZN => n63);
   U191 : NOR2_X1 port map( A1 => n38, A2 => n64, ZN => Als(15));
   U192 : INV_X1 port map( A => A(15), ZN => n64);
   U193 : NOR2_X1 port map( A1 => n38, A2 => n65, ZN => Als(14));
   U194 : INV_X1 port map( A => A(14), ZN => n65);
   U195 : NOR2_X1 port map( A1 => n38, A2 => n66, ZN => Als(13));
   U196 : INV_X1 port map( A => A(13), ZN => n66);
   U197 : NOR2_X1 port map( A1 => n38, A2 => n67, ZN => Als(12));
   U198 : INV_X1 port map( A => A(12), ZN => n67);
   U199 : NOR2_X1 port map( A1 => n38, A2 => n68, ZN => Als(11));
   U200 : INV_X1 port map( A => A(11), ZN => n68);
   U201 : NOR2_X1 port map( A1 => n38, A2 => n69, ZN => Als(10));
   U202 : INV_X1 port map( A => A(10), ZN => n69);
   U203 : NOR2_X1 port map( A1 => n38, A2 => n70, ZN => Als(0));
   U204 : INV_X1 port map( A => A(0), ZN => n70);
   U205 : OAI21_X1 port map( B1 => FUNC(3), B2 => n71, A => FUNC(2), ZN => n75)
                           ;
   U206 : INV_X1 port map( A => FUNC(1), ZN => n71);
   U207 : INV_X1 port map( A => FUNC(0), ZN => n72);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity comparator_bits32 is

   port( Cout, EN : in std_logic;  func : in std_logic_vector (0 to 3);  sum : 
         in std_logic_vector (31 downto 0);  set : out std_logic_vector (31 
         downto 0));

end comparator_bits32;

architecture SYN_BEHAVIORAL of comparator_bits32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, set_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18 : std_logic;

begin
   set <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, set_0_port 
      );
   
   X_Logic0_port <= '0';
   U2 : AND2_X1 port map( A1 => n1, A2 => EN, ZN => set_0_port);
   U3 : MUX2_X1 port map( A => n2, B => n3, S => func(1), Z => n1);
   U4 : AND4_X1 port map( A1 => n4, A2 => n5, A3 => func(3), A4 => func(2), ZN 
                           => n3);
   U5 : INV_X1 port map( A => n6, ZN => n5);
   U6 : NOR3_X1 port map( A1 => n4, A2 => func(2), A3 => n7, ZN => n2);
   U7 : XOR2_X1 port map( A => n8, B => Cout, Z => n7);
   U8 : OR2_X1 port map( A1 => func(3), A2 => n6, ZN => n8);
   U9 : NOR2_X1 port map( A1 => n9, A2 => n10, ZN => n6);
   U10 : NAND4_X1 port map( A1 => n11, A2 => n12, A3 => n13, A4 => n14, ZN => 
                           n10);
   U11 : NOR4_X1 port map( A1 => sum(23), A2 => sum(22), A3 => sum(21), A4 => 
                           sum(20), ZN => n14);
   U12 : NOR4_X1 port map( A1 => sum(1), A2 => sum(19), A3 => sum(18), A4 => 
                           sum(17), ZN => n13);
   U13 : NOR4_X1 port map( A1 => sum(16), A2 => sum(15), A3 => sum(14), A4 => 
                           sum(13), ZN => n12);
   U14 : NOR4_X1 port map( A1 => sum(12), A2 => sum(11), A3 => sum(10), A4 => 
                           sum(0), ZN => n11);
   U15 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           n9);
   U16 : NOR4_X1 port map( A1 => sum(9), A2 => sum(8), A3 => sum(7), A4 => 
                           sum(6), ZN => n18);
   U17 : NOR4_X1 port map( A1 => sum(5), A2 => sum(4), A3 => sum(3), A4 => 
                           sum(31), ZN => n17);
   U18 : NOR4_X1 port map( A1 => sum(30), A2 => sum(2), A3 => sum(29), A4 => 
                           sum(28), ZN => n16);
   U19 : NOR4_X1 port map( A1 => sum(27), A2 => sum(26), A3 => sum(25), A4 => 
                           sum(24), ZN => n15);
   U20 : INV_X1 port map( A => func(0), ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity outputSelect_nbits32 is

   port( FUNC : in std_logic_vector (0 to 3);  p4_out, LS_OUT, comp_out : in 
         std_logic_vector (31 downto 0);  outputSel : out std_logic_vector (31 
         downto 0));

end outputSelect_nbits32;

architecture SYN_BEHAVIORAL of outputSelect_nbits32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43 : 
      std_logic;

begin
   
   U2 : INV_X2 port map( A => n37, ZN => n5);
   U3 : AND2_X2 port map( A1 => n43, A2 => n42, ZN => n4);
   U4 : OR3_X1 port map( A1 => FUNC(1), A2 => FUNC(0), A3 => n41, ZN => n3);
   U5 : INV_X2 port map( A => n3, ZN => n1);
   U6 : INV_X1 port map( A => n2, ZN => outputSel(0));
   U7 : AOI222_X1 port map( A1 => p4_out(0), A2 => n1, B1 => LS_OUT(0), B2 => 
                           n4, C1 => comp_out(0), C2 => n5, ZN => n2);
   U8 : INV_X1 port map( A => n6, ZN => outputSel(5));
   U9 : AOI222_X1 port map( A1 => p4_out(5), A2 => n1, B1 => LS_OUT(5), B2 => 
                           n4, C1 => comp_out(5), C2 => n5, ZN => n6);
   U10 : INV_X1 port map( A => n7, ZN => outputSel(7));
   U11 : AOI222_X1 port map( A1 => p4_out(7), A2 => n1, B1 => LS_OUT(7), B2 => 
                           n4, C1 => comp_out(7), C2 => n5, ZN => n7);
   U12 : INV_X1 port map( A => n8, ZN => outputSel(6));
   U13 : AOI222_X1 port map( A1 => p4_out(6), A2 => n1, B1 => LS_OUT(6), B2 => 
                           n4, C1 => comp_out(6), C2 => n5, ZN => n8);
   U14 : INV_X1 port map( A => n9, ZN => outputSel(4));
   U15 : AOI222_X1 port map( A1 => p4_out(4), A2 => n1, B1 => LS_OUT(4), B2 => 
                           n4, C1 => comp_out(4), C2 => n5, ZN => n9);
   U16 : INV_X1 port map( A => n10, ZN => outputSel(9));
   U17 : AOI222_X1 port map( A1 => p4_out(9), A2 => n1, B1 => LS_OUT(9), B2 => 
                           n4, C1 => comp_out(9), C2 => n5, ZN => n10);
   U18 : INV_X1 port map( A => n11, ZN => outputSel(11));
   U19 : AOI222_X1 port map( A1 => p4_out(11), A2 => n1, B1 => LS_OUT(11), B2 
                           => n4, C1 => comp_out(11), C2 => n5, ZN => n11);
   U20 : INV_X1 port map( A => n12, ZN => outputSel(10));
   U21 : AOI222_X1 port map( A1 => p4_out(10), A2 => n1, B1 => LS_OUT(10), B2 
                           => n4, C1 => comp_out(10), C2 => n5, ZN => n12);
   U22 : INV_X1 port map( A => n13, ZN => outputSel(8));
   U23 : AOI222_X1 port map( A1 => p4_out(8), A2 => n1, B1 => LS_OUT(8), B2 => 
                           n4, C1 => comp_out(8), C2 => n5, ZN => n13);
   U24 : INV_X1 port map( A => n14, ZN => outputSel(13));
   U25 : AOI222_X1 port map( A1 => p4_out(13), A2 => n1, B1 => LS_OUT(13), B2 
                           => n4, C1 => comp_out(13), C2 => n5, ZN => n14);
   U26 : INV_X1 port map( A => n15, ZN => outputSel(15));
   U27 : AOI222_X1 port map( A1 => p4_out(15), A2 => n1, B1 => LS_OUT(15), B2 
                           => n4, C1 => comp_out(15), C2 => n5, ZN => n15);
   U28 : INV_X1 port map( A => n16, ZN => outputSel(14));
   U29 : AOI222_X1 port map( A1 => p4_out(14), A2 => n1, B1 => LS_OUT(14), B2 
                           => n4, C1 => comp_out(14), C2 => n5, ZN => n16);
   U30 : INV_X1 port map( A => n17, ZN => outputSel(12));
   U31 : AOI222_X1 port map( A1 => p4_out(12), A2 => n1, B1 => LS_OUT(12), B2 
                           => n4, C1 => comp_out(12), C2 => n5, ZN => n17);
   U32 : INV_X1 port map( A => n18, ZN => outputSel(17));
   U33 : AOI222_X1 port map( A1 => p4_out(17), A2 => n1, B1 => LS_OUT(17), B2 
                           => n4, C1 => comp_out(17), C2 => n5, ZN => n18);
   U34 : INV_X1 port map( A => n19, ZN => outputSel(19));
   U35 : AOI222_X1 port map( A1 => p4_out(19), A2 => n1, B1 => LS_OUT(19), B2 
                           => n4, C1 => comp_out(19), C2 => n5, ZN => n19);
   U36 : INV_X1 port map( A => n20, ZN => outputSel(18));
   U37 : AOI222_X1 port map( A1 => p4_out(18), A2 => n1, B1 => LS_OUT(18), B2 
                           => n4, C1 => comp_out(18), C2 => n5, ZN => n20);
   U38 : INV_X1 port map( A => n21, ZN => outputSel(16));
   U39 : AOI222_X1 port map( A1 => p4_out(16), A2 => n1, B1 => LS_OUT(16), B2 
                           => n4, C1 => comp_out(16), C2 => n5, ZN => n21);
   U40 : INV_X1 port map( A => n22, ZN => outputSel(21));
   U41 : AOI222_X1 port map( A1 => p4_out(21), A2 => n1, B1 => LS_OUT(21), B2 
                           => n4, C1 => comp_out(21), C2 => n5, ZN => n22);
   U42 : INV_X1 port map( A => n23, ZN => outputSel(23));
   U43 : AOI222_X1 port map( A1 => p4_out(23), A2 => n1, B1 => LS_OUT(23), B2 
                           => n4, C1 => comp_out(23), C2 => n5, ZN => n23);
   U44 : INV_X1 port map( A => n24, ZN => outputSel(22));
   U45 : AOI222_X1 port map( A1 => p4_out(22), A2 => n1, B1 => LS_OUT(22), B2 
                           => n4, C1 => comp_out(22), C2 => n5, ZN => n24);
   U46 : INV_X1 port map( A => n25, ZN => outputSel(20));
   U47 : AOI222_X1 port map( A1 => p4_out(20), A2 => n1, B1 => LS_OUT(20), B2 
                           => n4, C1 => comp_out(20), C2 => n5, ZN => n25);
   U48 : INV_X1 port map( A => n26, ZN => outputSel(25));
   U49 : AOI222_X1 port map( A1 => p4_out(25), A2 => n1, B1 => LS_OUT(25), B2 
                           => n4, C1 => comp_out(25), C2 => n5, ZN => n26);
   U50 : INV_X1 port map( A => n27, ZN => outputSel(27));
   U51 : AOI222_X1 port map( A1 => p4_out(27), A2 => n1, B1 => LS_OUT(27), B2 
                           => n4, C1 => comp_out(27), C2 => n5, ZN => n27);
   U52 : INV_X1 port map( A => n28, ZN => outputSel(26));
   U53 : AOI222_X1 port map( A1 => p4_out(26), A2 => n1, B1 => LS_OUT(26), B2 
                           => n4, C1 => comp_out(26), C2 => n5, ZN => n28);
   U54 : INV_X1 port map( A => n29, ZN => outputSel(24));
   U55 : AOI222_X1 port map( A1 => p4_out(24), A2 => n1, B1 => LS_OUT(24), B2 
                           => n4, C1 => comp_out(24), C2 => n5, ZN => n29);
   U56 : INV_X1 port map( A => n30, ZN => outputSel(29));
   U57 : AOI222_X1 port map( A1 => p4_out(29), A2 => n1, B1 => LS_OUT(29), B2 
                           => n4, C1 => comp_out(29), C2 => n5, ZN => n30);
   U58 : INV_X1 port map( A => n31, ZN => outputSel(31));
   U59 : AOI222_X1 port map( A1 => p4_out(31), A2 => n1, B1 => LS_OUT(31), B2 
                           => n4, C1 => comp_out(31), C2 => n5, ZN => n31);
   U60 : INV_X1 port map( A => n32, ZN => outputSel(30));
   U61 : AOI222_X1 port map( A1 => p4_out(30), A2 => n1, B1 => LS_OUT(30), B2 
                           => n4, C1 => comp_out(30), C2 => n5, ZN => n32);
   U62 : INV_X1 port map( A => n33, ZN => outputSel(28));
   U63 : AOI222_X1 port map( A1 => p4_out(28), A2 => n1, B1 => LS_OUT(28), B2 
                           => n4, C1 => comp_out(28), C2 => n5, ZN => n33);
   U64 : INV_X1 port map( A => n34, ZN => outputSel(3));
   U65 : AOI222_X1 port map( A1 => p4_out(3), A2 => n1, B1 => LS_OUT(3), B2 => 
                           n4, C1 => comp_out(3), C2 => n5, ZN => n34);
   U66 : INV_X1 port map( A => n35, ZN => outputSel(2));
   U67 : AOI222_X1 port map( A1 => p4_out(2), A2 => n1, B1 => LS_OUT(2), B2 => 
                           n4, C1 => comp_out(2), C2 => n5, ZN => n35);
   U68 : INV_X1 port map( A => n36, ZN => outputSel(1));
   U69 : AOI222_X1 port map( A1 => p4_out(1), A2 => n1, B1 => LS_OUT(1), B2 => 
                           n4, C1 => comp_out(1), C2 => n5, ZN => n36);
   U70 : MUX2_X1 port map( A => n38, B => n39, S => n40, Z => n37);
   U71 : NAND2_X1 port map( A1 => FUNC(0), A2 => n41, ZN => n39);
   U72 : NAND3_X1 port map( A1 => FUNC(2), A2 => n42, A3 => FUNC(3), ZN => n38)
                           ;
   U73 : INV_X1 port map( A => FUNC(0), ZN => n42);
   U74 : OAI21_X1 port map( B1 => FUNC(3), B2 => n40, A => FUNC(2), ZN => n43);
   U75 : INV_X1 port map( A => FUNC(1), ZN => n40);
   U76 : INV_X1 port map( A => FUNC(2), ZN => n41);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21;

architecture SYN_BEHAVIORAL of MUX21 is

   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X2 port map( A => B, B => A, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_0 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_0;

architecture SYN_ASYNCH_FD of FD_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n3, n4, n_1372 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CK, RN => n3, Q => Q_port, QN => 
                           n_1372);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n4);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n3);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity XNOR_logic is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR_logic;

architecture SYN_BEHAVIORAL of XNOR_logic is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity alu_nbits32 is

   port( FUNC : in std_logic_vector (0 to 3);  A, B : in std_logic_vector (31 
         downto 0);  OUTALU : out std_logic_vector (31 downto 0));

end alu_nbits32;

architecture SYN_STRUCTURAL of alu_nbits32 is

   component logic_and_shift_N32
      port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4_ADDER_NBITS32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component ctrl_alu_NBITS32
      port( A, B : in std_logic_vector (31 downto 0);  FUNC : in 
            std_logic_vector (0 to 3);  Ap4, Bp4 : out std_logic_vector (31 
            downto 0);  Cin : out std_logic;  Als, Bls : out std_logic_vector 
            (31 downto 0);  enableComp : out std_logic);
   end component;
   
   component comparator_bits32
      port( Cout, EN : in std_logic;  func : in std_logic_vector (0 to 3);  sum
            : in std_logic_vector (31 downto 0);  set : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component outputSelect_nbits32
      port( FUNC : in std_logic_vector (0 to 3);  p4_out, LS_OUT, comp_out : in
            std_logic_vector (31 downto 0);  outputSel : out std_logic_vector 
            (31 downto 0));
   end component;
   
   signal p4_outsig_31_port, p4_outsig_30_port, p4_outsig_29_port, 
      p4_outsig_28_port, p4_outsig_27_port, p4_outsig_26_port, 
      p4_outsig_25_port, p4_outsig_24_port, p4_outsig_23_port, 
      p4_outsig_22_port, p4_outsig_21_port, p4_outsig_20_port, 
      p4_outsig_19_port, p4_outsig_18_port, p4_outsig_17_port, 
      p4_outsig_16_port, p4_outsig_15_port, p4_outsig_14_port, 
      p4_outsig_13_port, p4_outsig_12_port, p4_outsig_11_port, 
      p4_outsig_10_port, p4_outsig_9_port, p4_outsig_8_port, p4_outsig_7_port, 
      p4_outsig_6_port, p4_outsig_5_port, p4_outsig_4_port, p4_outsig_3_port, 
      p4_outsig_2_port, p4_outsig_1_port, p4_outsig_0_port, LS_OUTsig_31_port, 
      LS_OUTsig_30_port, LS_OUTsig_29_port, LS_OUTsig_28_port, 
      LS_OUTsig_27_port, LS_OUTsig_26_port, LS_OUTsig_25_port, 
      LS_OUTsig_24_port, LS_OUTsig_23_port, LS_OUTsig_22_port, 
      LS_OUTsig_21_port, LS_OUTsig_20_port, LS_OUTsig_19_port, 
      LS_OUTsig_18_port, LS_OUTsig_17_port, LS_OUTsig_16_port, 
      LS_OUTsig_15_port, LS_OUTsig_14_port, LS_OUTsig_13_port, 
      LS_OUTsig_12_port, LS_OUTsig_11_port, LS_OUTsig_10_port, LS_OUTsig_9_port
      , LS_OUTsig_8_port, LS_OUTsig_7_port, LS_OUTsig_6_port, LS_OUTsig_5_port,
      LS_OUTsig_4_port, LS_OUTsig_3_port, LS_OUTsig_2_port, LS_OUTsig_1_port, 
      LS_OUTsig_0_port, comp_outsig_31_port, comp_outsig_30_port, 
      comp_outsig_29_port, comp_outsig_28_port, comp_outsig_27_port, 
      comp_outsig_26_port, comp_outsig_25_port, comp_outsig_24_port, 
      comp_outsig_23_port, comp_outsig_22_port, comp_outsig_21_port, 
      comp_outsig_20_port, comp_outsig_19_port, comp_outsig_18_port, 
      comp_outsig_17_port, comp_outsig_16_port, comp_outsig_15_port, 
      comp_outsig_14_port, comp_outsig_13_port, comp_outsig_12_port, 
      comp_outsig_11_port, comp_outsig_10_port, comp_outsig_9_port, 
      comp_outsig_8_port, comp_outsig_7_port, comp_outsig_6_port, 
      comp_outsig_5_port, comp_outsig_4_port, comp_outsig_3_port, 
      comp_outsig_2_port, comp_outsig_1_port, comp_outsig_0_port, p4_comp_Co, 
      enable_Comp, p4_ctrl_A_31_port, p4_ctrl_A_30_port, p4_ctrl_A_29_port, 
      p4_ctrl_A_28_port, p4_ctrl_A_27_port, p4_ctrl_A_26_port, 
      p4_ctrl_A_25_port, p4_ctrl_A_24_port, p4_ctrl_A_23_port, 
      p4_ctrl_A_22_port, p4_ctrl_A_21_port, p4_ctrl_A_20_port, 
      p4_ctrl_A_19_port, p4_ctrl_A_18_port, p4_ctrl_A_17_port, 
      p4_ctrl_A_16_port, p4_ctrl_A_15_port, p4_ctrl_A_14_port, 
      p4_ctrl_A_13_port, p4_ctrl_A_12_port, p4_ctrl_A_11_port, 
      p4_ctrl_A_10_port, p4_ctrl_A_9_port, p4_ctrl_A_8_port, p4_ctrl_A_7_port, 
      p4_ctrl_A_6_port, p4_ctrl_A_5_port, p4_ctrl_A_4_port, p4_ctrl_A_3_port, 
      p4_ctrl_A_2_port, p4_ctrl_A_1_port, p4_ctrl_A_0_port, p4_ctrl_B_31_port, 
      p4_ctrl_B_30_port, p4_ctrl_B_29_port, p4_ctrl_B_28_port, 
      p4_ctrl_B_27_port, p4_ctrl_B_26_port, p4_ctrl_B_25_port, 
      p4_ctrl_B_24_port, p4_ctrl_B_23_port, p4_ctrl_B_22_port, 
      p4_ctrl_B_21_port, p4_ctrl_B_20_port, p4_ctrl_B_19_port, 
      p4_ctrl_B_18_port, p4_ctrl_B_17_port, p4_ctrl_B_16_port, 
      p4_ctrl_B_15_port, p4_ctrl_B_14_port, p4_ctrl_B_13_port, 
      p4_ctrl_B_12_port, p4_ctrl_B_11_port, p4_ctrl_B_10_port, p4_ctrl_B_9_port
      , p4_ctrl_B_8_port, p4_ctrl_B_7_port, p4_ctrl_B_6_port, p4_ctrl_B_5_port,
      p4_ctrl_B_4_port, p4_ctrl_B_3_port, p4_ctrl_B_2_port, p4_ctrl_B_1_port, 
      p4_ctrl_B_0_port, p4_ctrl_Cin, ctrl_LS_A_31_port, ctrl_LS_A_30_port, 
      ctrl_LS_A_29_port, ctrl_LS_A_28_port, ctrl_LS_A_27_port, 
      ctrl_LS_A_26_port, ctrl_LS_A_25_port, ctrl_LS_A_24_port, 
      ctrl_LS_A_23_port, ctrl_LS_A_22_port, ctrl_LS_A_21_port, 
      ctrl_LS_A_20_port, ctrl_LS_A_19_port, ctrl_LS_A_18_port, 
      ctrl_LS_A_17_port, ctrl_LS_A_16_port, ctrl_LS_A_15_port, 
      ctrl_LS_A_14_port, ctrl_LS_A_13_port, ctrl_LS_A_12_port, 
      ctrl_LS_A_11_port, ctrl_LS_A_10_port, ctrl_LS_A_9_port, ctrl_LS_A_8_port,
      ctrl_LS_A_7_port, ctrl_LS_A_6_port, ctrl_LS_A_5_port, ctrl_LS_A_4_port, 
      ctrl_LS_A_3_port, ctrl_LS_A_2_port, ctrl_LS_A_1_port, ctrl_LS_A_0_port, 
      ctrl_LS_B_31_port, ctrl_LS_B_30_port, ctrl_LS_B_29_port, 
      ctrl_LS_B_28_port, ctrl_LS_B_27_port, ctrl_LS_B_26_port, 
      ctrl_LS_B_25_port, ctrl_LS_B_24_port, ctrl_LS_B_23_port, 
      ctrl_LS_B_22_port, ctrl_LS_B_21_port, ctrl_LS_B_20_port, 
      ctrl_LS_B_19_port, ctrl_LS_B_18_port, ctrl_LS_B_17_port, 
      ctrl_LS_B_16_port, ctrl_LS_B_15_port, ctrl_LS_B_14_port, 
      ctrl_LS_B_13_port, ctrl_LS_B_12_port, ctrl_LS_B_11_port, 
      ctrl_LS_B_10_port, ctrl_LS_B_9_port, ctrl_LS_B_8_port, ctrl_LS_B_7_port, 
      ctrl_LS_B_6_port, ctrl_LS_B_5_port, ctrl_LS_B_4_port, ctrl_LS_B_3_port, 
      ctrl_LS_B_2_port, ctrl_LS_B_1_port, ctrl_LS_B_0_port, n_1373, n_1374, 
      n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, 
      n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, 
      n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, 
      n_1402, n_1403 : std_logic;

begin
   
   SELOUT : outputSelect_nbits32 port map( FUNC(0) => FUNC(0), FUNC(1) => 
                           FUNC(1), FUNC(2) => FUNC(2), FUNC(3) => FUNC(3), 
                           p4_out(31) => p4_outsig_31_port, p4_out(30) => 
                           p4_outsig_30_port, p4_out(29) => p4_outsig_29_port, 
                           p4_out(28) => p4_outsig_28_port, p4_out(27) => 
                           p4_outsig_27_port, p4_out(26) => p4_outsig_26_port, 
                           p4_out(25) => p4_outsig_25_port, p4_out(24) => 
                           p4_outsig_24_port, p4_out(23) => p4_outsig_23_port, 
                           p4_out(22) => p4_outsig_22_port, p4_out(21) => 
                           p4_outsig_21_port, p4_out(20) => p4_outsig_20_port, 
                           p4_out(19) => p4_outsig_19_port, p4_out(18) => 
                           p4_outsig_18_port, p4_out(17) => p4_outsig_17_port, 
                           p4_out(16) => p4_outsig_16_port, p4_out(15) => 
                           p4_outsig_15_port, p4_out(14) => p4_outsig_14_port, 
                           p4_out(13) => p4_outsig_13_port, p4_out(12) => 
                           p4_outsig_12_port, p4_out(11) => p4_outsig_11_port, 
                           p4_out(10) => p4_outsig_10_port, p4_out(9) => 
                           p4_outsig_9_port, p4_out(8) => p4_outsig_8_port, 
                           p4_out(7) => p4_outsig_7_port, p4_out(6) => 
                           p4_outsig_6_port, p4_out(5) => p4_outsig_5_port, 
                           p4_out(4) => p4_outsig_4_port, p4_out(3) => 
                           p4_outsig_3_port, p4_out(2) => p4_outsig_2_port, 
                           p4_out(1) => p4_outsig_1_port, p4_out(0) => 
                           p4_outsig_0_port, LS_OUT(31) => LS_OUTsig_31_port, 
                           LS_OUT(30) => LS_OUTsig_30_port, LS_OUT(29) => 
                           LS_OUTsig_29_port, LS_OUT(28) => LS_OUTsig_28_port, 
                           LS_OUT(27) => LS_OUTsig_27_port, LS_OUT(26) => 
                           LS_OUTsig_26_port, LS_OUT(25) => LS_OUTsig_25_port, 
                           LS_OUT(24) => LS_OUTsig_24_port, LS_OUT(23) => 
                           LS_OUTsig_23_port, LS_OUT(22) => LS_OUTsig_22_port, 
                           LS_OUT(21) => LS_OUTsig_21_port, LS_OUT(20) => 
                           LS_OUTsig_20_port, LS_OUT(19) => LS_OUTsig_19_port, 
                           LS_OUT(18) => LS_OUTsig_18_port, LS_OUT(17) => 
                           LS_OUTsig_17_port, LS_OUT(16) => LS_OUTsig_16_port, 
                           LS_OUT(15) => LS_OUTsig_15_port, LS_OUT(14) => 
                           LS_OUTsig_14_port, LS_OUT(13) => LS_OUTsig_13_port, 
                           LS_OUT(12) => LS_OUTsig_12_port, LS_OUT(11) => 
                           LS_OUTsig_11_port, LS_OUT(10) => LS_OUTsig_10_port, 
                           LS_OUT(9) => LS_OUTsig_9_port, LS_OUT(8) => 
                           LS_OUTsig_8_port, LS_OUT(7) => LS_OUTsig_7_port, 
                           LS_OUT(6) => LS_OUTsig_6_port, LS_OUT(5) => 
                           LS_OUTsig_5_port, LS_OUT(4) => LS_OUTsig_4_port, 
                           LS_OUT(3) => LS_OUTsig_3_port, LS_OUT(2) => 
                           LS_OUTsig_2_port, LS_OUT(1) => LS_OUTsig_1_port, 
                           LS_OUT(0) => LS_OUTsig_0_port, comp_out(31) => 
                           comp_outsig_31_port, comp_out(30) => 
                           comp_outsig_30_port, comp_out(29) => 
                           comp_outsig_29_port, comp_out(28) => 
                           comp_outsig_28_port, comp_out(27) => 
                           comp_outsig_27_port, comp_out(26) => 
                           comp_outsig_26_port, comp_out(25) => 
                           comp_outsig_25_port, comp_out(24) => 
                           comp_outsig_24_port, comp_out(23) => 
                           comp_outsig_23_port, comp_out(22) => 
                           comp_outsig_22_port, comp_out(21) => 
                           comp_outsig_21_port, comp_out(20) => 
                           comp_outsig_20_port, comp_out(19) => 
                           comp_outsig_19_port, comp_out(18) => 
                           comp_outsig_18_port, comp_out(17) => 
                           comp_outsig_17_port, comp_out(16) => 
                           comp_outsig_16_port, comp_out(15) => 
                           comp_outsig_15_port, comp_out(14) => 
                           comp_outsig_14_port, comp_out(13) => 
                           comp_outsig_13_port, comp_out(12) => 
                           comp_outsig_12_port, comp_out(11) => 
                           comp_outsig_11_port, comp_out(10) => 
                           comp_outsig_10_port, comp_out(9) => 
                           comp_outsig_9_port, comp_out(8) => 
                           comp_outsig_8_port, comp_out(7) => 
                           comp_outsig_7_port, comp_out(6) => 
                           comp_outsig_6_port, comp_out(5) => 
                           comp_outsig_5_port, comp_out(4) => 
                           comp_outsig_4_port, comp_out(3) => 
                           comp_outsig_3_port, comp_out(2) => 
                           comp_outsig_2_port, comp_out(1) => 
                           comp_outsig_1_port, comp_out(0) => 
                           comp_outsig_0_port, outputSel(31) => OUTALU(31), 
                           outputSel(30) => OUTALU(30), outputSel(29) => 
                           OUTALU(29), outputSel(28) => OUTALU(28), 
                           outputSel(27) => OUTALU(27), outputSel(26) => 
                           OUTALU(26), outputSel(25) => OUTALU(25), 
                           outputSel(24) => OUTALU(24), outputSel(23) => 
                           OUTALU(23), outputSel(22) => OUTALU(22), 
                           outputSel(21) => OUTALU(21), outputSel(20) => 
                           OUTALU(20), outputSel(19) => OUTALU(19), 
                           outputSel(18) => OUTALU(18), outputSel(17) => 
                           OUTALU(17), outputSel(16) => OUTALU(16), 
                           outputSel(15) => OUTALU(15), outputSel(14) => 
                           OUTALU(14), outputSel(13) => OUTALU(13), 
                           outputSel(12) => OUTALU(12), outputSel(11) => 
                           OUTALU(11), outputSel(10) => OUTALU(10), 
                           outputSel(9) => OUTALU(9), outputSel(8) => OUTALU(8)
                           , outputSel(7) => OUTALU(7), outputSel(6) => 
                           OUTALU(6), outputSel(5) => OUTALU(5), outputSel(4) 
                           => OUTALU(4), outputSel(3) => OUTALU(3), 
                           outputSel(2) => OUTALU(2), outputSel(1) => OUTALU(1)
                           , outputSel(0) => OUTALU(0));
   COMP : comparator_bits32 port map( Cout => p4_comp_Co, EN => enable_Comp, 
                           func(0) => FUNC(0), func(1) => FUNC(1), func(2) => 
                           FUNC(2), func(3) => FUNC(3), sum(31) => 
                           p4_outsig_31_port, sum(30) => p4_outsig_30_port, 
                           sum(29) => p4_outsig_29_port, sum(28) => 
                           p4_outsig_28_port, sum(27) => p4_outsig_27_port, 
                           sum(26) => p4_outsig_26_port, sum(25) => 
                           p4_outsig_25_port, sum(24) => p4_outsig_24_port, 
                           sum(23) => p4_outsig_23_port, sum(22) => 
                           p4_outsig_22_port, sum(21) => p4_outsig_21_port, 
                           sum(20) => p4_outsig_20_port, sum(19) => 
                           p4_outsig_19_port, sum(18) => p4_outsig_18_port, 
                           sum(17) => p4_outsig_17_port, sum(16) => 
                           p4_outsig_16_port, sum(15) => p4_outsig_15_port, 
                           sum(14) => p4_outsig_14_port, sum(13) => 
                           p4_outsig_13_port, sum(12) => p4_outsig_12_port, 
                           sum(11) => p4_outsig_11_port, sum(10) => 
                           p4_outsig_10_port, sum(9) => p4_outsig_9_port, 
                           sum(8) => p4_outsig_8_port, sum(7) => 
                           p4_outsig_7_port, sum(6) => p4_outsig_6_port, sum(5)
                           => p4_outsig_5_port, sum(4) => p4_outsig_4_port, 
                           sum(3) => p4_outsig_3_port, sum(2) => 
                           p4_outsig_2_port, sum(1) => p4_outsig_1_port, sum(0)
                           => p4_outsig_0_port, set(31) => n_1373, set(30) => 
                           n_1374, set(29) => n_1375, set(28) => n_1376, 
                           set(27) => n_1377, set(26) => n_1378, set(25) => 
                           n_1379, set(24) => n_1380, set(23) => n_1381, 
                           set(22) => n_1382, set(21) => n_1383, set(20) => 
                           n_1384, set(19) => n_1385, set(18) => n_1386, 
                           set(17) => n_1387, set(16) => n_1388, set(15) => 
                           n_1389, set(14) => n_1390, set(13) => n_1391, 
                           set(12) => n_1392, set(11) => n_1393, set(10) => 
                           n_1394, set(9) => n_1395, set(8) => n_1396, set(7) 
                           => n_1397, set(6) => n_1398, set(5) => n_1399, 
                           set(4) => n_1400, set(3) => n_1401, set(2) => n_1402
                           , set(1) => n_1403, set(0) => comp_outsig_0_port);
   CTRLALU : ctrl_alu_NBITS32 port map( A(31) => A(31), A(30) => A(30), A(29) 
                           => A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), FUNC(0) => FUNC(0), FUNC(1) => FUNC(1), 
                           FUNC(2) => FUNC(2), FUNC(3) => FUNC(3), Ap4(31) => 
                           p4_ctrl_A_31_port, Ap4(30) => p4_ctrl_A_30_port, 
                           Ap4(29) => p4_ctrl_A_29_port, Ap4(28) => 
                           p4_ctrl_A_28_port, Ap4(27) => p4_ctrl_A_27_port, 
                           Ap4(26) => p4_ctrl_A_26_port, Ap4(25) => 
                           p4_ctrl_A_25_port, Ap4(24) => p4_ctrl_A_24_port, 
                           Ap4(23) => p4_ctrl_A_23_port, Ap4(22) => 
                           p4_ctrl_A_22_port, Ap4(21) => p4_ctrl_A_21_port, 
                           Ap4(20) => p4_ctrl_A_20_port, Ap4(19) => 
                           p4_ctrl_A_19_port, Ap4(18) => p4_ctrl_A_18_port, 
                           Ap4(17) => p4_ctrl_A_17_port, Ap4(16) => 
                           p4_ctrl_A_16_port, Ap4(15) => p4_ctrl_A_15_port, 
                           Ap4(14) => p4_ctrl_A_14_port, Ap4(13) => 
                           p4_ctrl_A_13_port, Ap4(12) => p4_ctrl_A_12_port, 
                           Ap4(11) => p4_ctrl_A_11_port, Ap4(10) => 
                           p4_ctrl_A_10_port, Ap4(9) => p4_ctrl_A_9_port, 
                           Ap4(8) => p4_ctrl_A_8_port, Ap4(7) => 
                           p4_ctrl_A_7_port, Ap4(6) => p4_ctrl_A_6_port, Ap4(5)
                           => p4_ctrl_A_5_port, Ap4(4) => p4_ctrl_A_4_port, 
                           Ap4(3) => p4_ctrl_A_3_port, Ap4(2) => 
                           p4_ctrl_A_2_port, Ap4(1) => p4_ctrl_A_1_port, Ap4(0)
                           => p4_ctrl_A_0_port, Bp4(31) => p4_ctrl_B_31_port, 
                           Bp4(30) => p4_ctrl_B_30_port, Bp4(29) => 
                           p4_ctrl_B_29_port, Bp4(28) => p4_ctrl_B_28_port, 
                           Bp4(27) => p4_ctrl_B_27_port, Bp4(26) => 
                           p4_ctrl_B_26_port, Bp4(25) => p4_ctrl_B_25_port, 
                           Bp4(24) => p4_ctrl_B_24_port, Bp4(23) => 
                           p4_ctrl_B_23_port, Bp4(22) => p4_ctrl_B_22_port, 
                           Bp4(21) => p4_ctrl_B_21_port, Bp4(20) => 
                           p4_ctrl_B_20_port, Bp4(19) => p4_ctrl_B_19_port, 
                           Bp4(18) => p4_ctrl_B_18_port, Bp4(17) => 
                           p4_ctrl_B_17_port, Bp4(16) => p4_ctrl_B_16_port, 
                           Bp4(15) => p4_ctrl_B_15_port, Bp4(14) => 
                           p4_ctrl_B_14_port, Bp4(13) => p4_ctrl_B_13_port, 
                           Bp4(12) => p4_ctrl_B_12_port, Bp4(11) => 
                           p4_ctrl_B_11_port, Bp4(10) => p4_ctrl_B_10_port, 
                           Bp4(9) => p4_ctrl_B_9_port, Bp4(8) => 
                           p4_ctrl_B_8_port, Bp4(7) => p4_ctrl_B_7_port, Bp4(6)
                           => p4_ctrl_B_6_port, Bp4(5) => p4_ctrl_B_5_port, 
                           Bp4(4) => p4_ctrl_B_4_port, Bp4(3) => 
                           p4_ctrl_B_3_port, Bp4(2) => p4_ctrl_B_2_port, Bp4(1)
                           => p4_ctrl_B_1_port, Bp4(0) => p4_ctrl_B_0_port, Cin
                           => p4_ctrl_Cin, Als(31) => ctrl_LS_A_31_port, 
                           Als(30) => ctrl_LS_A_30_port, Als(29) => 
                           ctrl_LS_A_29_port, Als(28) => ctrl_LS_A_28_port, 
                           Als(27) => ctrl_LS_A_27_port, Als(26) => 
                           ctrl_LS_A_26_port, Als(25) => ctrl_LS_A_25_port, 
                           Als(24) => ctrl_LS_A_24_port, Als(23) => 
                           ctrl_LS_A_23_port, Als(22) => ctrl_LS_A_22_port, 
                           Als(21) => ctrl_LS_A_21_port, Als(20) => 
                           ctrl_LS_A_20_port, Als(19) => ctrl_LS_A_19_port, 
                           Als(18) => ctrl_LS_A_18_port, Als(17) => 
                           ctrl_LS_A_17_port, Als(16) => ctrl_LS_A_16_port, 
                           Als(15) => ctrl_LS_A_15_port, Als(14) => 
                           ctrl_LS_A_14_port, Als(13) => ctrl_LS_A_13_port, 
                           Als(12) => ctrl_LS_A_12_port, Als(11) => 
                           ctrl_LS_A_11_port, Als(10) => ctrl_LS_A_10_port, 
                           Als(9) => ctrl_LS_A_9_port, Als(8) => 
                           ctrl_LS_A_8_port, Als(7) => ctrl_LS_A_7_port, Als(6)
                           => ctrl_LS_A_6_port, Als(5) => ctrl_LS_A_5_port, 
                           Als(4) => ctrl_LS_A_4_port, Als(3) => 
                           ctrl_LS_A_3_port, Als(2) => ctrl_LS_A_2_port, Als(1)
                           => ctrl_LS_A_1_port, Als(0) => ctrl_LS_A_0_port, 
                           Bls(31) => ctrl_LS_B_31_port, Bls(30) => 
                           ctrl_LS_B_30_port, Bls(29) => ctrl_LS_B_29_port, 
                           Bls(28) => ctrl_LS_B_28_port, Bls(27) => 
                           ctrl_LS_B_27_port, Bls(26) => ctrl_LS_B_26_port, 
                           Bls(25) => ctrl_LS_B_25_port, Bls(24) => 
                           ctrl_LS_B_24_port, Bls(23) => ctrl_LS_B_23_port, 
                           Bls(22) => ctrl_LS_B_22_port, Bls(21) => 
                           ctrl_LS_B_21_port, Bls(20) => ctrl_LS_B_20_port, 
                           Bls(19) => ctrl_LS_B_19_port, Bls(18) => 
                           ctrl_LS_B_18_port, Bls(17) => ctrl_LS_B_17_port, 
                           Bls(16) => ctrl_LS_B_16_port, Bls(15) => 
                           ctrl_LS_B_15_port, Bls(14) => ctrl_LS_B_14_port, 
                           Bls(13) => ctrl_LS_B_13_port, Bls(12) => 
                           ctrl_LS_B_12_port, Bls(11) => ctrl_LS_B_11_port, 
                           Bls(10) => ctrl_LS_B_10_port, Bls(9) => 
                           ctrl_LS_B_9_port, Bls(8) => ctrl_LS_B_8_port, Bls(7)
                           => ctrl_LS_B_7_port, Bls(6) => ctrl_LS_B_6_port, 
                           Bls(5) => ctrl_LS_B_5_port, Bls(4) => 
                           ctrl_LS_B_4_port, Bls(3) => ctrl_LS_B_3_port, Bls(2)
                           => ctrl_LS_B_2_port, Bls(1) => ctrl_LS_B_1_port, 
                           Bls(0) => ctrl_LS_B_0_port, enableComp => 
                           enable_Comp);
   ADDER_SUB : P4_ADDER_NBITS32 port map( A(31) => p4_ctrl_A_31_port, A(30) => 
                           p4_ctrl_A_30_port, A(29) => p4_ctrl_A_29_port, A(28)
                           => p4_ctrl_A_28_port, A(27) => p4_ctrl_A_27_port, 
                           A(26) => p4_ctrl_A_26_port, A(25) => 
                           p4_ctrl_A_25_port, A(24) => p4_ctrl_A_24_port, A(23)
                           => p4_ctrl_A_23_port, A(22) => p4_ctrl_A_22_port, 
                           A(21) => p4_ctrl_A_21_port, A(20) => 
                           p4_ctrl_A_20_port, A(19) => p4_ctrl_A_19_port, A(18)
                           => p4_ctrl_A_18_port, A(17) => p4_ctrl_A_17_port, 
                           A(16) => p4_ctrl_A_16_port, A(15) => 
                           p4_ctrl_A_15_port, A(14) => p4_ctrl_A_14_port, A(13)
                           => p4_ctrl_A_13_port, A(12) => p4_ctrl_A_12_port, 
                           A(11) => p4_ctrl_A_11_port, A(10) => 
                           p4_ctrl_A_10_port, A(9) => p4_ctrl_A_9_port, A(8) =>
                           p4_ctrl_A_8_port, A(7) => p4_ctrl_A_7_port, A(6) => 
                           p4_ctrl_A_6_port, A(5) => p4_ctrl_A_5_port, A(4) => 
                           p4_ctrl_A_4_port, A(3) => p4_ctrl_A_3_port, A(2) => 
                           p4_ctrl_A_2_port, A(1) => p4_ctrl_A_1_port, A(0) => 
                           p4_ctrl_A_0_port, B(31) => p4_ctrl_B_31_port, B(30) 
                           => p4_ctrl_B_30_port, B(29) => p4_ctrl_B_29_port, 
                           B(28) => p4_ctrl_B_28_port, B(27) => 
                           p4_ctrl_B_27_port, B(26) => p4_ctrl_B_26_port, B(25)
                           => p4_ctrl_B_25_port, B(24) => p4_ctrl_B_24_port, 
                           B(23) => p4_ctrl_B_23_port, B(22) => 
                           p4_ctrl_B_22_port, B(21) => p4_ctrl_B_21_port, B(20)
                           => p4_ctrl_B_20_port, B(19) => p4_ctrl_B_19_port, 
                           B(18) => p4_ctrl_B_18_port, B(17) => 
                           p4_ctrl_B_17_port, B(16) => p4_ctrl_B_16_port, B(15)
                           => p4_ctrl_B_15_port, B(14) => p4_ctrl_B_14_port, 
                           B(13) => p4_ctrl_B_13_port, B(12) => 
                           p4_ctrl_B_12_port, B(11) => p4_ctrl_B_11_port, B(10)
                           => p4_ctrl_B_10_port, B(9) => p4_ctrl_B_9_port, B(8)
                           => p4_ctrl_B_8_port, B(7) => p4_ctrl_B_7_port, B(6) 
                           => p4_ctrl_B_6_port, B(5) => p4_ctrl_B_5_port, B(4) 
                           => p4_ctrl_B_4_port, B(3) => p4_ctrl_B_3_port, B(2) 
                           => p4_ctrl_B_2_port, B(1) => p4_ctrl_B_1_port, B(0) 
                           => p4_ctrl_B_0_port, Ci => p4_ctrl_Cin, S(31) => 
                           p4_outsig_31_port, S(30) => p4_outsig_30_port, S(29)
                           => p4_outsig_29_port, S(28) => p4_outsig_28_port, 
                           S(27) => p4_outsig_27_port, S(26) => 
                           p4_outsig_26_port, S(25) => p4_outsig_25_port, S(24)
                           => p4_outsig_24_port, S(23) => p4_outsig_23_port, 
                           S(22) => p4_outsig_22_port, S(21) => 
                           p4_outsig_21_port, S(20) => p4_outsig_20_port, S(19)
                           => p4_outsig_19_port, S(18) => p4_outsig_18_port, 
                           S(17) => p4_outsig_17_port, S(16) => 
                           p4_outsig_16_port, S(15) => p4_outsig_15_port, S(14)
                           => p4_outsig_14_port, S(13) => p4_outsig_13_port, 
                           S(12) => p4_outsig_12_port, S(11) => 
                           p4_outsig_11_port, S(10) => p4_outsig_10_port, S(9) 
                           => p4_outsig_9_port, S(8) => p4_outsig_8_port, S(7) 
                           => p4_outsig_7_port, S(6) => p4_outsig_6_port, S(5) 
                           => p4_outsig_5_port, S(4) => p4_outsig_4_port, S(3) 
                           => p4_outsig_3_port, S(2) => p4_outsig_2_port, S(1) 
                           => p4_outsig_1_port, S(0) => p4_outsig_0_port, Co =>
                           p4_comp_Co);
   LOGIC_SHIFT : logic_and_shift_N32 port map( FUNC(0) => FUNC(0), FUNC(1) => 
                           FUNC(1), FUNC(2) => FUNC(2), FUNC(3) => FUNC(3), 
                           DATA1(31) => ctrl_LS_A_31_port, DATA1(30) => 
                           ctrl_LS_A_30_port, DATA1(29) => ctrl_LS_A_29_port, 
                           DATA1(28) => ctrl_LS_A_28_port, DATA1(27) => 
                           ctrl_LS_A_27_port, DATA1(26) => ctrl_LS_A_26_port, 
                           DATA1(25) => ctrl_LS_A_25_port, DATA1(24) => 
                           ctrl_LS_A_24_port, DATA1(23) => ctrl_LS_A_23_port, 
                           DATA1(22) => ctrl_LS_A_22_port, DATA1(21) => 
                           ctrl_LS_A_21_port, DATA1(20) => ctrl_LS_A_20_port, 
                           DATA1(19) => ctrl_LS_A_19_port, DATA1(18) => 
                           ctrl_LS_A_18_port, DATA1(17) => ctrl_LS_A_17_port, 
                           DATA1(16) => ctrl_LS_A_16_port, DATA1(15) => 
                           ctrl_LS_A_15_port, DATA1(14) => ctrl_LS_A_14_port, 
                           DATA1(13) => ctrl_LS_A_13_port, DATA1(12) => 
                           ctrl_LS_A_12_port, DATA1(11) => ctrl_LS_A_11_port, 
                           DATA1(10) => ctrl_LS_A_10_port, DATA1(9) => 
                           ctrl_LS_A_9_port, DATA1(8) => ctrl_LS_A_8_port, 
                           DATA1(7) => ctrl_LS_A_7_port, DATA1(6) => 
                           ctrl_LS_A_6_port, DATA1(5) => ctrl_LS_A_5_port, 
                           DATA1(4) => ctrl_LS_A_4_port, DATA1(3) => 
                           ctrl_LS_A_3_port, DATA1(2) => ctrl_LS_A_2_port, 
                           DATA1(1) => ctrl_LS_A_1_port, DATA1(0) => 
                           ctrl_LS_A_0_port, DATA2(31) => ctrl_LS_B_31_port, 
                           DATA2(30) => ctrl_LS_B_30_port, DATA2(29) => 
                           ctrl_LS_B_29_port, DATA2(28) => ctrl_LS_B_28_port, 
                           DATA2(27) => ctrl_LS_B_27_port, DATA2(26) => 
                           ctrl_LS_B_26_port, DATA2(25) => ctrl_LS_B_25_port, 
                           DATA2(24) => ctrl_LS_B_24_port, DATA2(23) => 
                           ctrl_LS_B_23_port, DATA2(22) => ctrl_LS_B_22_port, 
                           DATA2(21) => ctrl_LS_B_21_port, DATA2(20) => 
                           ctrl_LS_B_20_port, DATA2(19) => ctrl_LS_B_19_port, 
                           DATA2(18) => ctrl_LS_B_18_port, DATA2(17) => 
                           ctrl_LS_B_17_port, DATA2(16) => ctrl_LS_B_16_port, 
                           DATA2(15) => ctrl_LS_B_15_port, DATA2(14) => 
                           ctrl_LS_B_14_port, DATA2(13) => ctrl_LS_B_13_port, 
                           DATA2(12) => ctrl_LS_B_12_port, DATA2(11) => 
                           ctrl_LS_B_11_port, DATA2(10) => ctrl_LS_B_10_port, 
                           DATA2(9) => ctrl_LS_B_9_port, DATA2(8) => 
                           ctrl_LS_B_8_port, DATA2(7) => ctrl_LS_B_7_port, 
                           DATA2(6) => ctrl_LS_B_6_port, DATA2(5) => 
                           ctrl_LS_B_5_port, DATA2(4) => ctrl_LS_B_4_port, 
                           DATA2(3) => ctrl_LS_B_3_port, DATA2(2) => 
                           ctrl_LS_B_2_port, DATA2(1) => ctrl_LS_B_1_port, 
                           DATA2(0) => ctrl_LS_B_0_port, OUTALU(31) => 
                           LS_OUTsig_31_port, OUTALU(30) => LS_OUTsig_30_port, 
                           OUTALU(29) => LS_OUTsig_29_port, OUTALU(28) => 
                           LS_OUTsig_28_port, OUTALU(27) => LS_OUTsig_27_port, 
                           OUTALU(26) => LS_OUTsig_26_port, OUTALU(25) => 
                           LS_OUTsig_25_port, OUTALU(24) => LS_OUTsig_24_port, 
                           OUTALU(23) => LS_OUTsig_23_port, OUTALU(22) => 
                           LS_OUTsig_22_port, OUTALU(21) => LS_OUTsig_21_port, 
                           OUTALU(20) => LS_OUTsig_20_port, OUTALU(19) => 
                           LS_OUTsig_19_port, OUTALU(18) => LS_OUTsig_18_port, 
                           OUTALU(17) => LS_OUTsig_17_port, OUTALU(16) => 
                           LS_OUTsig_16_port, OUTALU(15) => LS_OUTsig_15_port, 
                           OUTALU(14) => LS_OUTsig_14_port, OUTALU(13) => 
                           LS_OUTsig_13_port, OUTALU(12) => LS_OUTsig_12_port, 
                           OUTALU(11) => LS_OUTsig_11_port, OUTALU(10) => 
                           LS_OUTsig_10_port, OUTALU(9) => LS_OUTsig_9_port, 
                           OUTALU(8) => LS_OUTsig_8_port, OUTALU(7) => 
                           LS_OUTsig_7_port, OUTALU(6) => LS_OUTsig_6_port, 
                           OUTALU(5) => LS_OUTsig_5_port, OUTALU(4) => 
                           LS_OUTsig_4_port, OUTALU(3) => LS_OUTsig_3_port, 
                           OUTALU(2) => LS_OUTsig_2_port, OUTALU(1) => 
                           LS_OUTsig_1_port, OUTALU(0) => LS_OUTsig_0_port);
   comp_outsig_1_port <= '0';
   comp_outsig_2_port <= '0';
   comp_outsig_3_port <= '0';
   comp_outsig_4_port <= '0';
   comp_outsig_5_port <= '0';
   comp_outsig_6_port <= '0';
   comp_outsig_7_port <= '0';
   comp_outsig_8_port <= '0';
   comp_outsig_9_port <= '0';
   comp_outsig_10_port <= '0';
   comp_outsig_11_port <= '0';
   comp_outsig_12_port <= '0';
   comp_outsig_13_port <= '0';
   comp_outsig_14_port <= '0';
   comp_outsig_15_port <= '0';
   comp_outsig_16_port <= '0';
   comp_outsig_17_port <= '0';
   comp_outsig_18_port <= '0';
   comp_outsig_19_port <= '0';
   comp_outsig_20_port <= '0';
   comp_outsig_21_port <= '0';
   comp_outsig_22_port <= '0';
   comp_outsig_23_port <= '0';
   comp_outsig_24_port <= '0';
   comp_outsig_25_port <= '0';
   comp_outsig_26_port <= '0';
   comp_outsig_27_port <= '0';
   comp_outsig_28_port <= '0';
   comp_outsig_29_port <= '0';
   comp_outsig_30_port <= '0';
   comp_outsig_31_port <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_0;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U5 : MUX2_X1 port map( A => B(4), B => A(4), S => S, Z => Y(4));
   U6 : MUX2_X1 port map( A => B(5), B => A(5), S => S, Z => Y(5));
   U7 : MUX2_X1 port map( A => B(6), B => A(6), S => S, Z => Y(6));
   U8 : MUX2_X1 port map( A => B(7), B => A(7), S => S, Z => Y(7));
   U9 : MUX2_X1 port map( A => B(8), B => A(8), S => S, Z => Y(8));
   U10 : MUX2_X1 port map( A => B(9), B => A(9), S => S, Z => Y(9));
   U11 : MUX2_X1 port map( A => B(10), B => A(10), S => S, Z => Y(10));
   U12 : MUX2_X1 port map( A => B(11), B => A(11), S => S, Z => Y(11));
   U13 : MUX2_X1 port map( A => B(12), B => A(12), S => S, Z => Y(12));
   U14 : MUX2_X1 port map( A => B(13), B => A(13), S => S, Z => Y(13));
   U15 : MUX2_X1 port map( A => B(14), B => A(14), S => S, Z => Y(14));
   U16 : MUX2_X1 port map( A => B(15), B => A(15), S => S, Z => Y(15));
   U17 : MUX2_X1 port map( A => B(16), B => A(16), S => S, Z => Y(16));
   U18 : MUX2_X1 port map( A => B(17), B => A(17), S => S, Z => Y(17));
   U19 : MUX2_X1 port map( A => B(18), B => A(18), S => S, Z => Y(18));
   U20 : MUX2_X1 port map( A => B(19), B => A(19), S => S, Z => Y(19));
   U21 : MUX2_X1 port map( A => B(20), B => A(20), S => S, Z => Y(20));
   U22 : MUX2_X1 port map( A => B(21), B => A(21), S => S, Z => Y(21));
   U23 : MUX2_X1 port map( A => B(22), B => A(22), S => S, Z => Y(22));
   U24 : MUX2_X1 port map( A => B(23), B => A(23), S => S, Z => Y(23));
   U25 : MUX2_X1 port map( A => B(24), B => A(24), S => S, Z => Y(24));
   U26 : MUX2_X1 port map( A => B(25), B => A(25), S => S, Z => Y(25));
   U27 : MUX2_X1 port map( A => B(26), B => A(26), S => S, Z => Y(26));
   U28 : MUX2_X1 port map( A => B(27), B => A(27), S => S, Z => Y(27));
   U29 : MUX2_X1 port map( A => B(28), B => A(28), S => S, Z => Y(28));
   U30 : MUX2_X1 port map( A => B(29), B => A(29), S => S, Z => Y(29));
   U31 : MUX2_X1 port map( A => B(30), B => A(30), S => S, Z => Y(30));
   U32 : MUX2_X1 port map( A => B(31), B => A(31), S => S, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ZERO_DEC_bits32 is

   port( data : in std_logic_vector (31 downto 0);  zero_detect : out std_logic
         );

end ZERO_DEC_bits32;

architecture SYN_BEHAVIORAL of ZERO_DEC_bits32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => zero_detect);
   U2 : NAND4_X1 port map( A1 => n3, A2 => n4, A3 => n5, A4 => n6, ZN => n2);
   U3 : NOR4_X1 port map( A1 => data(23), A2 => data(22), A3 => data(21), A4 =>
                           data(20), ZN => n6);
   U4 : NOR4_X1 port map( A1 => data(1), A2 => data(19), A3 => data(18), A4 => 
                           data(17), ZN => n5);
   U5 : NOR4_X1 port map( A1 => data(16), A2 => data(15), A3 => data(14), A4 =>
                           data(13), ZN => n4);
   U6 : NOR4_X1 port map( A1 => data(12), A2 => data(11), A3 => data(10), A4 =>
                           data(0), ZN => n3);
   U7 : NAND4_X1 port map( A1 => n7, A2 => n8, A3 => n9, A4 => n10, ZN => n1);
   U8 : NOR4_X1 port map( A1 => data(9), A2 => data(8), A3 => data(7), A4 => 
                           data(6), ZN => n10);
   U9 : NOR4_X1 port map( A1 => data(5), A2 => data(4), A3 => data(3), A4 => 
                           data(31), ZN => n9);
   U10 : NOR4_X1 port map( A1 => data(30), A2 => data(2), A3 => data(29), A4 =>
                           data(28), ZN => n8);
   U11 : NOR4_X1 port map( A1 => data(27), A2 => data(26), A3 => data(25), A4 
                           => data(24), ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity REGISTER_FILE_NBITS32_NREGISTERS32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end REGISTER_FILE_NBITS32_NREGISTERS32;

architecture SYN_BEHAVIORAL of REGISTER_FILE_NBITS32_NREGISTERS32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, 
      N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84
      , N85, N86, N87, N88, N89, N90, N91, N127, N128, N129, N130, N131, N132, 
      N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, 
      N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, 
      N157, N158, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311
      , n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, 
      n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, 
      n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, 
      n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, 
      n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, 
      n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, 
      n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, 
      n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, 
      n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
      n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, 
      n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
      n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
      n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, 
      n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, 
      n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, 
      n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, 
      n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, 
      n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, 
      n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, 
      n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, 
      n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
      n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, 
      n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, 
      n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, 
      n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, 
      n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, 
      n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, 
      n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, 
      n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, 
      n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, 
      n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, 
      n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, 
      n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, 
      n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, 
      n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, 
      n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, 
      n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, 
      n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, 
      n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, 
      n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, 
      n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, 
      n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, 
      n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, 
      n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, 
      n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, 
      n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, 
      n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, 
      n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, 
      n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, 
      n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, 
      n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, 
      n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, 
      n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, 
      n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, 
      n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, 
      n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, 
      n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, 
      n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, 
      n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, 
      n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, 
      n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, 
      n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, 
      n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, 
      n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, 
      n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, 
      n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, 
      n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, 
      n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, 
      n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, 
      n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, 
      n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, 
      n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, 
      n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, 
      n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, 
      n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, 
      n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, 
      n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, 
      n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, 
      n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, 
      n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, 
      n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, 
      n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, 
      n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, 
      n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, 
      n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, 
      n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, 
      n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, 
      n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, 
      n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, 
      n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, 
      n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, 
      n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, 
      n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, 
      n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, 
      n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, 
      n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, 
      n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, 
      n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, 
      n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, 
      n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, 
      n2322, n2323, n2324, n2325, n2326, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60_port, n61_port, n62_port, n63_port, 
      n64_port, n65_port, n66_port, n67_port, n68_port, n69_port, n70_port, 
      n71_port, n72_port, n73_port, n74_port, n75_port, n76_port, n77_port, 
      n78_port, n79_port, n80_port, n81_port, n82_port, n83_port, n84_port, 
      n85_port, n86_port, n87_port, n88_port, n89_port, n90_port, n91_port, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127_port, 
      n128_port, n129_port, n130_port, n131_port, n132_port, n133_port, 
      n134_port, n135_port, n136_port, n137_port, n138_port, n139_port, 
      n140_port, n141_port, n142_port, n143_port, n144_port, n145_port, 
      n146_port, n147_port, n148_port, n149_port, n150_port, n151_port, 
      n152_port, n153_port, n154_port, n155_port, n156_port, n157_port, 
      n158_port, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
      n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
      n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, 
      n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
      n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
      n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
      n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
      n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
      n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
      n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
      n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
      n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, 
      n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, 
      n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
      n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, 
      n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, 
      n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, 
      n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, 
      n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, 
      n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, 
      n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, 
      n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, 
      n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, 
      n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, 
      n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, 
      n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
      n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, 
      n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, 
      n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, 
      n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, 
      n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, 
      n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, 
      n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, 
      n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, 
      n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, 
      n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, 
      n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, 
      n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, 
      n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, 
      n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, 
      n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, 
      n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, 
      n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, 
      n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, 
      n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, 
      n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, 
      n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, 
      n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, 
      n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, 
      n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, 
      n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, 
      n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, 
      n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, 
      n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, 
      n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, 
      n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, 
      n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, 
      n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, 
      n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
      n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, 
      n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
      n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, 
      n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, 
      n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, 
      n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, 
      n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, 
      n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, 
      n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, 
      n1298, n1299, n1300, n1301, n1302, n2327, n2328, n2329, n2330, n2331, 
      n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, 
      n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, 
      n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, 
      n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, 
      n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, 
      n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, 
      n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, 
      n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, 
      n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, 
      n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, 
      n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, 
      n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, 
      n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, 
      n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, 
      n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, 
      n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, 
      n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, 
      n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, 
      n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, 
      n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, 
      n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, 
      n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, 
      n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, 
      n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, 
      n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, 
      n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
      n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, 
      n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, 
      n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, 
      n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
      n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, 
      n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, 
      n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, 
      n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, 
      n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, 
      n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, 
      n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, 
      n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, 
      n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, 
      n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, 
      n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, 
      n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, 
      n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, 
      n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, 
      n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, 
      n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, 
      n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, 
      n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, 
      n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, 
      n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, 
      n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, 
      n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, 
      n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, 
      n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, 
      n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, 
      n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, 
      n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
      n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, 
      n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, 
      n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, 
      n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, 
      n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, 
      n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, 
      n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, 
      n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, 
      n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, 
      n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, 
      n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, 
      n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, 
      n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, 
      n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, 
      n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, 
      n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, 
      n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, 
      n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, 
      n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
      n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, 
      n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, 
      n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, 
      n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, 
      n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, 
      n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, 
      n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, 
      n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, 
      n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, 
      n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, 
      n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, 
      n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, 
      n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, 
      n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, 
      n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, 
      n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, 
      n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, 
      n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, 
      n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
      n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, 
      n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, 
      n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, 
      n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, 
      n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, 
      n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, 
      n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, 
      n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, 
      n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, 
      n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, 
      n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, 
      n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, 
      n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, 
      n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, 
      n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, 
      n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, 
      n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, 
      n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, 
      n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, 
      n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, 
      n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, 
      n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, 
      n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, 
      n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, 
      n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, 
      n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, 
      n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, 
      n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, 
      n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, 
      n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, 
      n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, 
      n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, 
      n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, 
      n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, 
      n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, 
      n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, 
      n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, 
      n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, 
      n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, 
      n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, 
      n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, 
      n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, 
      n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, 
      n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, 
      n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, 
      n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, 
      n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, 
      n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, 
      n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, 
      n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, 
      n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, 
      n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, 
      n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, 
      n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, 
      n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, 
      n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, 
      n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, 
      n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, 
      n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, 
      n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, 
      n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, 
      n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, 
      n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, 
      n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, 
      n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, 
      n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, 
      n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, 
      n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, 
      n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, 
      n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, 
      n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, 
      n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, 
      n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, 
      n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, 
      n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, 
      n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, 
      n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, 
      n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, 
      n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, 
      n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, 
      n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, 
      n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, 
      n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, 
      n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, 
      n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, 
      n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, 
      n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, 
      n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, 
      n4162 : std_logic;

begin
   
   OUT2_reg_31_inst : DFF_X1 port map( D => n4130, CK => n293, Q => OUT2(31), 
                           QN => n3074);
   OUT2_reg_30_inst : DFF_X1 port map( D => n4129, CK => n320, Q => OUT2(30), 
                           QN => n3073);
   OUT2_reg_29_inst : DFF_X1 port map( D => n4128, CK => n314, Q => OUT2(29), 
                           QN => n3072);
   OUT2_reg_28_inst : DFF_X1 port map( D => n4127, CK => n323, Q => OUT2(28), 
                           QN => n3071);
   OUT2_reg_27_inst : DFF_X1 port map( D => n4126, CK => n327, Q => OUT2(27), 
                           QN => n3070);
   OUT2_reg_26_inst : DFF_X1 port map( D => n4125, CK => n330, Q => OUT2(26), 
                           QN => n3069);
   OUT2_reg_25_inst : DFF_X1 port map( D => n4124, CK => n305, Q => OUT2(25), 
                           QN => n3068);
   OUT2_reg_24_inst : DFF_X1 port map( D => n4123, CK => n333, Q => OUT2(24), 
                           QN => n3067);
   OUT2_reg_23_inst : DFF_X1 port map( D => n4122, CK => n336, Q => OUT2(23), 
                           QN => n3066);
   OUT2_reg_22_inst : DFF_X1 port map( D => n4121, CK => n339, Q => OUT2(22), 
                           QN => n3065);
   OUT2_reg_21_inst : DFF_X1 port map( D => n4120, CK => n293, Q => OUT2(21), 
                           QN => n3064);
   OUT2_reg_20_inst : DFF_X1 port map( D => n4119, CK => n342, Q => OUT2(20), 
                           QN => n3063);
   OUT2_reg_19_inst : DFF_X1 port map( D => n4118, CK => n345, Q => OUT2(19), 
                           QN => n3062);
   OUT2_reg_18_inst : DFF_X1 port map( D => n4117, CK => n348, Q => OUT2(18), 
                           QN => n3061);
   OUT2_reg_17_inst : DFF_X1 port map( D => n4116, CK => n293, Q => OUT2(17), 
                           QN => n3060);
   OUT2_reg_16_inst : DFF_X1 port map( D => n4115, CK => n351, Q => OUT2(16), 
                           QN => n3059);
   OUT2_reg_15_inst : DFF_X1 port map( D => n4114, CK => n354, Q => OUT2(15), 
                           QN => n3058);
   OUT2_reg_14_inst : DFF_X1 port map( D => n4113, CK => n357, Q => OUT2(14), 
                           QN => n3057);
   OUT2_reg_13_inst : DFF_X1 port map( D => n4112, CK => n296, Q => OUT2(13), 
                           QN => n3056);
   OUT2_reg_12_inst : DFF_X1 port map( D => n4111, CK => n361, Q => OUT2(12), 
                           QN => n3055);
   OUT2_reg_11_inst : DFF_X1 port map( D => n4110, CK => n364, Q => OUT2(11), 
                           QN => n3054);
   OUT2_reg_10_inst : DFF_X1 port map( D => n4109, CK => n367, Q => OUT2(10), 
                           QN => n3053);
   OUT2_reg_9_inst : DFF_X1 port map( D => n4108, CK => n308, Q => OUT2(9), QN 
                           => n3052);
   OUT2_reg_8_inst : DFF_X1 port map( D => n4107, CK => n370, Q => OUT2(8), QN 
                           => n3051);
   OUT2_reg_7_inst : DFF_X1 port map( D => n4106, CK => n373, Q => OUT2(7), QN 
                           => n3050);
   OUT2_reg_6_inst : DFF_X1 port map( D => n4105, CK => n376, Q => OUT2(6), QN 
                           => n3049);
   OUT2_reg_5_inst : DFF_X1 port map( D => n4104, CK => n293, Q => OUT2(5), QN 
                           => n3048);
   OUT2_reg_4_inst : DFF_X1 port map( D => n4103, CK => n379, Q => OUT2(4), QN 
                           => n3047);
   OUT2_reg_3_inst : DFF_X1 port map( D => n4102, CK => n382, Q => OUT2(3), QN 
                           => n3046);
   OUT2_reg_2_inst : DFF_X1 port map( D => n4101, CK => n385, Q => OUT2(2), QN 
                           => n3045);
   OUT2_reg_1_inst : DFF_X1 port map( D => n4100, CK => n311, Q => OUT2(1), QN 
                           => n3044);
   OUT2_reg_0_inst : DFF_X1 port map( D => n4099, CK => n388, Q => OUT2(0), QN 
                           => n3043);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2326, CK => n317, Q => 
                           REGISTERS_0_31_port, QN => n4098);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2325, CK => n321, Q => 
                           REGISTERS_0_30_port, QN => n4097);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2324, CK => n314, Q => 
                           REGISTERS_0_29_port, QN => n4096);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2323, CK => n324, Q => 
                           REGISTERS_0_28_port, QN => n4095);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2322, CK => n327, Q => 
                           REGISTERS_0_27_port, QN => n4094);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2321, CK => n330, Q => 
                           REGISTERS_0_26_port, QN => n4093);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2320, CK => n305, Q => 
                           REGISTERS_0_25_port, QN => n4092);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2319, CK => n333, Q => 
                           REGISTERS_0_24_port, QN => n4091);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2318, CK => n336, Q => 
                           REGISTERS_0_23_port, QN => n4090);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2317, CK => n339, Q => 
                           REGISTERS_0_22_port, QN => n4089);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2316, CK => n302, Q => 
                           REGISTERS_0_21_port, QN => n4088);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2315, CK => n342, Q => 
                           REGISTERS_0_20_port, QN => n4087);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2314, CK => n345, Q => 
                           REGISTERS_0_19_port, QN => n4086);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2313, CK => n348, Q => 
                           REGISTERS_0_18_port, QN => n4085);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2312, CK => n293, Q => 
                           REGISTERS_0_17_port, QN => n4084);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2311, CK => n351, Q => 
                           REGISTERS_0_16_port, QN => n4083);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2310, CK => n355, Q => 
                           REGISTERS_0_15_port, QN => n4082);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2309, CK => n358, Q => 
                           REGISTERS_0_14_port, QN => n4081);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2308, CK => n296, Q => 
                           REGISTERS_0_13_port, QN => n4080);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2307, CK => n361, Q => 
                           REGISTERS_0_12_port, QN => n4079);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2306, CK => n364, Q => 
                           REGISTERS_0_11_port, QN => n4078);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2305, CK => n367, Q => 
                           REGISTERS_0_10_port, QN => n4077);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2304, CK => n308, Q => 
                           REGISTERS_0_9_port, QN => n4076);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2303, CK => n370, Q => 
                           REGISTERS_0_8_port, QN => n4075);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2302, CK => n373, Q => 
                           REGISTERS_0_7_port, QN => n4074);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2301, CK => n376, Q => 
                           REGISTERS_0_6_port, QN => n4073);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2300, CK => n299, Q => 
                           REGISTERS_0_5_port, QN => n4072);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2299, CK => n379, Q => 
                           REGISTERS_0_4_port, QN => n4071);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2298, CK => n382, Q => 
                           REGISTERS_0_3_port, QN => n4070);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2297, CK => n385, Q => 
                           REGISTERS_0_2_port, QN => n4069);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2296, CK => n311, Q => 
                           REGISTERS_0_1_port, QN => n4068);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2295, CK => n389, Q => 
                           REGISTERS_0_0_port, QN => n4067);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2294, CK => n318, Q => 
                           REGISTERS_1_31_port, QN => n4066);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2293, CK => n321, Q => 
                           REGISTERS_1_30_port, QN => n4065);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2292, CK => n315, Q => 
                           REGISTERS_1_29_port, QN => n4064);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2291, CK => n324, Q => 
                           REGISTERS_1_28_port, QN => n4063);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2290, CK => n327, Q => 
                           REGISTERS_1_27_port, QN => n4062);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2289, CK => n330, Q => 
                           REGISTERS_1_26_port, QN => n4061);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2288, CK => n305, Q => 
                           REGISTERS_1_25_port, QN => n4060);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2287, CK => n333, Q => 
                           REGISTERS_1_24_port, QN => n4059);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2286, CK => n336, Q => 
                           REGISTERS_1_23_port, QN => n4058);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2285, CK => n339, Q => 
                           REGISTERS_1_22_port, QN => n4057);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2284, CK => n302, Q => 
                           REGISTERS_1_21_port, QN => n4056);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2283, CK => n342, Q => 
                           REGISTERS_1_20_port, QN => n4055);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2282, CK => n345, Q => 
                           REGISTERS_1_19_port, QN => n4054);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2281, CK => n348, Q => 
                           REGISTERS_1_18_port, QN => n4053);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2280, CK => n293, Q => 
                           REGISTERS_1_17_port, QN => n4052);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2279, CK => n352, Q => 
                           REGISTERS_1_16_port, QN => n4051);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2278, CK => n355, Q => 
                           REGISTERS_1_15_port, QN => n4050);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2277, CK => n358, Q => 
                           REGISTERS_1_14_port, QN => n4049);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2276, CK => n296, Q => 
                           REGISTERS_1_13_port, QN => n4048);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2275, CK => n361, Q => 
                           REGISTERS_1_12_port, QN => n4047);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2274, CK => n364, Q => 
                           REGISTERS_1_11_port, QN => n4046);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2273, CK => n367, Q => 
                           REGISTERS_1_10_port, QN => n4045);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2272, CK => n308, Q => 
                           REGISTERS_1_9_port, QN => n4044);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2271, CK => n370, Q => 
                           REGISTERS_1_8_port, QN => n4043);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2270, CK => n373, Q => 
                           REGISTERS_1_7_port, QN => n4042);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2269, CK => n376, Q => 
                           REGISTERS_1_6_port, QN => n4041);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2268, CK => n299, Q => 
                           REGISTERS_1_5_port, QN => n4040);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2267, CK => n379, Q => 
                           REGISTERS_1_4_port, QN => n4039);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2266, CK => n382, Q => 
                           REGISTERS_1_3_port, QN => n4038);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2265, CK => n386, Q => 
                           REGISTERS_1_2_port, QN => n4037);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2264, CK => n311, Q => 
                           REGISTERS_1_1_port, QN => n4036);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2263, CK => n389, Q => 
                           REGISTERS_1_0_port, QN => n4035);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2262, CK => n318, Q => 
                           REGISTERS_2_31_port, QN => n4034);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2261, CK => n321, Q => 
                           REGISTERS_2_30_port, QN => n4033);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2260, CK => n315, Q => 
                           REGISTERS_2_29_port, QN => n4032);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2259, CK => n324, Q => 
                           REGISTERS_2_28_port, QN => n4031);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2258, CK => n327, Q => 
                           REGISTERS_2_27_port, QN => n4030);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2257, CK => n330, Q => 
                           REGISTERS_2_26_port, QN => n4029);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2256, CK => n305, Q => 
                           REGISTERS_2_25_port, QN => n4028);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2255, CK => n333, Q => 
                           REGISTERS_2_24_port, QN => n4027);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2254, CK => n336, Q => 
                           REGISTERS_2_23_port, QN => n4026);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2253, CK => n339, Q => 
                           REGISTERS_2_22_port, QN => n4025);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2252, CK => n302, Q => 
                           REGISTERS_2_21_port, QN => n4024);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2251, CK => n342, Q => 
                           REGISTERS_2_20_port, QN => n4023);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2250, CK => n345, Q => 
                           REGISTERS_2_19_port, QN => n4022);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2249, CK => n349, Q => 
                           REGISTERS_2_18_port, QN => n4021);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2248, CK => n293, Q => 
                           REGISTERS_2_17_port, QN => n4020);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2247, CK => n352, Q => 
                           REGISTERS_2_16_port, QN => n4019);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2246, CK => n355, Q => 
                           REGISTERS_2_15_port, QN => n4018);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2245, CK => n358, Q => 
                           REGISTERS_2_14_port, QN => n4017);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2244, CK => n296, Q => 
                           REGISTERS_2_13_port, QN => n4016);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2243, CK => n361, Q => 
                           REGISTERS_2_12_port, QN => n4015);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2242, CK => n364, Q => 
                           REGISTERS_2_11_port, QN => n4014);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2241, CK => n367, Q => 
                           REGISTERS_2_10_port, QN => n4013);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2240, CK => n308, Q => 
                           REGISTERS_2_9_port, QN => n4012);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2239, CK => n370, Q => 
                           REGISTERS_2_8_port, QN => n4011);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2238, CK => n373, Q => 
                           REGISTERS_2_7_port, QN => n4010);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2237, CK => n376, Q => 
                           REGISTERS_2_6_port, QN => n4009);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2236, CK => n299, Q => 
                           REGISTERS_2_5_port, QN => n4008);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2235, CK => n379, Q => 
                           REGISTERS_2_4_port, QN => n4007);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2234, CK => n383, Q => 
                           REGISTERS_2_3_port, QN => n4006);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2233, CK => n386, Q => 
                           REGISTERS_2_2_port, QN => n4005);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2232, CK => n312, Q => 
                           REGISTERS_2_1_port, QN => n4004);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2231, CK => n389, Q => 
                           REGISTERS_2_0_port, QN => n4003);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2230, CK => n318, Q => 
                           REGISTERS_3_31_port, QN => n4002);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2229, CK => n321, Q => 
                           REGISTERS_3_30_port, QN => n4001);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2228, CK => n315, Q => 
                           REGISTERS_3_29_port, QN => n4000);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2227, CK => n324, Q => 
                           REGISTERS_3_28_port, QN => n3999);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2226, CK => n327, Q => 
                           REGISTERS_3_27_port, QN => n3998);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2225, CK => n330, Q => 
                           REGISTERS_3_26_port, QN => n3997);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2224, CK => n305, Q => 
                           REGISTERS_3_25_port, QN => n3996);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2223, CK => n333, Q => 
                           REGISTERS_3_24_port, QN => n3995);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2222, CK => n336, Q => 
                           REGISTERS_3_23_port, QN => n3994);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2221, CK => n339, Q => 
                           REGISTERS_3_22_port, QN => n3993);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2220, CK => n302, Q => 
                           REGISTERS_3_21_port, QN => n3992);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2219, CK => n342, Q => 
                           REGISTERS_3_20_port, QN => n3991);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2218, CK => n346, Q => 
                           REGISTERS_3_19_port, QN => n3990);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2217, CK => n349, Q => 
                           REGISTERS_3_18_port, QN => n3989);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2216, CK => n293, Q => 
                           REGISTERS_3_17_port, QN => n3988);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2215, CK => n352, Q => 
                           REGISTERS_3_16_port, QN => n3987);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2214, CK => n355, Q => 
                           REGISTERS_3_15_port, QN => n3986);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2213, CK => n358, Q => 
                           REGISTERS_3_14_port, QN => n3985);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2212, CK => n296, Q => 
                           REGISTERS_3_13_port, QN => n3984);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2211, CK => n361, Q => 
                           REGISTERS_3_12_port, QN => n3983);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2210, CK => n364, Q => 
                           REGISTERS_3_11_port, QN => n3982);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2209, CK => n367, Q => 
                           REGISTERS_3_10_port, QN => n3981);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2208, CK => n309, Q => 
                           REGISTERS_3_9_port, QN => n3980);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2207, CK => n370, Q => 
                           REGISTERS_3_8_port, QN => n3979);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2206, CK => n373, Q => 
                           REGISTERS_3_7_port, QN => n3978);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2205, CK => n376, Q => 
                           REGISTERS_3_6_port, QN => n3977);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2204, CK => n299, Q => 
                           REGISTERS_3_5_port, QN => n3976);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2203, CK => n380, Q => 
                           REGISTERS_3_4_port, QN => n3975);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2202, CK => n383, Q => 
                           REGISTERS_3_3_port, QN => n3974);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2201, CK => n386, Q => 
                           REGISTERS_3_2_port, QN => n3973);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2200, CK => n312, Q => 
                           REGISTERS_3_1_port, QN => n3972);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2199, CK => n389, Q => 
                           REGISTERS_3_0_port, QN => n3971);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2198, CK => n318, Q => 
                           REGISTERS_4_31_port, QN => n3970);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2197, CK => n321, Q => 
                           REGISTERS_4_30_port, QN => n3969);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2196, CK => n315, Q => 
                           REGISTERS_4_29_port, QN => n3968);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2195, CK => n324, Q => 
                           REGISTERS_4_28_port, QN => n3967);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2194, CK => n327, Q => 
                           REGISTERS_4_27_port, QN => n3966);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2193, CK => n330, Q => 
                           REGISTERS_4_26_port, QN => n3965);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2192, CK => n306, Q => 
                           REGISTERS_4_25_port, QN => n3964);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2191, CK => n333, Q => 
                           REGISTERS_4_24_port, QN => n3963);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2190, CK => n336, Q => 
                           REGISTERS_4_23_port, QN => n3962);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2189, CK => n339, Q => 
                           REGISTERS_4_22_port, QN => n3961);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2188, CK => n302, Q => 
                           REGISTERS_4_21_port, QN => n3960);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2187, CK => n343, Q => 
                           REGISTERS_4_20_port, QN => n3959);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2186, CK => n346, Q => 
                           REGISTERS_4_19_port, QN => n3958);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2185, CK => n349, Q => 
                           REGISTERS_4_18_port, QN => n3957);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2184, CK => n293, Q => 
                           REGISTERS_4_17_port, QN => n3956);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2183, CK => n352, Q => 
                           REGISTERS_4_16_port, QN => n3955);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2182, CK => n355, Q => 
                           REGISTERS_4_15_port, QN => n3954);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2181, CK => n358, Q => 
                           REGISTERS_4_14_port, QN => n3953);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2180, CK => n296, Q => 
                           REGISTERS_4_13_port, QN => n3952);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2179, CK => n361, Q => 
                           REGISTERS_4_12_port, QN => n3951);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2178, CK => n364, Q => 
                           REGISTERS_4_11_port, QN => n3950);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2177, CK => n367, Q => 
                           REGISTERS_4_10_port, QN => n3949);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2176, CK => n309, Q => 
                           REGISTERS_4_9_port, QN => n3948);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2175, CK => n370, Q => 
                           REGISTERS_4_8_port, QN => n3947);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2174, CK => n373, Q => 
                           REGISTERS_4_7_port, QN => n3946);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2173, CK => n377, Q => 
                           REGISTERS_4_6_port, QN => n3945);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2172, CK => n299, Q => 
                           REGISTERS_4_5_port, QN => n3944);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2171, CK => n380, Q => 
                           REGISTERS_4_4_port, QN => n3943);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2170, CK => n383, Q => 
                           REGISTERS_4_3_port, QN => n3942);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2169, CK => n386, Q => 
                           REGISTERS_4_2_port, QN => n3941);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2168, CK => n312, Q => 
                           REGISTERS_4_1_port, QN => n3940);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2167, CK => n389, Q => 
                           REGISTERS_4_0_port, QN => n3939);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2166, CK => n318, Q => 
                           REGISTERS_5_31_port, QN => n3938);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2165, CK => n321, Q => 
                           REGISTERS_5_30_port, QN => n3937);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2164, CK => n315, Q => 
                           REGISTERS_5_29_port, QN => n3936);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2163, CK => n324, Q => 
                           REGISTERS_5_28_port, QN => n3935);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2162, CK => n327, Q => 
                           REGISTERS_5_27_port, QN => n3934);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2161, CK => n330, Q => 
                           REGISTERS_5_26_port, QN => n3933);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2160, CK => n306, Q => 
                           REGISTERS_5_25_port, QN => n3932);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n2159, CK => n333, Q => 
                           REGISTERS_5_24_port, QN => n3931);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n2158, CK => n336, Q => 
                           REGISTERS_5_23_port, QN => n3930);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n2157, CK => n340, Q => 
                           REGISTERS_5_22_port, QN => n3929);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n2156, CK => n303, Q => 
                           REGISTERS_5_21_port, QN => n3928);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n2155, CK => n343, Q => 
                           REGISTERS_5_20_port, QN => n3927);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n2154, CK => n346, Q => 
                           REGISTERS_5_19_port, QN => n3926);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n2153, CK => n349, Q => 
                           REGISTERS_5_18_port, QN => n3925);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n2152, CK => n293, Q => 
                           REGISTERS_5_17_port, QN => n3924);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n2151, CK => n352, Q => 
                           REGISTERS_5_16_port, QN => n3923);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n2150, CK => n355, Q => 
                           REGISTERS_5_15_port, QN => n3922);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n2149, CK => n358, Q => 
                           REGISTERS_5_14_port, QN => n3921);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n2148, CK => n297, Q => 
                           REGISTERS_5_13_port, QN => n3920);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n2147, CK => n361, Q => 
                           REGISTERS_5_12_port, QN => n3919);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n2146, CK => n364, Q => 
                           REGISTERS_5_11_port, QN => n3918);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n2145, CK => n367, Q => 
                           REGISTERS_5_10_port, QN => n3917);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n2144, CK => n309, Q => 
                           REGISTERS_5_9_port, QN => n3916);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n2143, CK => n370, Q => 
                           REGISTERS_5_8_port, QN => n3915);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n2142, CK => n374, Q => 
                           REGISTERS_5_7_port, QN => n3914);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n2141, CK => n377, Q => 
                           REGISTERS_5_6_port, QN => n3913);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n2140, CK => n300, Q => 
                           REGISTERS_5_5_port, QN => n3912);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n2139, CK => n380, Q => 
                           REGISTERS_5_4_port, QN => n3911);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n2138, CK => n383, Q => 
                           REGISTERS_5_3_port, QN => n3910);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n2137, CK => n386, Q => 
                           REGISTERS_5_2_port, QN => n3909);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n2136, CK => n312, Q => 
                           REGISTERS_5_1_port, QN => n3908);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n2135, CK => n389, Q => 
                           REGISTERS_5_0_port, QN => n3907);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n2134, CK => n318, Q => 
                           REGISTERS_6_31_port, QN => n3906);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n2133, CK => n321, Q => 
                           REGISTERS_6_30_port, QN => n3905);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n2132, CK => n315, Q => 
                           REGISTERS_6_29_port, QN => n3904);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n2131, CK => n324, Q => 
                           REGISTERS_6_28_port, QN => n3903);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n2130, CK => n327, Q => 
                           REGISTERS_6_27_port, QN => n3902);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n2129, CK => n330, Q => 
                           REGISTERS_6_26_port, QN => n3901);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n2128, CK => n306, Q => 
                           REGISTERS_6_25_port, QN => n3900);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n2127, CK => n333, Q => 
                           REGISTERS_6_24_port, QN => n3899);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n2126, CK => n337, Q => 
                           REGISTERS_6_23_port, QN => n3898);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n2125, CK => n340, Q => 
                           REGISTERS_6_22_port, QN => n3897);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n2124, CK => n303, Q => 
                           REGISTERS_6_21_port, QN => n3896);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n2123, CK => n343, Q => 
                           REGISTERS_6_20_port, QN => n3895);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n2122, CK => n346, Q => 
                           REGISTERS_6_19_port, QN => n3894);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n2121, CK => n349, Q => 
                           REGISTERS_6_18_port, QN => n3893);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n2120, CK => n294, Q => 
                           REGISTERS_6_17_port, QN => n3892);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n2119, CK => n352, Q => 
                           REGISTERS_6_16_port, QN => n3891);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n2118, CK => n355, Q => 
                           REGISTERS_6_15_port, QN => n3890);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n2117, CK => n358, Q => 
                           REGISTERS_6_14_port, QN => n3889);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n2116, CK => n297, Q => 
                           REGISTERS_6_13_port, QN => n3888);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n2115, CK => n361, Q => 
                           REGISTERS_6_12_port, QN => n3887);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n2114, CK => n364, Q => 
                           REGISTERS_6_11_port, QN => n3886);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n2113, CK => n367, Q => 
                           REGISTERS_6_10_port, QN => n3885);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n2112, CK => n309, Q => 
                           REGISTERS_6_9_port, QN => n3884);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n2111, CK => n371, Q => 
                           REGISTERS_6_8_port, QN => n3883);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n2110, CK => n374, Q => 
                           REGISTERS_6_7_port, QN => n3882);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n2109, CK => n377, Q => 
                           REGISTERS_6_6_port, QN => n3881);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n2108, CK => n300, Q => 
                           REGISTERS_6_5_port, QN => n3880);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n2107, CK => n380, Q => 
                           REGISTERS_6_4_port, QN => n3879);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n2106, CK => n383, Q => 
                           REGISTERS_6_3_port, QN => n3878);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n2105, CK => n386, Q => 
                           REGISTERS_6_2_port, QN => n3877);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n2104, CK => n312, Q => 
                           REGISTERS_6_1_port, QN => n3876);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n2103, CK => n389, Q => 
                           REGISTERS_6_0_port, QN => n3875);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n2102, CK => n318, Q => 
                           REGISTERS_7_31_port, QN => n3874);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n2101, CK => n321, Q => 
                           REGISTERS_7_30_port, QN => n3873);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n2100, CK => n315, Q => 
                           REGISTERS_7_29_port, QN => n3872);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n2099, CK => n324, Q => 
                           REGISTERS_7_28_port, QN => n3871);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n2098, CK => n327, Q => 
                           REGISTERS_7_27_port, QN => n3870);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n2097, CK => n330, Q => 
                           REGISTERS_7_26_port, QN => n3869);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n2096, CK => n306, Q => 
                           REGISTERS_7_25_port, QN => n3868);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n2095, CK => n334, Q => 
                           REGISTERS_7_24_port, QN => n3867);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n2094, CK => n337, Q => 
                           REGISTERS_7_23_port, QN => n3866);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n2093, CK => n340, Q => 
                           REGISTERS_7_22_port, QN => n3865);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n2092, CK => n303, Q => 
                           REGISTERS_7_21_port, QN => n3864);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n2091, CK => n343, Q => 
                           REGISTERS_7_20_port, QN => n3863);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n2090, CK => n346, Q => 
                           REGISTERS_7_19_port, QN => n3862);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n2089, CK => n349, Q => 
                           REGISTERS_7_18_port, QN => n3861);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n2088, CK => n294, Q => 
                           REGISTERS_7_17_port, QN => n3860);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n2087, CK => n352, Q => 
                           REGISTERS_7_16_port, QN => n3859);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n2086, CK => n355, Q => 
                           REGISTERS_7_15_port, QN => n3858);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n2085, CK => n358, Q => 
                           REGISTERS_7_14_port, QN => n3857);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n2084, CK => n297, Q => 
                           REGISTERS_7_13_port, QN => n3856);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n2083, CK => n361, Q => 
                           REGISTERS_7_12_port, QN => n3855);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n2082, CK => n364, Q => 
                           REGISTERS_7_11_port, QN => n3854);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n2081, CK => n368, Q => 
                           REGISTERS_7_10_port, QN => n3853);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n2080, CK => n309, Q => 
                           REGISTERS_7_9_port, QN => n3852);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n2079, CK => n371, Q => 
                           REGISTERS_7_8_port, QN => n3851);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n2078, CK => n374, Q => 
                           REGISTERS_7_7_port, QN => n3850);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n2077, CK => n377, Q => 
                           REGISTERS_7_6_port, QN => n3849);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n2076, CK => n300, Q => 
                           REGISTERS_7_5_port, QN => n3848);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n2075, CK => n380, Q => 
                           REGISTERS_7_4_port, QN => n3847);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n2074, CK => n383, Q => 
                           REGISTERS_7_3_port, QN => n3846);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n2073, CK => n386, Q => 
                           REGISTERS_7_2_port, QN => n3845);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n2072, CK => n312, Q => 
                           REGISTERS_7_1_port, QN => n3844);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n2071, CK => n389, Q => 
                           REGISTERS_7_0_port, QN => n3843);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n2070, CK => n318, Q => 
                           REGISTERS_8_31_port, QN => n3842);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n2069, CK => n321, Q => 
                           REGISTERS_8_30_port, QN => n3841);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n2068, CK => n315, Q => 
                           REGISTERS_8_29_port, QN => n3840);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n2067, CK => n324, Q => 
                           REGISTERS_8_28_port, QN => n3839);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n2066, CK => n327, Q => 
                           REGISTERS_8_27_port, QN => n3838);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n2065, CK => n331, Q => 
                           REGISTERS_8_26_port, QN => n3837);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n2064, CK => n306, Q => 
                           REGISTERS_8_25_port, QN => n3836);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n2063, CK => n334, Q => 
                           REGISTERS_8_24_port, QN => n3835);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n2062, CK => n337, Q => 
                           REGISTERS_8_23_port, QN => n3834);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n2061, CK => n340, Q => 
                           REGISTERS_8_22_port, QN => n3833);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n2060, CK => n303, Q => 
                           REGISTERS_8_21_port, QN => n3832);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n2059, CK => n343, Q => 
                           REGISTERS_8_20_port, QN => n3831);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n2058, CK => n346, Q => 
                           REGISTERS_8_19_port, QN => n3830);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n2057, CK => n349, Q => 
                           REGISTERS_8_18_port, QN => n3829);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n2056, CK => n294, Q => 
                           REGISTERS_8_17_port, QN => n3828);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n2055, CK => n352, Q => 
                           REGISTERS_8_16_port, QN => n3827);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n2054, CK => n355, Q => 
                           REGISTERS_8_15_port, QN => n3826);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n2053, CK => n358, Q => 
                           REGISTERS_8_14_port, QN => n3825);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n2052, CK => n297, Q => 
                           REGISTERS_8_13_port, QN => n3824);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n2051, CK => n361, Q => 
                           REGISTERS_8_12_port, QN => n3823);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n2050, CK => n365, Q => 
                           REGISTERS_8_11_port, QN => n3822);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n2049, CK => n368, Q => 
                           REGISTERS_8_10_port, QN => n3821);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n2048, CK => n309, Q => 
                           REGISTERS_8_9_port, QN => n3820);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n2047, CK => n371, Q => 
                           REGISTERS_8_8_port, QN => n3819);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n2046, CK => n374, Q => 
                           REGISTERS_8_7_port, QN => n3818);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n2045, CK => n377, Q => 
                           REGISTERS_8_6_port, QN => n3817);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n2044, CK => n300, Q => 
                           REGISTERS_8_5_port, QN => n3816);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n2043, CK => n380, Q => 
                           REGISTERS_8_4_port, QN => n3815);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n2042, CK => n383, Q => 
                           REGISTERS_8_3_port, QN => n3814);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n2041, CK => n386, Q => 
                           REGISTERS_8_2_port, QN => n3813);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n2040, CK => n312, Q => 
                           REGISTERS_8_1_port, QN => n3812);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n2039, CK => n389, Q => 
                           REGISTERS_8_0_port, QN => n3811);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n2038, CK => n318, Q => 
                           REGISTERS_9_31_port, QN => n3810);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n2037, CK => n321, Q => 
                           REGISTERS_9_30_port, QN => n3809);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n2036, CK => n315, Q => 
                           REGISTERS_9_29_port, QN => n3808);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n2035, CK => n324, Q => 
                           REGISTERS_9_28_port, QN => n3807);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n2034, CK => n328, Q => 
                           REGISTERS_9_27_port, QN => n3806);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n2033, CK => n331, Q => 
                           REGISTERS_9_26_port, QN => n3805);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n2032, CK => n306, Q => 
                           REGISTERS_9_25_port, QN => n3804);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n2031, CK => n334, Q => 
                           REGISTERS_9_24_port, QN => n3803);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n2030, CK => n337, Q => 
                           REGISTERS_9_23_port, QN => n3802);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n2029, CK => n340, Q => 
                           REGISTERS_9_22_port, QN => n3801);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n2028, CK => n303, Q => 
                           REGISTERS_9_21_port, QN => n3800);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n2027, CK => n343, Q => 
                           REGISTERS_9_20_port, QN => n3799);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n2026, CK => n346, Q => 
                           REGISTERS_9_19_port, QN => n3798);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n2025, CK => n349, Q => 
                           REGISTERS_9_18_port, QN => n3797);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n2024, CK => n294, Q => 
                           REGISTERS_9_17_port, QN => n3796);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n2023, CK => n352, Q => 
                           REGISTERS_9_16_port, QN => n3795);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n2022, CK => n355, Q => 
                           REGISTERS_9_15_port, QN => n3794);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n2021, CK => n358, Q => 
                           REGISTERS_9_14_port, QN => n3793);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n2020, CK => n297, Q => 
                           REGISTERS_9_13_port, QN => n3792);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n2019, CK => n362, Q => 
                           REGISTERS_9_12_port, QN => n3791);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n2018, CK => n365, Q => 
                           REGISTERS_9_11_port, QN => n3790);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n2017, CK => n368, Q => 
                           REGISTERS_9_10_port, QN => n3789);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n2016, CK => n309, Q => 
                           REGISTERS_9_9_port, QN => n3788);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n2015, CK => n371, Q => 
                           REGISTERS_9_8_port, QN => n3787);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n2014, CK => n374, Q => 
                           REGISTERS_9_7_port, QN => n3786);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n2013, CK => n377, Q => 
                           REGISTERS_9_6_port, QN => n3785);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n2012, CK => n300, Q => 
                           REGISTERS_9_5_port, QN => n3784);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n2011, CK => n380, Q => 
                           REGISTERS_9_4_port, QN => n3783);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n2010, CK => n383, Q => 
                           REGISTERS_9_3_port, QN => n3782);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n2009, CK => n386, Q => 
                           REGISTERS_9_2_port, QN => n3781);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n2008, CK => n312, Q => 
                           REGISTERS_9_1_port, QN => n3780);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n2007, CK => n389, Q => 
                           REGISTERS_9_0_port, QN => n3779);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n2006, CK => n318, Q => 
                           REGISTERS_10_31_port, QN => n3778);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n2005, CK => n321, Q => 
                           REGISTERS_10_30_port, QN => n3777);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n2004, CK => n315, Q => 
                           REGISTERS_10_29_port, QN => n3776);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n2003, CK => n325, Q => 
                           REGISTERS_10_28_port, QN => n3775);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n2002, CK => n328, Q => 
                           REGISTERS_10_27_port, QN => n3774);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n2001, CK => n331, Q => 
                           REGISTERS_10_26_port, QN => n3773);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n2000, CK => n306, Q => 
                           REGISTERS_10_25_port, QN => n3772);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1999, CK => n334, Q => 
                           REGISTERS_10_24_port, QN => n3771);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1998, CK => n337, Q => 
                           REGISTERS_10_23_port, QN => n3770);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1997, CK => n340, Q => 
                           REGISTERS_10_22_port, QN => n3769);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1996, CK => n303, Q => 
                           REGISTERS_10_21_port, QN => n3768);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1995, CK => n343, Q => 
                           REGISTERS_10_20_port, QN => n3767);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1994, CK => n346, Q => 
                           REGISTERS_10_19_port, QN => n3766);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1993, CK => n349, Q => 
                           REGISTERS_10_18_port, QN => n3765);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1992, CK => n294, Q => 
                           REGISTERS_10_17_port, QN => n3764);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1991, CK => n352, Q => 
                           REGISTERS_10_16_port, QN => n3763);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1990, CK => n355, Q => 
                           REGISTERS_10_15_port, QN => n3762);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1989, CK => n359, Q => 
                           REGISTERS_10_14_port, QN => n3761);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1988, CK => n297, Q => 
                           REGISTERS_10_13_port, QN => n3760);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1987, CK => n362, Q => 
                           REGISTERS_10_12_port, QN => n3759);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1986, CK => n365, Q => 
                           REGISTERS_10_11_port, QN => n3758);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1985, CK => n368, Q => 
                           REGISTERS_10_10_port, QN => n3757);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1984, CK => n309, Q => 
                           REGISTERS_10_9_port, QN => n3756);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1983, CK => n371, Q => 
                           REGISTERS_10_8_port, QN => n3755);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1982, CK => n374, Q => 
                           REGISTERS_10_7_port, QN => n3754);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1981, CK => n377, Q => 
                           REGISTERS_10_6_port, QN => n3753);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1980, CK => n300, Q => 
                           REGISTERS_10_5_port, QN => n3752);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1979, CK => n380, Q => 
                           REGISTERS_10_4_port, QN => n3751);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1978, CK => n383, Q => 
                           REGISTERS_10_3_port, QN => n3750);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1977, CK => n386, Q => 
                           REGISTERS_10_2_port, QN => n3749);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1976, CK => n312, Q => 
                           REGISTERS_10_1_port, QN => n3748);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1975, CK => n389, Q => 
                           REGISTERS_10_0_port, QN => n3747);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1974, CK => n318, Q => 
                           REGISTERS_11_31_port, QN => n3746);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1973, CK => n322, Q => 
                           REGISTERS_11_30_port, QN => n3745);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1972, CK => n315, Q => 
                           REGISTERS_11_29_port, QN => n3744);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1971, CK => n325, Q => 
                           REGISTERS_11_28_port, QN => n3743);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1970, CK => n328, Q => 
                           REGISTERS_11_27_port, QN => n3742);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1969, CK => n331, Q => 
                           REGISTERS_11_26_port, QN => n3741);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1968, CK => n306, Q => 
                           REGISTERS_11_25_port, QN => n3740);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1967, CK => n334, Q => 
                           REGISTERS_11_24_port, QN => n3739);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1966, CK => n337, Q => 
                           REGISTERS_11_23_port, QN => n3738);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1965, CK => n340, Q => 
                           REGISTERS_11_22_port, QN => n3737);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1964, CK => n303, Q => 
                           REGISTERS_11_21_port, QN => n3736);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1963, CK => n343, Q => 
                           REGISTERS_11_20_port, QN => n3735);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1962, CK => n346, Q => 
                           REGISTERS_11_19_port, QN => n3734);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1961, CK => n349, Q => 
                           REGISTERS_11_18_port, QN => n3733);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1960, CK => n294, Q => 
                           REGISTERS_11_17_port, QN => n3732);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1959, CK => n352, Q => 
                           REGISTERS_11_16_port, QN => n3731);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1958, CK => n356, Q => 
                           REGISTERS_11_15_port, QN => n3730);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1957, CK => n359, Q => 
                           REGISTERS_11_14_port, QN => n3729);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1956, CK => n297, Q => 
                           REGISTERS_11_13_port, QN => n3728);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1955, CK => n362, Q => 
                           REGISTERS_11_12_port, QN => n3727);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1954, CK => n365, Q => 
                           REGISTERS_11_11_port, QN => n3726);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1953, CK => n368, Q => 
                           REGISTERS_11_10_port, QN => n3725);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1952, CK => n309, Q => 
                           REGISTERS_11_9_port, QN => n3724);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1951, CK => n371, Q => 
                           REGISTERS_11_8_port, QN => n3723);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1950, CK => n374, Q => 
                           REGISTERS_11_7_port, QN => n3722);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1949, CK => n377, Q => 
                           REGISTERS_11_6_port, QN => n3721);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1948, CK => n300, Q => 
                           REGISTERS_11_5_port, QN => n3720);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1947, CK => n380, Q => 
                           REGISTERS_11_4_port, QN => n3719);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1946, CK => n383, Q => 
                           REGISTERS_11_3_port, QN => n3718);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1945, CK => n386, Q => 
                           REGISTERS_11_2_port, QN => n3717);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1944, CK => n312, Q => 
                           REGISTERS_11_1_port, QN => n3716);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1943, CK => n390, Q => 
                           REGISTERS_11_0_port, QN => n3715);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1942, CK => n319, Q => 
                           REGISTERS_12_31_port, QN => n3714);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1941, CK => n322, Q => 
                           REGISTERS_12_30_port, QN => n3713);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1940, CK => n316, Q => 
                           REGISTERS_12_29_port, QN => n3712);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1939, CK => n325, Q => 
                           REGISTERS_12_28_port, QN => n3711);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1938, CK => n328, Q => 
                           REGISTERS_12_27_port, QN => n3710);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1937, CK => n331, Q => 
                           REGISTERS_12_26_port, QN => n3709);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1936, CK => n306, Q => 
                           REGISTERS_12_25_port, QN => n3708);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1935, CK => n334, Q => 
                           REGISTERS_12_24_port, QN => n3707);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1934, CK => n337, Q => 
                           REGISTERS_12_23_port, QN => n3706);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1933, CK => n340, Q => 
                           REGISTERS_12_22_port, QN => n3705);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1932, CK => n303, Q => 
                           REGISTERS_12_21_port, QN => n3704);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1931, CK => n343, Q => 
                           REGISTERS_12_20_port, QN => n3703);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1930, CK => n346, Q => 
                           REGISTERS_12_19_port, QN => n3702);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1929, CK => n349, Q => 
                           REGISTERS_12_18_port, QN => n3701);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1928, CK => n294, Q => 
                           REGISTERS_12_17_port, QN => n3700);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1927, CK => n353, Q => 
                           REGISTERS_12_16_port, QN => n3699);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1926, CK => n356, Q => 
                           REGISTERS_12_15_port, QN => n3698);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1925, CK => n359, Q => 
                           REGISTERS_12_14_port, QN => n3697);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1924, CK => n297, Q => 
                           REGISTERS_12_13_port, QN => n3696);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1923, CK => n362, Q => 
                           REGISTERS_12_12_port, QN => n3695);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1922, CK => n365, Q => 
                           REGISTERS_12_11_port, QN => n3694);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1921, CK => n368, Q => 
                           REGISTERS_12_10_port, QN => n3693);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1920, CK => n309, Q => 
                           REGISTERS_12_9_port, QN => n3692);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1919, CK => n371, Q => 
                           REGISTERS_12_8_port, QN => n3691);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1918, CK => n374, Q => 
                           REGISTERS_12_7_port, QN => n3690);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1917, CK => n377, Q => 
                           REGISTERS_12_6_port, QN => n3689);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1916, CK => n300, Q => 
                           REGISTERS_12_5_port, QN => n3688);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1915, CK => n380, Q => 
                           REGISTERS_12_4_port, QN => n3687);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1914, CK => n383, Q => 
                           REGISTERS_12_3_port, QN => n3686);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1913, CK => n387, Q => 
                           REGISTERS_12_2_port, QN => n3685);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1912, CK => n312, Q => 
                           REGISTERS_12_1_port, QN => n3684);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1911, CK => n390, Q => 
                           REGISTERS_12_0_port, QN => n3683);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1910, CK => n319, Q => 
                           REGISTERS_13_31_port, QN => n3682);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1909, CK => n322, Q => 
                           REGISTERS_13_30_port, QN => n3681);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1908, CK => n316, Q => 
                           REGISTERS_13_29_port, QN => n3680);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1907, CK => n325, Q => 
                           REGISTERS_13_28_port, QN => n3679);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1906, CK => n328, Q => 
                           REGISTERS_13_27_port, QN => n3678);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1905, CK => n331, Q => 
                           REGISTERS_13_26_port, QN => n3677);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1904, CK => n306, Q => 
                           REGISTERS_13_25_port, QN => n3676);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1903, CK => n334, Q => 
                           REGISTERS_13_24_port, QN => n3675);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1902, CK => n337, Q => 
                           REGISTERS_13_23_port, QN => n3674);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1901, CK => n340, Q => 
                           REGISTERS_13_22_port, QN => n3673);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1900, CK => n303, Q => 
                           REGISTERS_13_21_port, QN => n3672);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1899, CK => n343, Q => 
                           REGISTERS_13_20_port, QN => n3671);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1898, CK => n346, Q => 
                           REGISTERS_13_19_port, QN => n3670);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1897, CK => n350, Q => 
                           REGISTERS_13_18_port, QN => n3669);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1896, CK => n294, Q => 
                           REGISTERS_13_17_port, QN => n3668);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1895, CK => n353, Q => 
                           REGISTERS_13_16_port, QN => n3667);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1894, CK => n356, Q => 
                           REGISTERS_13_15_port, QN => n3666);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1893, CK => n359, Q => 
                           REGISTERS_13_14_port, QN => n3665);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1892, CK => n297, Q => 
                           REGISTERS_13_13_port, QN => n3664);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1891, CK => n362, Q => 
                           REGISTERS_13_12_port, QN => n3663);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1890, CK => n365, Q => 
                           REGISTERS_13_11_port, QN => n3662);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1889, CK => n368, Q => 
                           REGISTERS_13_10_port, QN => n3661);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1888, CK => n309, Q => 
                           REGISTERS_13_9_port, QN => n3660);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1887, CK => n371, Q => 
                           REGISTERS_13_8_port, QN => n3659);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1886, CK => n374, Q => 
                           REGISTERS_13_7_port, QN => n3658);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1885, CK => n377, Q => 
                           REGISTERS_13_6_port, QN => n3657);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1884, CK => n300, Q => 
                           REGISTERS_13_5_port, QN => n3656);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1883, CK => n380, Q => 
                           REGISTERS_13_4_port, QN => n3655);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1882, CK => n384, Q => 
                           REGISTERS_13_3_port, QN => n3654);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1881, CK => n387, Q => 
                           REGISTERS_13_2_port, QN => n3653);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1880, CK => n313, Q => 
                           REGISTERS_13_1_port, QN => n3652);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1879, CK => n390, Q => 
                           REGISTERS_13_0_port, QN => n3651);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1878, CK => n319, Q => 
                           REGISTERS_14_31_port, QN => n3650);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1877, CK => n322, Q => 
                           REGISTERS_14_30_port, QN => n3649);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1876, CK => n316, Q => 
                           REGISTERS_14_29_port, QN => n3648);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1875, CK => n325, Q => 
                           REGISTERS_14_28_port, QN => n3647);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1874, CK => n328, Q => 
                           REGISTERS_14_27_port, QN => n3646);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1873, CK => n331, Q => 
                           REGISTERS_14_26_port, QN => n3645);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1872, CK => n306, Q => 
                           REGISTERS_14_25_port, QN => n3644);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1871, CK => n334, Q => 
                           REGISTERS_14_24_port, QN => n3643);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1870, CK => n337, Q => 
                           REGISTERS_14_23_port, QN => n3642);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1869, CK => n340, Q => 
                           REGISTERS_14_22_port, QN => n3641);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1868, CK => n303, Q => 
                           REGISTERS_14_21_port, QN => n3640);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1867, CK => n343, Q => 
                           REGISTERS_14_20_port, QN => n3639);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1866, CK => n347, Q => 
                           REGISTERS_14_19_port, QN => n3638);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1865, CK => n350, Q => 
                           REGISTERS_14_18_port, QN => n3637);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1864, CK => n294, Q => 
                           REGISTERS_14_17_port, QN => n3636);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1863, CK => n353, Q => 
                           REGISTERS_14_16_port, QN => n3635);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1862, CK => n356, Q => 
                           REGISTERS_14_15_port, QN => n3634);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1861, CK => n359, Q => 
                           REGISTERS_14_14_port, QN => n3633);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1860, CK => n297, Q => 
                           REGISTERS_14_13_port, QN => n3632);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1859, CK => n362, Q => 
                           REGISTERS_14_12_port, QN => n3631);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1858, CK => n365, Q => 
                           REGISTERS_14_11_port, QN => n3630);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1857, CK => n368, Q => 
                           REGISTERS_14_10_port, QN => n3629);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1856, CK => n310, Q => 
                           REGISTERS_14_9_port, QN => n3628);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1855, CK => n371, Q => 
                           REGISTERS_14_8_port, QN => n3627);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1854, CK => n374, Q => 
                           REGISTERS_14_7_port, QN => n3626);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1853, CK => n377, Q => 
                           REGISTERS_14_6_port, QN => n3625);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1852, CK => n300, Q => 
                           REGISTERS_14_5_port, QN => n3624);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1851, CK => n381, Q => 
                           REGISTERS_14_4_port, QN => n3623);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1850, CK => n384, Q => 
                           REGISTERS_14_3_port, QN => n3622);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1849, CK => n387, Q => 
                           REGISTERS_14_2_port, QN => n3621);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1848, CK => n313, Q => 
                           REGISTERS_14_1_port, QN => n3620);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1847, CK => n390, Q => 
                           REGISTERS_14_0_port, QN => n3619);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1846, CK => n319, Q => 
                           REGISTERS_15_31_port, QN => n3618);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1845, CK => n322, Q => 
                           REGISTERS_15_30_port, QN => n3617);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1844, CK => n316, Q => 
                           REGISTERS_15_29_port, QN => n3616);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1843, CK => n325, Q => 
                           REGISTERS_15_28_port, QN => n3615);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1842, CK => n328, Q => 
                           REGISTERS_15_27_port, QN => n3614);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1841, CK => n331, Q => 
                           REGISTERS_15_26_port, QN => n3613);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1840, CK => n307, Q => 
                           REGISTERS_15_25_port, QN => n3612);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1839, CK => n334, Q => 
                           REGISTERS_15_24_port, QN => n3611);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1838, CK => n337, Q => 
                           REGISTERS_15_23_port, QN => n3610);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1837, CK => n340, Q => 
                           REGISTERS_15_22_port, QN => n3609);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1836, CK => n303, Q => 
                           REGISTERS_15_21_port, QN => n3608);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1835, CK => n344, Q => 
                           REGISTERS_15_20_port, QN => n3607);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1834, CK => n347, Q => 
                           REGISTERS_15_19_port, QN => n3606);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1833, CK => n350, Q => 
                           REGISTERS_15_18_port, QN => n3605);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1832, CK => n294, Q => 
                           REGISTERS_15_17_port, QN => n3604);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1831, CK => n353, Q => 
                           REGISTERS_15_16_port, QN => n3603);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1830, CK => n356, Q => 
                           REGISTERS_15_15_port, QN => n3602);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1829, CK => n359, Q => 
                           REGISTERS_15_14_port, QN => n3601);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1828, CK => n297, Q => 
                           REGISTERS_15_13_port, QN => n3600);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1827, CK => n362, Q => 
                           REGISTERS_15_12_port, QN => n3599);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1826, CK => n365, Q => 
                           REGISTERS_15_11_port, QN => n3598);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1825, CK => n368, Q => 
                           REGISTERS_15_10_port, QN => n3597);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1824, CK => n310, Q => 
                           REGISTERS_15_9_port, QN => n3596);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1823, CK => n371, Q => 
                           REGISTERS_15_8_port, QN => n3595);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1822, CK => n374, Q => 
                           REGISTERS_15_7_port, QN => n3594);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1821, CK => n378, Q => 
                           REGISTERS_15_6_port, QN => n3593);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1820, CK => n300, Q => 
                           REGISTERS_15_5_port, QN => n3592);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1819, CK => n381, Q => 
                           REGISTERS_15_4_port, QN => n3591);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1818, CK => n384, Q => 
                           REGISTERS_15_3_port, QN => n3590);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1817, CK => n387, Q => 
                           REGISTERS_15_2_port, QN => n3589);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1816, CK => n313, Q => 
                           REGISTERS_15_1_port, QN => n3588);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1815, CK => n390, Q => 
                           REGISTERS_15_0_port, QN => n3587);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1814, CK => n319, Q => 
                           REGISTERS_16_31_port, QN => n3586);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1813, CK => n322, Q => 
                           REGISTERS_16_30_port, QN => n3585);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1812, CK => n316, Q => 
                           REGISTERS_16_29_port, QN => n3584);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1811, CK => n325, Q => 
                           REGISTERS_16_28_port, QN => n3583);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1810, CK => n328, Q => 
                           REGISTERS_16_27_port, QN => n3582);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1809, CK => n331, Q => 
                           REGISTERS_16_26_port, QN => n3581);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1808, CK => n307, Q => 
                           REGISTERS_16_25_port, QN => n3580);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1807, CK => n334, Q => 
                           REGISTERS_16_24_port, QN => n3579);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1806, CK => n337, Q => 
                           REGISTERS_16_23_port, QN => n3578);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1805, CK => n341, Q => 
                           REGISTERS_16_22_port, QN => n3577);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1804, CK => n304, Q => 
                           REGISTERS_16_21_port, QN => n3576);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1803, CK => n344, Q => 
                           REGISTERS_16_20_port, QN => n3575);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1802, CK => n347, Q => 
                           REGISTERS_16_19_port, QN => n3574);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1801, CK => n350, Q => 
                           REGISTERS_16_18_port, QN => n3573);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1800, CK => n294, Q => 
                           REGISTERS_16_17_port, QN => n3572);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1799, CK => n353, Q => 
                           REGISTERS_16_16_port, QN => n3571);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1798, CK => n356, Q => 
                           REGISTERS_16_15_port, QN => n3570);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1797, CK => n359, Q => 
                           REGISTERS_16_14_port, QN => n3569);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1796, CK => n298, Q => 
                           REGISTERS_16_13_port, QN => n3568);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1795, CK => n362, Q => 
                           REGISTERS_16_12_port, QN => n3567);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1794, CK => n365, Q => 
                           REGISTERS_16_11_port, QN => n3566);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1793, CK => n368, Q => 
                           REGISTERS_16_10_port, QN => n3565);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1792, CK => n310, Q => 
                           REGISTERS_16_9_port, QN => n3564);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1791, CK => n371, Q => 
                           REGISTERS_16_8_port, QN => n3563);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1790, CK => n375, Q => 
                           REGISTERS_16_7_port, QN => n3562);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1789, CK => n378, Q => 
                           REGISTERS_16_6_port, QN => n3561);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1788, CK => n301, Q => 
                           REGISTERS_16_5_port, QN => n3560);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1787, CK => n381, Q => 
                           REGISTERS_16_4_port, QN => n3559);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1786, CK => n384, Q => 
                           REGISTERS_16_3_port, QN => n3558);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1785, CK => n387, Q => 
                           REGISTERS_16_2_port, QN => n3557);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1784, CK => n313, Q => 
                           REGISTERS_16_1_port, QN => n3556);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1783, CK => n390, Q => 
                           REGISTERS_16_0_port, QN => n3555);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1782, CK => n319, Q => 
                           REGISTERS_17_31_port, QN => n3554);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1781, CK => n322, Q => 
                           REGISTERS_17_30_port, QN => n3553);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1780, CK => n316, Q => 
                           REGISTERS_17_29_port, QN => n3552);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1779, CK => n325, Q => 
                           REGISTERS_17_28_port, QN => n3551);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1778, CK => n328, Q => 
                           REGISTERS_17_27_port, QN => n3550);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1777, CK => n331, Q => 
                           REGISTERS_17_26_port, QN => n3549);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1776, CK => n307, Q => 
                           REGISTERS_17_25_port, QN => n3548);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1775, CK => n334, Q => 
                           REGISTERS_17_24_port, QN => n3547);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1774, CK => n338, Q => 
                           REGISTERS_17_23_port, QN => n3546);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1773, CK => n341, Q => 
                           REGISTERS_17_22_port, QN => n3545);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1772, CK => n304, Q => 
                           REGISTERS_17_21_port, QN => n3544);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1771, CK => n344, Q => 
                           REGISTERS_17_20_port, QN => n3543);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1770, CK => n347, Q => 
                           REGISTERS_17_19_port, QN => n3542);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1769, CK => n350, Q => 
                           REGISTERS_17_18_port, QN => n3541);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1768, CK => n295, Q => 
                           REGISTERS_17_17_port, QN => n3540);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1767, CK => n353, Q => 
                           REGISTERS_17_16_port, QN => n3539);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1766, CK => n356, Q => 
                           REGISTERS_17_15_port, QN => n3538);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1765, CK => n359, Q => 
                           REGISTERS_17_14_port, QN => n3537);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1764, CK => n298, Q => 
                           REGISTERS_17_13_port, QN => n3536);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1763, CK => n362, Q => 
                           REGISTERS_17_12_port, QN => n3535);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1762, CK => n365, Q => 
                           REGISTERS_17_11_port, QN => n3534);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1761, CK => n368, Q => 
                           REGISTERS_17_10_port, QN => n3533);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1760, CK => n310, Q => 
                           REGISTERS_17_9_port, QN => n3532);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1759, CK => n372, Q => 
                           REGISTERS_17_8_port, QN => n3531);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1758, CK => n375, Q => 
                           REGISTERS_17_7_port, QN => n3530);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1757, CK => n378, Q => 
                           REGISTERS_17_6_port, QN => n3529);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1756, CK => n301, Q => 
                           REGISTERS_17_5_port, QN => n3528);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1755, CK => n381, Q => 
                           REGISTERS_17_4_port, QN => n3527);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1754, CK => n384, Q => 
                           REGISTERS_17_3_port, QN => n3526);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1753, CK => n387, Q => 
                           REGISTERS_17_2_port, QN => n3525);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1752, CK => n313, Q => 
                           REGISTERS_17_1_port, QN => n3524);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1751, CK => n390, Q => 
                           REGISTERS_17_0_port, QN => n3523);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1750, CK => n319, Q => 
                           REGISTERS_18_31_port, QN => n3522);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1749, CK => n322, Q => 
                           REGISTERS_18_30_port, QN => n3521);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1748, CK => n316, Q => 
                           REGISTERS_18_29_port, QN => n3520);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1747, CK => n325, Q => 
                           REGISTERS_18_28_port, QN => n3519);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1746, CK => n328, Q => 
                           REGISTERS_18_27_port, QN => n3518);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1745, CK => n331, Q => 
                           REGISTERS_18_26_port, QN => n3517);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1744, CK => n307, Q => 
                           REGISTERS_18_25_port, QN => n3516);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1743, CK => n335, Q => 
                           REGISTERS_18_24_port, QN => n3515);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1742, CK => n338, Q => 
                           REGISTERS_18_23_port, QN => n3514);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1741, CK => n341, Q => 
                           REGISTERS_18_22_port, QN => n3513);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1740, CK => n304, Q => 
                           REGISTERS_18_21_port, QN => n3512);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1739, CK => n344, Q => 
                           REGISTERS_18_20_port, QN => n3511);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1738, CK => n347, Q => 
                           REGISTERS_18_19_port, QN => n3510);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1737, CK => n350, Q => 
                           REGISTERS_18_18_port, QN => n3509);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1736, CK => n295, Q => 
                           REGISTERS_18_17_port, QN => n3508);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1735, CK => n353, Q => 
                           REGISTERS_18_16_port, QN => n3507);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1734, CK => n356, Q => 
                           REGISTERS_18_15_port, QN => n3506);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1733, CK => n359, Q => 
                           REGISTERS_18_14_port, QN => n3505);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1732, CK => n298, Q => 
                           REGISTERS_18_13_port, QN => n3504);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1731, CK => n362, Q => 
                           REGISTERS_18_12_port, QN => n3503);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1730, CK => n365, Q => 
                           REGISTERS_18_11_port, QN => n3502);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1729, CK => n369, Q => 
                           REGISTERS_18_10_port, QN => n3501);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1728, CK => n310, Q => 
                           REGISTERS_18_9_port, QN => n3500);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1727, CK => n372, Q => 
                           REGISTERS_18_8_port, QN => n3499);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1726, CK => n375, Q => 
                           REGISTERS_18_7_port, QN => n3498);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1725, CK => n378, Q => 
                           REGISTERS_18_6_port, QN => n3497);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1724, CK => n301, Q => 
                           REGISTERS_18_5_port, QN => n3496);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1723, CK => n381, Q => 
                           REGISTERS_18_4_port, QN => n3495);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1722, CK => n384, Q => 
                           REGISTERS_18_3_port, QN => n3494);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1721, CK => n387, Q => 
                           REGISTERS_18_2_port, QN => n3493);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1720, CK => n313, Q => 
                           REGISTERS_18_1_port, QN => n3492);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1719, CK => n390, Q => 
                           REGISTERS_18_0_port, QN => n3491);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1718, CK => n319, Q => 
                           REGISTERS_19_31_port, QN => n3490);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1717, CK => n322, Q => 
                           REGISTERS_19_30_port, QN => n3489);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1716, CK => n316, Q => 
                           REGISTERS_19_29_port, QN => n3488);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1715, CK => n325, Q => 
                           REGISTERS_19_28_port, QN => n3487);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1714, CK => n328, Q => 
                           REGISTERS_19_27_port, QN => n3486);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1713, CK => n332, Q => 
                           REGISTERS_19_26_port, QN => n3485);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1712, CK => n307, Q => 
                           REGISTERS_19_25_port, QN => n3484);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1711, CK => n335, Q => 
                           REGISTERS_19_24_port, QN => n3483);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1710, CK => n338, Q => 
                           REGISTERS_19_23_port, QN => n3482);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1709, CK => n341, Q => 
                           REGISTERS_19_22_port, QN => n3481);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1708, CK => n304, Q => 
                           REGISTERS_19_21_port, QN => n3480);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1707, CK => n344, Q => 
                           REGISTERS_19_20_port, QN => n3479);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1706, CK => n347, Q => 
                           REGISTERS_19_19_port, QN => n3478);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1705, CK => n350, Q => 
                           REGISTERS_19_18_port, QN => n3477);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1704, CK => n295, Q => 
                           REGISTERS_19_17_port, QN => n3476);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1703, CK => n353, Q => 
                           REGISTERS_19_16_port, QN => n3475);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1702, CK => n356, Q => 
                           REGISTERS_19_15_port, QN => n3474);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1701, CK => n359, Q => 
                           REGISTERS_19_14_port, QN => n3473);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1700, CK => n298, Q => 
                           REGISTERS_19_13_port, QN => n3472);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1699, CK => n362, Q => 
                           REGISTERS_19_12_port, QN => n3471);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1698, CK => n366, Q => 
                           REGISTERS_19_11_port, QN => n3470);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1697, CK => n369, Q => 
                           REGISTERS_19_10_port, QN => n3469);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1696, CK => n310, Q => 
                           REGISTERS_19_9_port, QN => n3468);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1695, CK => n372, Q => 
                           REGISTERS_19_8_port, QN => n3467);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1694, CK => n375, Q => 
                           REGISTERS_19_7_port, QN => n3466);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1693, CK => n378, Q => 
                           REGISTERS_19_6_port, QN => n3465);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1692, CK => n301, Q => 
                           REGISTERS_19_5_port, QN => n3464);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1691, CK => n381, Q => 
                           REGISTERS_19_4_port, QN => n3463);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1690, CK => n384, Q => 
                           REGISTERS_19_3_port, QN => n3462);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1689, CK => n387, Q => 
                           REGISTERS_19_2_port, QN => n3461);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1688, CK => n313, Q => 
                           REGISTERS_19_1_port, QN => n3460);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1687, CK => n390, Q => 
                           REGISTERS_19_0_port, QN => n3459);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1686, CK => n319, Q => 
                           REGISTERS_20_31_port, QN => n3458);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1685, CK => n322, Q => 
                           REGISTERS_20_30_port, QN => n3457);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1684, CK => n316, Q => 
                           REGISTERS_20_29_port, QN => n3456);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1683, CK => n325, Q => 
                           REGISTERS_20_28_port, QN => n3455);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1682, CK => n329, Q => 
                           REGISTERS_20_27_port, QN => n3454);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1681, CK => n332, Q => 
                           REGISTERS_20_26_port, QN => n3453);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1680, CK => n307, Q => 
                           REGISTERS_20_25_port, QN => n3452);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1679, CK => n335, Q => 
                           REGISTERS_20_24_port, QN => n3451);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1678, CK => n338, Q => 
                           REGISTERS_20_23_port, QN => n3450);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1677, CK => n341, Q => 
                           REGISTERS_20_22_port, QN => n3449);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1676, CK => n304, Q => 
                           REGISTERS_20_21_port, QN => n3448);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1675, CK => n344, Q => 
                           REGISTERS_20_20_port, QN => n3447);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1674, CK => n347, Q => 
                           REGISTERS_20_19_port, QN => n3446);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1673, CK => n350, Q => 
                           REGISTERS_20_18_port, QN => n3445);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1672, CK => n295, Q => 
                           REGISTERS_20_17_port, QN => n3444);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1671, CK => n353, Q => 
                           REGISTERS_20_16_port, QN => n3443);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1670, CK => n356, Q => 
                           REGISTERS_20_15_port, QN => n3442);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1669, CK => n359, Q => 
                           REGISTERS_20_14_port, QN => n3441);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1668, CK => n298, Q => 
                           REGISTERS_20_13_port, QN => n3440);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1667, CK => n363, Q => 
                           REGISTERS_20_12_port, QN => n3439);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1666, CK => n366, Q => 
                           REGISTERS_20_11_port, QN => n3438);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1665, CK => n369, Q => 
                           REGISTERS_20_10_port, QN => n3437);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1664, CK => n310, Q => 
                           REGISTERS_20_9_port, QN => n3436);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1663, CK => n372, Q => 
                           REGISTERS_20_8_port, QN => n3435);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1662, CK => n375, Q => 
                           REGISTERS_20_7_port, QN => n3434);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1661, CK => n378, Q => 
                           REGISTERS_20_6_port, QN => n3433);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1660, CK => n301, Q => 
                           REGISTERS_20_5_port, QN => n3432);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1659, CK => n381, Q => 
                           REGISTERS_20_4_port, QN => n3431);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1658, CK => n384, Q => 
                           REGISTERS_20_3_port, QN => n3430);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1657, CK => n387, Q => 
                           REGISTERS_20_2_port, QN => n3429);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1656, CK => n313, Q => 
                           REGISTERS_20_1_port, QN => n3428);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1655, CK => n390, Q => 
                           REGISTERS_20_0_port, QN => n3427);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1654, CK => n319, Q => 
                           REGISTERS_21_31_port, QN => n3426);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1653, CK => n322, Q => 
                           REGISTERS_21_30_port, QN => n3425);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1652, CK => n316, Q => 
                           REGISTERS_21_29_port, QN => n3424);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1651, CK => n326, Q => 
                           REGISTERS_21_28_port, QN => n3423);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1650, CK => n329, Q => 
                           REGISTERS_21_27_port, QN => n3422);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1649, CK => n332, Q => 
                           REGISTERS_21_26_port, QN => n3421);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1648, CK => n307, Q => 
                           REGISTERS_21_25_port, QN => n3420);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1647, CK => n335, Q => 
                           REGISTERS_21_24_port, QN => n3419);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1646, CK => n338, Q => 
                           REGISTERS_21_23_port, QN => n3418);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1645, CK => n341, Q => 
                           REGISTERS_21_22_port, QN => n3417);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1644, CK => n304, Q => 
                           REGISTERS_21_21_port, QN => n3416);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1643, CK => n344, Q => 
                           REGISTERS_21_20_port, QN => n3415);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1642, CK => n347, Q => 
                           REGISTERS_21_19_port, QN => n3414);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1641, CK => n350, Q => 
                           REGISTERS_21_18_port, QN => n3413);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1640, CK => n295, Q => 
                           REGISTERS_21_17_port, QN => n3412);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1639, CK => n353, Q => 
                           REGISTERS_21_16_port, QN => n3411);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1638, CK => n356, Q => 
                           REGISTERS_21_15_port, QN => n3410);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1637, CK => n360, Q => 
                           REGISTERS_21_14_port, QN => n3409);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1636, CK => n298, Q => 
                           REGISTERS_21_13_port, QN => n3408);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1635, CK => n363, Q => 
                           REGISTERS_21_12_port, QN => n3407);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1634, CK => n366, Q => 
                           REGISTERS_21_11_port, QN => n3406);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1633, CK => n369, Q => 
                           REGISTERS_21_10_port, QN => n3405);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1632, CK => n310, Q => 
                           REGISTERS_21_9_port, QN => n3404);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1631, CK => n372, Q => 
                           REGISTERS_21_8_port, QN => n3403);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1630, CK => n375, Q => 
                           REGISTERS_21_7_port, QN => n3402);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1629, CK => n378, Q => 
                           REGISTERS_21_6_port, QN => n3401);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1628, CK => n301, Q => 
                           REGISTERS_21_5_port, QN => n3400);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1627, CK => n381, Q => 
                           REGISTERS_21_4_port, QN => n3399);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1626, CK => n384, Q => 
                           REGISTERS_21_3_port, QN => n3398);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1625, CK => n387, Q => 
                           REGISTERS_21_2_port, QN => n3397);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1624, CK => n313, Q => 
                           REGISTERS_21_1_port, QN => n3396);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1623, CK => n390, Q => 
                           REGISTERS_21_0_port, QN => n3395);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1622, CK => n319, Q => 
                           REGISTERS_22_31_port, QN => n3394);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1621, CK => n323, Q => 
                           REGISTERS_22_30_port, QN => n3393);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1620, CK => n316, Q => 
                           REGISTERS_22_29_port, QN => n3392);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1619, CK => n326, Q => 
                           REGISTERS_22_28_port, QN => n3391);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1618, CK => n329, Q => 
                           REGISTERS_22_27_port, QN => n3390);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1617, CK => n332, Q => 
                           REGISTERS_22_26_port, QN => n3389);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1616, CK => n307, Q => 
                           REGISTERS_22_25_port, QN => n3388);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1615, CK => n335, Q => 
                           REGISTERS_22_24_port, QN => n3387);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1614, CK => n338, Q => 
                           REGISTERS_22_23_port, QN => n3386);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1613, CK => n341, Q => 
                           REGISTERS_22_22_port, QN => n3385);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1612, CK => n304, Q => 
                           REGISTERS_22_21_port, QN => n3384);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1611, CK => n344, Q => 
                           REGISTERS_22_20_port, QN => n3383);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1610, CK => n347, Q => 
                           REGISTERS_22_19_port, QN => n3382);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1609, CK => n350, Q => 
                           REGISTERS_22_18_port, QN => n3381);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1608, CK => n295, Q => 
                           REGISTERS_22_17_port, QN => n3380);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1607, CK => n353, Q => 
                           REGISTERS_22_16_port, QN => n3379);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1606, CK => n357, Q => 
                           REGISTERS_22_15_port, QN => n3378);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1605, CK => n360, Q => 
                           REGISTERS_22_14_port, QN => n3377);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1604, CK => n298, Q => 
                           REGISTERS_22_13_port, QN => n3376);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1603, CK => n363, Q => 
                           REGISTERS_22_12_port, QN => n3375);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1602, CK => n366, Q => 
                           REGISTERS_22_11_port, QN => n3374);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1601, CK => n369, Q => 
                           REGISTERS_22_10_port, QN => n3373);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1600, CK => n310, Q => 
                           REGISTERS_22_9_port, QN => n3372);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1599, CK => n372, Q => 
                           REGISTERS_22_8_port, QN => n3371);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1598, CK => n375, Q => 
                           REGISTERS_22_7_port, QN => n3370);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1597, CK => n378, Q => 
                           REGISTERS_22_6_port, QN => n3369);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1596, CK => n301, Q => 
                           REGISTERS_22_5_port, QN => n3368);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1595, CK => n381, Q => 
                           REGISTERS_22_4_port, QN => n3367);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1594, CK => n384, Q => 
                           REGISTERS_22_3_port, QN => n3366);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1593, CK => n387, Q => 
                           REGISTERS_22_2_port, QN => n3365);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1592, CK => n313, Q => 
                           REGISTERS_22_1_port, QN => n3364);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1591, CK => n391, Q => 
                           REGISTERS_22_0_port, QN => n3363);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1590, CK => n320, Q => 
                           REGISTERS_23_31_port, QN => n3362);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1589, CK => n323, Q => 
                           REGISTERS_23_30_port, QN => n3361);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1588, CK => n317, Q => 
                           REGISTERS_23_29_port, QN => n3360);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1587, CK => n326, Q => 
                           REGISTERS_23_28_port, QN => n3359);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1586, CK => n329, Q => 
                           REGISTERS_23_27_port, QN => n3358);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1585, CK => n332, Q => 
                           REGISTERS_23_26_port, QN => n3357);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1584, CK => n307, Q => 
                           REGISTERS_23_25_port, QN => n3356);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1583, CK => n335, Q => 
                           REGISTERS_23_24_port, QN => n3355);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1582, CK => n338, Q => 
                           REGISTERS_23_23_port, QN => n3354);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1581, CK => n341, Q => 
                           REGISTERS_23_22_port, QN => n3353);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1580, CK => n304, Q => 
                           REGISTERS_23_21_port, QN => n3352);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1579, CK => n344, Q => 
                           REGISTERS_23_20_port, QN => n3351);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1578, CK => n347, Q => 
                           REGISTERS_23_19_port, QN => n3350);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1577, CK => n350, Q => 
                           REGISTERS_23_18_port, QN => n3349);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1576, CK => n295, Q => 
                           REGISTERS_23_17_port, QN => n3348);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1575, CK => n354, Q => 
                           REGISTERS_23_16_port, QN => n3347);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1574, CK => n357, Q => 
                           REGISTERS_23_15_port, QN => n3346);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1573, CK => n360, Q => 
                           REGISTERS_23_14_port, QN => n3345);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1572, CK => n298, Q => 
                           REGISTERS_23_13_port, QN => n3344);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1571, CK => n363, Q => 
                           REGISTERS_23_12_port, QN => n3343);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1570, CK => n366, Q => 
                           REGISTERS_23_11_port, QN => n3342);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1569, CK => n369, Q => 
                           REGISTERS_23_10_port, QN => n3341);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1568, CK => n310, Q => 
                           REGISTERS_23_9_port, QN => n3340);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1567, CK => n372, Q => 
                           REGISTERS_23_8_port, QN => n3339);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1566, CK => n375, Q => 
                           REGISTERS_23_7_port, QN => n3338);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1565, CK => n378, Q => 
                           REGISTERS_23_6_port, QN => n3337);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1564, CK => n301, Q => 
                           REGISTERS_23_5_port, QN => n3336);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1563, CK => n381, Q => 
                           REGISTERS_23_4_port, QN => n3335);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1562, CK => n384, Q => 
                           REGISTERS_23_3_port, QN => n3334);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1561, CK => n388, Q => 
                           REGISTERS_23_2_port, QN => n3333);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1560, CK => n313, Q => 
                           REGISTERS_23_1_port, QN => n3332);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1559, CK => n391, Q => 
                           REGISTERS_23_0_port, QN => n3331);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1558, CK => n320, Q => 
                           REGISTERS_24_31_port, QN => n3330);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1557, CK => n323, Q => 
                           REGISTERS_24_30_port, QN => n3329);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1556, CK => n317, Q => 
                           REGISTERS_24_29_port, QN => n3328);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1555, CK => n326, Q => 
                           REGISTERS_24_28_port, QN => n3327);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1554, CK => n329, Q => 
                           REGISTERS_24_27_port, QN => n3326);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1553, CK => n332, Q => 
                           REGISTERS_24_26_port, QN => n3325);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1552, CK => n307, Q => 
                           REGISTERS_24_25_port, QN => n3324);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1551, CK => n335, Q => 
                           REGISTERS_24_24_port, QN => n3323);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1550, CK => n338, Q => 
                           REGISTERS_24_23_port, QN => n3322);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1549, CK => n341, Q => 
                           REGISTERS_24_22_port, QN => n3321);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1548, CK => n304, Q => 
                           REGISTERS_24_21_port, QN => n3320);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1547, CK => n344, Q => 
                           REGISTERS_24_20_port, QN => n3319);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1546, CK => n347, Q => 
                           REGISTERS_24_19_port, QN => n3318);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1545, CK => n351, Q => 
                           REGISTERS_24_18_port, QN => n3317);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1544, CK => n295, Q => 
                           REGISTERS_24_17_port, QN => n3316);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1543, CK => n354, Q => 
                           REGISTERS_24_16_port, QN => n3315);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1542, CK => n357, Q => 
                           REGISTERS_24_15_port, QN => n3314);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1541, CK => n360, Q => 
                           REGISTERS_24_14_port, QN => n3313);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1540, CK => n298, Q => 
                           REGISTERS_24_13_port, QN => n3312);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1539, CK => n363, Q => 
                           REGISTERS_24_12_port, QN => n3311);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1538, CK => n366, Q => 
                           REGISTERS_24_11_port, QN => n3310);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1537, CK => n369, Q => 
                           REGISTERS_24_10_port, QN => n3309);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1536, CK => n310, Q => 
                           REGISTERS_24_9_port, QN => n3308);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1535, CK => n372, Q => 
                           REGISTERS_24_8_port, QN => n3307);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1534, CK => n375, Q => 
                           REGISTERS_24_7_port, QN => n3306);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1533, CK => n378, Q => 
                           REGISTERS_24_6_port, QN => n3305);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1532, CK => n301, Q => 
                           REGISTERS_24_5_port, QN => n3304);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1531, CK => n381, Q => 
                           REGISTERS_24_4_port, QN => n3303);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1530, CK => n385, Q => 
                           REGISTERS_24_3_port, QN => n3302);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1529, CK => n388, Q => 
                           REGISTERS_24_2_port, QN => n3301);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1528, CK => n314, Q => 
                           REGISTERS_24_1_port, QN => n3300);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1527, CK => n391, Q => 
                           REGISTERS_24_0_port, QN => n3299);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1526, CK => n320, Q => 
                           REGISTERS_25_31_port, QN => n3298);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1525, CK => n323, Q => 
                           REGISTERS_25_30_port, QN => n3297);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1524, CK => n317, Q => 
                           REGISTERS_25_29_port, QN => n3296);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1523, CK => n326, Q => 
                           REGISTERS_25_28_port, QN => n3295);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1522, CK => n329, Q => 
                           REGISTERS_25_27_port, QN => n3294);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1521, CK => n332, Q => 
                           REGISTERS_25_26_port, QN => n3293);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1520, CK => n307, Q => 
                           REGISTERS_25_25_port, QN => n3292);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1519, CK => n335, Q => 
                           REGISTERS_25_24_port, QN => n3291);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1518, CK => n338, Q => 
                           REGISTERS_25_23_port, QN => n3290);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1517, CK => n341, Q => 
                           REGISTERS_25_22_port, QN => n3289);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1516, CK => n304, Q => 
                           REGISTERS_25_21_port, QN => n3288);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1515, CK => n344, Q => 
                           REGISTERS_25_20_port, QN => n3287);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1514, CK => n348, Q => 
                           REGISTERS_25_19_port, QN => n3286);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1513, CK => n351, Q => 
                           REGISTERS_25_18_port, QN => n3285);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1512, CK => n295, Q => 
                           REGISTERS_25_17_port, QN => n3284);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1511, CK => n354, Q => 
                           REGISTERS_25_16_port, QN => n3283);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1510, CK => n357, Q => 
                           REGISTERS_25_15_port, QN => n3282);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1509, CK => n360, Q => 
                           REGISTERS_25_14_port, QN => n3281);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1508, CK => n298, Q => 
                           REGISTERS_25_13_port, QN => n3280);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1507, CK => n363, Q => 
                           REGISTERS_25_12_port, QN => n3279);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1506, CK => n366, Q => 
                           REGISTERS_25_11_port, QN => n3278);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1505, CK => n369, Q => 
                           REGISTERS_25_10_port, QN => n3277);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1504, CK => n311, Q => 
                           REGISTERS_25_9_port, QN => n3276);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1503, CK => n372, Q => 
                           REGISTERS_25_8_port, QN => n3275);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1502, CK => n375, Q => 
                           REGISTERS_25_7_port, QN => n3274);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1501, CK => n378, Q => 
                           REGISTERS_25_6_port, QN => n3273);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1500, CK => n301, Q => 
                           REGISTERS_25_5_port, QN => n3272);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1499, CK => n382, Q => 
                           REGISTERS_25_4_port, QN => n3271);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1498, CK => n385, Q => 
                           REGISTERS_25_3_port, QN => n3270);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1497, CK => n388, Q => 
                           REGISTERS_25_2_port, QN => n3269);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1496, CK => n314, Q => 
                           REGISTERS_25_1_port, QN => n3268);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1495, CK => n391, Q => 
                           REGISTERS_25_0_port, QN => n3267);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1494, CK => n320, Q => 
                           REGISTERS_26_31_port, QN => n3266);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1493, CK => n323, Q => 
                           REGISTERS_26_30_port, QN => n3265);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1492, CK => n317, Q => 
                           REGISTERS_26_29_port, QN => n3264);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1491, CK => n326, Q => 
                           REGISTERS_26_28_port, QN => n3263);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1490, CK => n329, Q => 
                           REGISTERS_26_27_port, QN => n3262);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1489, CK => n332, Q => 
                           REGISTERS_26_26_port, QN => n3261);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1488, CK => n308, Q => 
                           REGISTERS_26_25_port, QN => n3260);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1487, CK => n335, Q => 
                           REGISTERS_26_24_port, QN => n3259);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1486, CK => n338, Q => 
                           REGISTERS_26_23_port, QN => n3258);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1485, CK => n341, Q => 
                           REGISTERS_26_22_port, QN => n3257);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1484, CK => n304, Q => 
                           REGISTERS_26_21_port, QN => n3256);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1483, CK => n345, Q => 
                           REGISTERS_26_20_port, QN => n3255);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1482, CK => n348, Q => 
                           REGISTERS_26_19_port, QN => n3254);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1481, CK => n351, Q => 
                           REGISTERS_26_18_port, QN => n3253);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1480, CK => n295, Q => 
                           REGISTERS_26_17_port, QN => n3252);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1479, CK => n354, Q => 
                           REGISTERS_26_16_port, QN => n3251);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1478, CK => n357, Q => 
                           REGISTERS_26_15_port, QN => n3250);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1477, CK => n360, Q => 
                           REGISTERS_26_14_port, QN => n3249);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1476, CK => n298, Q => 
                           REGISTERS_26_13_port, QN => n3248);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1475, CK => n363, Q => 
                           REGISTERS_26_12_port, QN => n3247);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1474, CK => n366, Q => 
                           REGISTERS_26_11_port, QN => n3246);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1473, CK => n369, Q => 
                           REGISTERS_26_10_port, QN => n3245);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1472, CK => n311, Q => 
                           REGISTERS_26_9_port, QN => n3244);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1471, CK => n372, Q => 
                           REGISTERS_26_8_port, QN => n3243);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1470, CK => n375, Q => 
                           REGISTERS_26_7_port, QN => n3242);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1469, CK => n379, Q => 
                           REGISTERS_26_6_port, QN => n3241);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1468, CK => n301, Q => 
                           REGISTERS_26_5_port, QN => n3240);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1467, CK => n382, Q => 
                           REGISTERS_26_4_port, QN => n3239);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1466, CK => n385, Q => 
                           REGISTERS_26_3_port, QN => n3238);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1465, CK => n388, Q => 
                           REGISTERS_26_2_port, QN => n3237);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1464, CK => n314, Q => 
                           REGISTERS_26_1_port, QN => n3236);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1463, CK => n391, Q => 
                           REGISTERS_26_0_port, QN => n3235);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1462, CK => n320, Q => 
                           REGISTERS_27_31_port, QN => n3234);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1461, CK => n323, Q => 
                           REGISTERS_27_30_port, QN => n3233);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1460, CK => n317, Q => 
                           REGISTERS_27_29_port, QN => n3232);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1459, CK => n326, Q => 
                           REGISTERS_27_28_port, QN => n3231);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1458, CK => n329, Q => 
                           REGISTERS_27_27_port, QN => n3230);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1457, CK => n332, Q => 
                           REGISTERS_27_26_port, QN => n3229);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1456, CK => n308, Q => 
                           REGISTERS_27_25_port, QN => n3228);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1455, CK => n335, Q => 
                           REGISTERS_27_24_port, QN => n3227);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1454, CK => n338, Q => 
                           REGISTERS_27_23_port, QN => n3226);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1453, CK => n342, Q => 
                           REGISTERS_27_22_port, QN => n3225);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1452, CK => n305, Q => 
                           REGISTERS_27_21_port, QN => n3224);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1451, CK => n345, Q => 
                           REGISTERS_27_20_port, QN => n3223);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1450, CK => n348, Q => 
                           REGISTERS_27_19_port, QN => n3222);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1449, CK => n351, Q => 
                           REGISTERS_27_18_port, QN => n3221);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1448, CK => n295, Q => 
                           REGISTERS_27_17_port, QN => n3220);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1447, CK => n354, Q => 
                           REGISTERS_27_16_port, QN => n3219);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1446, CK => n357, Q => 
                           REGISTERS_27_15_port, QN => n3218);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1445, CK => n360, Q => 
                           REGISTERS_27_14_port, QN => n3217);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1444, CK => n299, Q => 
                           REGISTERS_27_13_port, QN => n3216);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1443, CK => n363, Q => 
                           REGISTERS_27_12_port, QN => n3215);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1442, CK => n366, Q => 
                           REGISTERS_27_11_port, QN => n3214);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1441, CK => n369, Q => 
                           REGISTERS_27_10_port, QN => n3213);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1440, CK => n311, Q => 
                           REGISTERS_27_9_port, QN => n3212);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1439, CK => n372, Q => 
                           REGISTERS_27_8_port, QN => n3211);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1438, CK => n376, Q => 
                           REGISTERS_27_7_port, QN => n3210);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1437, CK => n379, Q => 
                           REGISTERS_27_6_port, QN => n3209);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1436, CK => n302, Q => 
                           REGISTERS_27_5_port, QN => n3208);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1435, CK => n382, Q => 
                           REGISTERS_27_4_port, QN => n3207);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1434, CK => n385, Q => 
                           REGISTERS_27_3_port, QN => n3206);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1433, CK => n388, Q => 
                           REGISTERS_27_2_port, QN => n3205);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1432, CK => n314, Q => 
                           REGISTERS_27_1_port, QN => n3204);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1431, CK => n391, Q => 
                           REGISTERS_27_0_port, QN => n3203);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1430, CK => n320, Q => 
                           REGISTERS_28_31_port, QN => n3202);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1429, CK => n323, Q => 
                           REGISTERS_28_30_port, QN => n3201);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1428, CK => n317, Q => 
                           REGISTERS_28_29_port, QN => n3200);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1427, CK => n326, Q => 
                           REGISTERS_28_28_port, QN => n3199);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1426, CK => n329, Q => 
                           REGISTERS_28_27_port, QN => n3198);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1425, CK => n332, Q => 
                           REGISTERS_28_26_port, QN => n3197);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1424, CK => n308, Q => 
                           REGISTERS_28_25_port, QN => n3196);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1423, CK => n335, Q => 
                           REGISTERS_28_24_port, QN => n3195);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1422, CK => n339, Q => 
                           REGISTERS_28_23_port, QN => n3194);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1421, CK => n342, Q => 
                           REGISTERS_28_22_port, QN => n3193);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1420, CK => n305, Q => 
                           REGISTERS_28_21_port, QN => n3192);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1419, CK => n345, Q => 
                           REGISTERS_28_20_port, QN => n3191);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1418, CK => n348, Q => 
                           REGISTERS_28_19_port, QN => n3190);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1417, CK => n351, Q => 
                           REGISTERS_28_18_port, QN => n3189);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1416, CK => n296, Q => 
                           REGISTERS_28_17_port, QN => n3188);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1415, CK => n354, Q => 
                           REGISTERS_28_16_port, QN => n3187);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1414, CK => n357, Q => 
                           REGISTERS_28_15_port, QN => n3186);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1413, CK => n360, Q => 
                           REGISTERS_28_14_port, QN => n3185);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1412, CK => n299, Q => 
                           REGISTERS_28_13_port, QN => n3184);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1411, CK => n363, Q => 
                           REGISTERS_28_12_port, QN => n3183);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1410, CK => n366, Q => 
                           REGISTERS_28_11_port, QN => n3182);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1409, CK => n369, Q => 
                           REGISTERS_28_10_port, QN => n3181);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1408, CK => n311, Q => 
                           REGISTERS_28_9_port, QN => n3180);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1407, CK => n373, Q => 
                           REGISTERS_28_8_port, QN => n3179);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1406, CK => n376, Q => 
                           REGISTERS_28_7_port, QN => n3178);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1405, CK => n379, Q => 
                           REGISTERS_28_6_port, QN => n3177);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1404, CK => n302, Q => 
                           REGISTERS_28_5_port, QN => n3176);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1403, CK => n382, Q => 
                           REGISTERS_28_4_port, QN => n3175);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1402, CK => n385, Q => 
                           REGISTERS_28_3_port, QN => n3174);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1401, CK => n388, Q => 
                           REGISTERS_28_2_port, QN => n3173);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1400, CK => n314, Q => 
                           REGISTERS_28_1_port, QN => n3172);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1399, CK => n391, Q => 
                           REGISTERS_28_0_port, QN => n3171);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1398, CK => n320, Q => 
                           REGISTERS_29_31_port, QN => n3170);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1397, CK => n323, Q => 
                           REGISTERS_29_30_port, QN => n3169);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1396, CK => n317, Q => 
                           REGISTERS_29_29_port, QN => n3168);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1395, CK => n326, Q => 
                           REGISTERS_29_28_port, QN => n3167);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1394, CK => n329, Q => 
                           REGISTERS_29_27_port, QN => n3166);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1393, CK => n332, Q => 
                           REGISTERS_29_26_port, QN => n3165);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1392, CK => n308, Q => 
                           REGISTERS_29_25_port, QN => n3164);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1391, CK => n336, Q => 
                           REGISTERS_29_24_port, QN => n3163);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1390, CK => n339, Q => 
                           REGISTERS_29_23_port, QN => n3162);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1389, CK => n342, Q => 
                           REGISTERS_29_22_port, QN => n3161);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1388, CK => n305, Q => 
                           REGISTERS_29_21_port, QN => n3160);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1387, CK => n345, Q => 
                           REGISTERS_29_20_port, QN => n3159);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1386, CK => n348, Q => 
                           REGISTERS_29_19_port, QN => n3158);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1385, CK => n351, Q => 
                           REGISTERS_29_18_port, QN => n3157);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1384, CK => n296, Q => 
                           REGISTERS_29_17_port, QN => n3156);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1383, CK => n354, Q => 
                           REGISTERS_29_16_port, QN => n3155);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1382, CK => n357, Q => 
                           REGISTERS_29_15_port, QN => n3154);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1381, CK => n360, Q => 
                           REGISTERS_29_14_port, QN => n3153);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1380, CK => n299, Q => 
                           REGISTERS_29_13_port, QN => n3152);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1379, CK => n363, Q => 
                           REGISTERS_29_12_port, QN => n3151);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1378, CK => n366, Q => 
                           REGISTERS_29_11_port, QN => n3150);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1377, CK => n370, Q => 
                           REGISTERS_29_10_port, QN => n3149);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1376, CK => n311, Q => 
                           REGISTERS_29_9_port, QN => n3148);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1375, CK => n373, Q => 
                           REGISTERS_29_8_port, QN => n3147);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1374, CK => n376, Q => 
                           REGISTERS_29_7_port, QN => n3146);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1373, CK => n379, Q => 
                           REGISTERS_29_6_port, QN => n3145);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1372, CK => n302, Q => 
                           REGISTERS_29_5_port, QN => n3144);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1371, CK => n382, Q => 
                           REGISTERS_29_4_port, QN => n3143);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1370, CK => n385, Q => 
                           REGISTERS_29_3_port, QN => n3142);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1369, CK => n388, Q => 
                           REGISTERS_29_2_port, QN => n3141);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1368, CK => n314, Q => 
                           REGISTERS_29_1_port, QN => n3140);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1367, CK => n391, Q => 
                           REGISTERS_29_0_port, QN => n3139);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1366, CK => n320, Q => 
                           REGISTERS_30_31_port, QN => n3138);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1365, CK => n323, Q => 
                           REGISTERS_30_30_port, QN => n3137);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1364, CK => n317, Q => 
                           REGISTERS_30_29_port, QN => n3136);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1363, CK => n326, Q => 
                           REGISTERS_30_28_port, QN => n3135);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1362, CK => n329, Q => 
                           REGISTERS_30_27_port, QN => n3134);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1361, CK => n333, Q => 
                           REGISTERS_30_26_port, QN => n3133);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1360, CK => n308, Q => 
                           REGISTERS_30_25_port, QN => n3132);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1359, CK => n336, Q => 
                           REGISTERS_30_24_port, QN => n3131);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1358, CK => n339, Q => 
                           REGISTERS_30_23_port, QN => n3130);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1357, CK => n342, Q => 
                           REGISTERS_30_22_port, QN => n3129);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1356, CK => n305, Q => 
                           REGISTERS_30_21_port, QN => n3128);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1355, CK => n345, Q => 
                           REGISTERS_30_20_port, QN => n3127);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1354, CK => n348, Q => 
                           REGISTERS_30_19_port, QN => n3126);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1353, CK => n351, Q => 
                           REGISTERS_30_18_port, QN => n3125);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1352, CK => n296, Q => 
                           REGISTERS_30_17_port, QN => n3124);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1351, CK => n354, Q => 
                           REGISTERS_30_16_port, QN => n3123);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1350, CK => n357, Q => 
                           REGISTERS_30_15_port, QN => n3122);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1349, CK => n360, Q => 
                           REGISTERS_30_14_port, QN => n3121);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1348, CK => n299, Q => 
                           REGISTERS_30_13_port, QN => n3120);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1347, CK => n363, Q => 
                           REGISTERS_30_12_port, QN => n3119);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1346, CK => n367, Q => 
                           REGISTERS_30_11_port, QN => n3118);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1345, CK => n370, Q => 
                           REGISTERS_30_10_port, QN => n3117);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1344, CK => n311, Q => 
                           REGISTERS_30_9_port, QN => n3116);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1343, CK => n373, Q => 
                           REGISTERS_30_8_port, QN => n3115);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1342, CK => n376, Q => 
                           REGISTERS_30_7_port, QN => n3114);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1341, CK => n379, Q => 
                           REGISTERS_30_6_port, QN => n3113);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1340, CK => n302, Q => 
                           REGISTERS_30_5_port, QN => n3112);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1339, CK => n382, Q => 
                           REGISTERS_30_4_port, QN => n3111);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1338, CK => n385, Q => 
                           REGISTERS_30_3_port, QN => n3110);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1337, CK => n388, Q => 
                           REGISTERS_30_2_port, QN => n3109);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1336, CK => n314, Q => 
                           REGISTERS_30_1_port, QN => n3108);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1335, CK => n391, Q => 
                           REGISTERS_30_0_port, QN => n3107);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1334, CK => n320, Q => 
                           REGISTERS_31_31_port, QN => n3106);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1333, CK => n323, Q => 
                           REGISTERS_31_30_port, QN => n3105);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1332, CK => n317, Q => 
                           REGISTERS_31_29_port, QN => n3104);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1331, CK => n326, Q => 
                           REGISTERS_31_28_port, QN => n3103);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1330, CK => n330, Q => 
                           REGISTERS_31_27_port, QN => n3102);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1329, CK => n333, Q => 
                           REGISTERS_31_26_port, QN => n3101);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1328, CK => n308, Q => 
                           REGISTERS_31_25_port, QN => n3100);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1327, CK => n336, Q => 
                           REGISTERS_31_24_port, QN => n3099);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1326, CK => n339, Q => 
                           REGISTERS_31_23_port, QN => n3098);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1325, CK => n342, Q => 
                           REGISTERS_31_22_port, QN => n3097);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1324, CK => n305, Q => 
                           REGISTERS_31_21_port, QN => n3096);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1323, CK => n345, Q => 
                           REGISTERS_31_20_port, QN => n3095);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1322, CK => n348, Q => 
                           REGISTERS_31_19_port, QN => n3094);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1321, CK => n351, Q => 
                           REGISTERS_31_18_port, QN => n3093);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1320, CK => n296, Q => 
                           REGISTERS_31_17_port, QN => n3092);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1319, CK => n354, Q => 
                           REGISTERS_31_16_port, QN => n3091);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1318, CK => n357, Q => 
                           REGISTERS_31_15_port, QN => n3090);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1317, CK => n360, Q => 
                           REGISTERS_31_14_port, QN => n3089);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1316, CK => n299, Q => 
                           REGISTERS_31_13_port, QN => n3088);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1315, CK => n364, Q => 
                           REGISTERS_31_12_port, QN => n3087);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1314, CK => n367, Q => 
                           REGISTERS_31_11_port, QN => n3086);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1313, CK => n370, Q => 
                           REGISTERS_31_10_port, QN => n3085);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1312, CK => n311, Q => 
                           REGISTERS_31_9_port, QN => n3084);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1311, CK => n373, Q => 
                           REGISTERS_31_8_port, QN => n3083);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1310, CK => n376, Q => 
                           REGISTERS_31_7_port, QN => n3082);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1309, CK => n379, Q => 
                           REGISTERS_31_6_port, QN => n3081);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1308, CK => n302, Q => 
                           REGISTERS_31_5_port, QN => n3080);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1307, CK => n382, Q => 
                           REGISTERS_31_4_port, QN => n3079);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1306, CK => n385, Q => 
                           REGISTERS_31_3_port, QN => n3078);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1305, CK => n388, Q => 
                           REGISTERS_31_2_port, QN => n3077);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1304, CK => n314, Q => 
                           REGISTERS_31_1_port, QN => n3076);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1303, CK => n391, Q => 
                           REGISTERS_31_0_port, QN => n3075);
   OUT1_reg_31_inst : DFF_X1 port map( D => n4162, CK => n317, Q => OUT1(31), 
                           QN => n3042);
   OUT1_reg_30_inst : DFF_X1 port map( D => n4161, CK => n320, Q => OUT1(30), 
                           QN => n3041);
   OUT1_reg_29_inst : DFF_X1 port map( D => n4160, CK => n314, Q => OUT1(29), 
                           QN => n3040);
   OUT1_reg_28_inst : DFF_X1 port map( D => n4159, CK => n324, Q => OUT1(28), 
                           QN => n3039);
   OUT1_reg_27_inst : DFF_X1 port map( D => n4158, CK => n327, Q => OUT1(27), 
                           QN => n3038);
   OUT1_reg_26_inst : DFF_X1 port map( D => n4157, CK => n330, Q => OUT1(26), 
                           QN => n3037);
   OUT1_reg_25_inst : DFF_X1 port map( D => n4156, CK => n305, Q => OUT1(25), 
                           QN => n3036);
   OUT1_reg_24_inst : DFF_X1 port map( D => n4155, CK => n333, Q => OUT1(24), 
                           QN => n3035);
   OUT1_reg_23_inst : DFF_X1 port map( D => n4154, CK => n336, Q => OUT1(23), 
                           QN => n3034);
   OUT1_reg_22_inst : DFF_X1 port map( D => n4153, CK => n339, Q => OUT1(22), 
                           QN => n3033);
   OUT1_reg_21_inst : DFF_X1 port map( D => n4152, CK => n302, Q => OUT1(21), 
                           QN => n3032);
   OUT1_reg_20_inst : DFF_X1 port map( D => n4151, CK => n342, Q => OUT1(20), 
                           QN => n3031);
   OUT1_reg_19_inst : DFF_X1 port map( D => n4150, CK => n345, Q => OUT1(19), 
                           QN => n3030);
   OUT1_reg_18_inst : DFF_X1 port map( D => n4149, CK => n348, Q => OUT1(18), 
                           QN => n3029);
   OUT1_reg_17_inst : DFF_X1 port map( D => n4148, CK => n293, Q => OUT1(17), 
                           QN => n3028);
   OUT1_reg_16_inst : DFF_X1 port map( D => n4147, CK => n351, Q => OUT1(16), 
                           QN => n3027);
   OUT1_reg_15_inst : DFF_X1 port map( D => n4146, CK => n354, Q => OUT1(15), 
                           QN => n3026);
   OUT1_reg_14_inst : DFF_X1 port map( D => n4145, CK => n358, Q => OUT1(14), 
                           QN => n3025);
   OUT1_reg_13_inst : DFF_X1 port map( D => n4144, CK => n296, Q => OUT1(13), 
                           QN => n3024);
   OUT1_reg_12_inst : DFF_X1 port map( D => n4143, CK => n361, Q => OUT1(12), 
                           QN => n3023);
   OUT1_reg_11_inst : DFF_X1 port map( D => n4142, CK => n364, Q => OUT1(11), 
                           QN => n3022);
   OUT1_reg_10_inst : DFF_X1 port map( D => n4141, CK => n367, Q => OUT1(10), 
                           QN => n3021);
   OUT1_reg_9_inst : DFF_X1 port map( D => n4140, CK => n308, Q => OUT1(9), QN 
                           => n3020);
   OUT1_reg_8_inst : DFF_X1 port map( D => n4139, CK => n370, Q => OUT1(8), QN 
                           => n3019);
   OUT1_reg_7_inst : DFF_X1 port map( D => n4138, CK => n373, Q => OUT1(7), QN 
                           => n3018);
   OUT1_reg_6_inst : DFF_X1 port map( D => n4137, CK => n376, Q => OUT1(6), QN 
                           => n3017);
   OUT1_reg_5_inst : DFF_X1 port map( D => n4136, CK => n299, Q => OUT1(5), QN 
                           => n3016);
   OUT1_reg_4_inst : DFF_X1 port map( D => n4135, CK => n379, Q => OUT1(4), QN 
                           => n3015);
   OUT1_reg_3_inst : DFF_X1 port map( D => n4134, CK => n382, Q => OUT1(3), QN 
                           => n3014);
   OUT1_reg_2_inst : DFF_X1 port map( D => n4133, CK => n385, Q => OUT1(2), QN 
                           => n3013);
   OUT1_reg_1_inst : DFF_X1 port map( D => n4132, CK => n311, Q => OUT1(1), QN 
                           => n3012);
   OUT1_reg_0_inst : DFF_X1 port map( D => n4131, CK => n388, Q => OUT1(0), QN 
                           => n3011);
   U3 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n437, ZN => n1);
   U4 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => n1121, ZN => n2);
   U5 : AND2_X1 port map( A1 => n437, A2 => n1119, ZN => n3);
   U6 : AND2_X1 port map( A1 => n1121, A2 => n2827, ZN => n4);
   U7 : AND2_X1 port map( A1 => n436, A2 => ADD_RD1(0), ZN => n5);
   U8 : AND2_X1 port map( A1 => n439, A2 => ADD_RD1(0), ZN => n6);
   U9 : AND2_X1 port map( A1 => n438, A2 => ADD_RD1(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n436, A2 => n1119, ZN => n8);
   U11 : AND2_X1 port map( A1 => n439, A2 => n1119, ZN => n9);
   U12 : AND2_X1 port map( A1 => n438, A2 => n1119, ZN => n10);
   U13 : AND2_X1 port map( A1 => n1120, A2 => ADD_RD2(0), ZN => n11);
   U14 : AND2_X1 port map( A1 => n1123, A2 => ADD_RD2(0), ZN => n12);
   U15 : AND2_X1 port map( A1 => n1122, A2 => ADD_RD2(0), ZN => n13);
   U16 : AND2_X1 port map( A1 => n1120, A2 => n2827, ZN => n14);
   U17 : AND2_X1 port map( A1 => n1123, A2 => n2827, ZN => n15);
   U18 : AND2_X1 port map( A1 => n1122, A2 => n2827, ZN => n16);
   U19 : NAND2_X2 port map( A1 => n2940, A2 => n291, ZN => n2941);
   U20 : NAND2_X2 port map( A1 => n2943, A2 => n291, ZN => n2944);
   U21 : NAND2_X2 port map( A1 => n2949, A2 => n291, ZN => n2950);
   U22 : NAND2_X2 port map( A1 => n2934, A2 => n291, ZN => n2935);
   U23 : NAND2_X2 port map( A1 => n2937, A2 => n291, ZN => n2938);
   U24 : NAND2_X2 port map( A1 => n2952, A2 => n291, ZN => n2953);
   U25 : NAND2_X2 port map( A1 => n2958, A2 => n290, ZN => n2959);
   U26 : NAND2_X2 port map( A1 => n2961, A2 => n290, ZN => n2962);
   U27 : NAND2_X2 port map( A1 => n2963, A2 => n290, ZN => n2964);
   U28 : NAND2_X2 port map( A1 => n2965, A2 => n290, ZN => n2966);
   U29 : NAND2_X2 port map( A1 => n2971, A2 => n290, ZN => n2972);
   U30 : NAND2_X2 port map( A1 => n2973, A2 => n290, ZN => n2974);
   U31 : NAND2_X2 port map( A1 => n2975, A2 => n290, ZN => n2976);
   U32 : NAND2_X2 port map( A1 => n2978, A2 => n290, ZN => n2979);
   U33 : NAND2_X2 port map( A1 => n2980, A2 => n290, ZN => n2981);
   U34 : NAND2_X2 port map( A1 => n2982, A2 => n290, ZN => n2983);
   U35 : NAND2_X2 port map( A1 => n2984, A2 => n289, ZN => n2985);
   U36 : NAND2_X2 port map( A1 => n2986, A2 => n289, ZN => n2987);
   U37 : NAND2_X2 port map( A1 => n2988, A2 => n289, ZN => n2989);
   U38 : NAND2_X2 port map( A1 => n2990, A2 => n289, ZN => n2991);
   U39 : NAND2_X2 port map( A1 => n2992, A2 => n289, ZN => n2993);
   U40 : NAND2_X2 port map( A1 => n2942, A2 => n2933, ZN => n2940);
   U41 : NAND2_X2 port map( A1 => n2960, A2 => n2939, ZN => n2963);
   U42 : NAND2_X2 port map( A1 => n2977, A2 => n2936, ZN => n2978);
   U43 : NAND2_X2 port map( A1 => n2994, A2 => n2932, ZN => n2992);
   U44 : NAND2_X2 port map( A1 => n2995, A2 => n289, ZN => n2996);
   U45 : NAND2_X2 port map( A1 => n2939, A2 => n2933, ZN => n2937);
   U46 : NAND2_X2 port map( A1 => n2960, A2 => n2942, ZN => n2965);
   U47 : NAND2_X2 port map( A1 => n2977, A2 => n2932, ZN => n2975);
   U48 : NAND2_X2 port map( A1 => n2994, A2 => n2936, ZN => n2995);
   U49 : NAND2_X2 port map( A1 => n2998, A2 => n289, ZN => n2999);
   U50 : NAND2_X2 port map( A1 => n2936, A2 => n2933, ZN => n2934);
   U51 : NAND2_X2 port map( A1 => n2960, A2 => n2932, ZN => n2958);
   U52 : NAND2_X2 port map( A1 => n2977, A2 => n2942, ZN => n2982);
   U53 : NAND2_X2 port map( A1 => n2994, A2 => n2939, ZN => n2998);
   U54 : NAND2_X2 port map( A1 => n3001, A2 => n289, ZN => n3002);
   U55 : NAND2_X2 port map( A1 => n2945, A2 => n2933, ZN => n2943);
   U56 : NAND2_X2 port map( A1 => n2960, A2 => n2936, ZN => n2961);
   U57 : NAND2_X2 port map( A1 => n2977, A2 => n2939, ZN => n2980);
   U58 : NAND2_X2 port map( A1 => n2994, A2 => n2942, ZN => n3001);
   U59 : NAND2_X2 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n2820);
   U60 : NAND2_X2 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n1112);
   U61 : NAND2_X2 port map( A1 => n2862, A2 => n291, ZN => n2828);
   U62 : NAND2_X2 port map( A1 => n3003, A2 => n289, ZN => n3004);
   U63 : NAND2_X2 port map( A1 => n2954, A2 => n2933, ZN => n2952);
   U64 : NAND2_X2 port map( A1 => n2960, A2 => n2951, ZN => n2971);
   U65 : NAND2_X2 port map( A1 => n2977, A2 => n2948, ZN => n2986);
   U66 : NAND2_X2 port map( A1 => n2994, A2 => n2945, ZN => n3003);
   U67 : NAND2_X2 port map( A1 => n2897, A2 => n291, ZN => n2863);
   U68 : NAND2_X2 port map( A1 => n3005, A2 => n289, ZN => n3006);
   U69 : NAND2_X2 port map( A1 => ADD_RD2(4), A2 => n2824, ZN => n2822);
   U70 : NAND2_X2 port map( A1 => ADD_RD1(4), A2 => n1116, ZN => n1114);
   U71 : NAND2_X2 port map( A1 => n2951, A2 => n2933, ZN => n2949);
   U72 : NAND2_X2 port map( A1 => n2960, A2 => n2954, ZN => n2973);
   U73 : NAND2_X2 port map( A1 => n2977, A2 => n2945, ZN => n2984);
   U74 : NAND2_X2 port map( A1 => n2994, A2 => n2948, ZN => n3005);
   U75 : NAND2_X2 port map( A1 => n2946, A2 => n291, ZN => n2947);
   U76 : NAND2_X2 port map( A1 => n2967, A2 => n290, ZN => n2968);
   U77 : NAND2_X2 port map( A1 => n3007, A2 => n289, ZN => n3008);
   U78 : NAND2_X2 port map( A1 => n2948, A2 => n2933, ZN => n2946);
   U79 : NAND2_X2 port map( A1 => n2960, A2 => n2945, ZN => n2967);
   U80 : NAND2_X2 port map( A1 => n2977, A2 => n2954, ZN => n2990);
   U81 : NAND2_X2 port map( A1 => n2994, A2 => n2951, ZN => n3007);
   U82 : NOR2_X4 port map( A1 => n2824, A2 => ADD_RD2(4), ZN => n2816);
   U83 : NOR2_X4 port map( A1 => n1116, A2 => ADD_RD1(4), ZN => n1108);
   U84 : NAND2_X2 port map( A1 => n2898, A2 => n291, ZN => n2900);
   U85 : NAND2_X2 port map( A1 => n2969, A2 => n290, ZN => n2970);
   U86 : NAND2_X2 port map( A1 => n3009, A2 => n289, ZN => n3010);
   U87 : INV_X2 port map( A => n2862, ZN => n2830);
   U88 : INV_X2 port map( A => n2897, ZN => n2865);
   U89 : INV_X2 port map( A => DATAIN(31), ZN => n2899);
   U90 : INV_X2 port map( A => DATAIN(30), ZN => n2901);
   U91 : INV_X2 port map( A => DATAIN(29), ZN => n2902);
   U92 : INV_X2 port map( A => DATAIN(28), ZN => n2903);
   U93 : INV_X2 port map( A => DATAIN(27), ZN => n2904);
   U94 : INV_X2 port map( A => DATAIN(26), ZN => n2905);
   U95 : INV_X2 port map( A => DATAIN(25), ZN => n2906);
   U96 : INV_X2 port map( A => DATAIN(24), ZN => n2907);
   U97 : INV_X2 port map( A => DATAIN(23), ZN => n2908);
   U98 : INV_X2 port map( A => DATAIN(22), ZN => n2909);
   U99 : INV_X2 port map( A => DATAIN(21), ZN => n2910);
   U100 : INV_X2 port map( A => DATAIN(20), ZN => n2911);
   U101 : INV_X2 port map( A => DATAIN(19), ZN => n2912);
   U102 : INV_X2 port map( A => DATAIN(18), ZN => n2913);
   U103 : INV_X2 port map( A => DATAIN(17), ZN => n2914);
   U104 : INV_X2 port map( A => DATAIN(16), ZN => n2915);
   U105 : INV_X2 port map( A => DATAIN(15), ZN => n2916);
   U106 : INV_X2 port map( A => DATAIN(14), ZN => n2917);
   U107 : INV_X2 port map( A => DATAIN(13), ZN => n2918);
   U108 : INV_X2 port map( A => DATAIN(12), ZN => n2919);
   U109 : INV_X2 port map( A => DATAIN(11), ZN => n2920);
   U110 : INV_X2 port map( A => DATAIN(10), ZN => n2921);
   U111 : INV_X2 port map( A => DATAIN(9), ZN => n2922);
   U112 : INV_X2 port map( A => DATAIN(8), ZN => n2923);
   U113 : INV_X2 port map( A => DATAIN(7), ZN => n2924);
   U114 : INV_X2 port map( A => DATAIN(6), ZN => n2925);
   U115 : INV_X2 port map( A => DATAIN(5), ZN => n2926);
   U116 : INV_X2 port map( A => DATAIN(4), ZN => n2927);
   U117 : INV_X2 port map( A => DATAIN(3), ZN => n2928);
   U118 : INV_X2 port map( A => DATAIN(2), ZN => n2929);
   U119 : INV_X2 port map( A => DATAIN(1), ZN => n2930);
   U120 : INV_X2 port map( A => DATAIN(0), ZN => n2931);
   U121 : NAND2_X2 port map( A1 => n2960, A2 => n2948, ZN => n2969);
   U122 : NAND2_X2 port map( A1 => n2977, A2 => n2951, ZN => n2988);
   U123 : NAND2_X2 port map( A1 => n2994, A2 => n2954, ZN => n3009);
   U124 : NAND2_X2 port map( A1 => n2932, A2 => n2933, ZN => n2898);
   U125 : NOR2_X4 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n2818);
   U126 : NOR2_X4 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n1110);
   U127 : BUF_X1 port map( A => n432, Z => n430);
   U128 : BUF_X1 port map( A => n432, Z => n429);
   U129 : BUF_X1 port map( A => n433, Z => n428);
   U130 : BUF_X1 port map( A => n433, Z => n427);
   U131 : BUF_X1 port map( A => n433, Z => n426);
   U132 : BUF_X1 port map( A => n434, Z => n425);
   U133 : BUF_X1 port map( A => n435, Z => n433);
   U134 : BUF_X1 port map( A => n435, Z => n432);
   U135 : BUF_X1 port map( A => n151_port, Z => n149_port);
   U136 : BUF_X1 port map( A => n134_port, Z => n132_port);
   U137 : BUF_X1 port map( A => n151_port, Z => n148_port);
   U138 : BUF_X1 port map( A => n134_port, Z => n131_port);
   U139 : BUF_X1 port map( A => n287, Z => n285);
   U140 : BUF_X1 port map( A => n270, Z => n268);
   U141 : BUF_X1 port map( A => n287, Z => n284);
   U142 : BUF_X1 port map( A => n270, Z => n267);
   U143 : BUF_X1 port map( A => n117, Z => n115);
   U144 : BUF_X1 port map( A => n100, Z => n98);
   U145 : BUF_X1 port map( A => n117, Z => n114);
   U146 : BUF_X1 port map( A => n100, Z => n97);
   U147 : BUF_X1 port map( A => n253, Z => n251);
   U148 : BUF_X1 port map( A => n236, Z => n234);
   U149 : BUF_X1 port map( A => n253, Z => n250);
   U150 : BUF_X1 port map( A => n236, Z => n233);
   U151 : BUF_X1 port map( A => CLK, Z => n435);
   U152 : BUF_X1 port map( A => n10, Z => n151_port);
   U153 : BUF_X1 port map( A => n9, Z => n134_port);
   U154 : BUF_X1 port map( A => n16, Z => n287);
   U155 : BUF_X1 port map( A => n15, Z => n270);
   U156 : BUF_X1 port map( A => n8, Z => n117);
   U157 : BUF_X1 port map( A => n3, Z => n100);
   U158 : BUF_X1 port map( A => n14, Z => n253);
   U159 : BUF_X1 port map( A => n4, Z => n236);
   U160 : BUF_X1 port map( A => n83_port, Z => n81_port);
   U161 : BUF_X1 port map( A => n66_port, Z => n64_port);
   U162 : BUF_X1 port map( A => n49, Z => n47);
   U163 : BUF_X1 port map( A => n32, Z => n30);
   U164 : BUF_X1 port map( A => n83_port, Z => n80_port);
   U165 : BUF_X1 port map( A => n66_port, Z => n63_port);
   U166 : BUF_X1 port map( A => n49, Z => n46);
   U167 : BUF_X1 port map( A => n32, Z => n29);
   U168 : BUF_X1 port map( A => n219, Z => n217);
   U169 : BUF_X1 port map( A => n202, Z => n200);
   U170 : BUF_X1 port map( A => n185, Z => n183);
   U171 : BUF_X1 port map( A => n168, Z => n166);
   U172 : BUF_X1 port map( A => n219, Z => n216);
   U173 : BUF_X1 port map( A => n202, Z => n199);
   U174 : BUF_X1 port map( A => n185, Z => n182);
   U175 : BUF_X1 port map( A => n168, Z => n165);
   U176 : BUF_X1 port map( A => n152_port, Z => n147_port);
   U177 : BUF_X1 port map( A => n135_port, Z => n130_port);
   U178 : BUF_X1 port map( A => n288, Z => n283);
   U179 : BUF_X1 port map( A => n271, Z => n266);
   U180 : BUF_X1 port map( A => n118, Z => n113);
   U181 : BUF_X1 port map( A => n101, Z => n96);
   U182 : BUF_X1 port map( A => n254, Z => n249);
   U183 : BUF_X1 port map( A => n237, Z => n232);
   U184 : BUF_X1 port map( A => n7, Z => n83_port);
   U185 : BUF_X1 port map( A => n6, Z => n66_port);
   U186 : BUF_X1 port map( A => n5, Z => n49);
   U187 : BUF_X1 port map( A => n1, Z => n32);
   U188 : BUF_X1 port map( A => n13, Z => n219);
   U189 : BUF_X1 port map( A => n12, Z => n202);
   U190 : BUF_X1 port map( A => n11, Z => n185);
   U191 : BUF_X1 port map( A => n2, Z => n168);
   U192 : BUF_X1 port map( A => n84_port, Z => n79_port);
   U193 : BUF_X1 port map( A => n67_port, Z => n62_port);
   U194 : BUF_X1 port map( A => n50, Z => n45);
   U195 : BUF_X1 port map( A => n33, Z => n28);
   U196 : BUF_X1 port map( A => n220, Z => n215);
   U197 : BUF_X1 port map( A => n203, Z => n198);
   U198 : BUF_X1 port map( A => n186, Z => n181);
   U199 : BUF_X1 port map( A => n169, Z => n164);
   U200 : BUF_X1 port map( A => n402, Z => n360);
   U201 : BUF_X1 port map( A => n413, Z => n326);
   U202 : BUF_X1 port map( A => n401, Z => n363);
   U203 : BUF_X1 port map( A => n412, Z => n329);
   U204 : BUF_X1 port map( A => n400, Z => n366);
   U205 : BUF_X1 port map( A => n411, Z => n332);
   U206 : BUF_X1 port map( A => n399, Z => n369);
   U207 : BUF_X1 port map( A => n410, Z => n335);
   U208 : BUF_X1 port map( A => n398, Z => n372);
   U209 : BUF_X1 port map( A => n409, Z => n338);
   U210 : BUF_X1 port map( A => n397, Z => n375);
   U211 : BUF_X1 port map( A => n408, Z => n341);
   U212 : BUF_X1 port map( A => n396, Z => n378);
   U213 : BUF_X1 port map( A => n407, Z => n344);
   U214 : BUF_X1 port map( A => n395, Z => n381);
   U215 : BUF_X1 port map( A => n419, Z => n310);
   U216 : BUF_X1 port map( A => n406, Z => n347);
   U217 : BUF_X1 port map( A => n418, Z => n313);
   U218 : BUF_X1 port map( A => n394, Z => n384);
   U219 : BUF_X1 port map( A => n405, Z => n350);
   U220 : BUF_X1 port map( A => n393, Z => n387);
   U221 : BUF_X1 port map( A => n404, Z => n353);
   U222 : BUF_X1 port map( A => n417, Z => n316);
   U223 : BUF_X1 port map( A => n416, Z => n319);
   U224 : BUF_X1 port map( A => n392, Z => n390);
   U225 : BUF_X1 port map( A => n403, Z => n356);
   U226 : BUF_X1 port map( A => n415, Z => n322);
   U227 : BUF_X1 port map( A => n402, Z => n359);
   U228 : BUF_X1 port map( A => n414, Z => n325);
   U229 : BUF_X1 port map( A => n401, Z => n362);
   U230 : BUF_X1 port map( A => n413, Z => n328);
   U231 : BUF_X1 port map( A => n400, Z => n365);
   U232 : BUF_X1 port map( A => n412, Z => n331);
   U233 : BUF_X1 port map( A => n399, Z => n368);
   U234 : BUF_X1 port map( A => n411, Z => n334);
   U235 : BUF_X1 port map( A => n398, Z => n371);
   U236 : BUF_X1 port map( A => n410, Z => n337);
   U237 : BUF_X1 port map( A => n397, Z => n374);
   U238 : BUF_X1 port map( A => n409, Z => n340);
   U239 : BUF_X1 port map( A => n396, Z => n377);
   U240 : BUF_X1 port map( A => n408, Z => n343);
   U241 : BUF_X1 port map( A => n395, Z => n380);
   U242 : BUF_X1 port map( A => n419, Z => n309);
   U243 : BUF_X1 port map( A => n407, Z => n346);
   U244 : BUF_X1 port map( A => n418, Z => n312);
   U245 : BUF_X1 port map( A => n394, Z => n383);
   U246 : BUF_X1 port map( A => n406, Z => n349);
   U247 : BUF_X1 port map( A => n393, Z => n386);
   U248 : BUF_X1 port map( A => n405, Z => n352);
   U249 : BUF_X1 port map( A => n417, Z => n315);
   U250 : BUF_X1 port map( A => n416, Z => n318);
   U251 : BUF_X1 port map( A => n392, Z => n389);
   U252 : BUF_X1 port map( A => n403, Z => n358);
   U253 : BUF_X1 port map( A => n404, Z => n355);
   U254 : BUF_X1 port map( A => n414, Z => n324);
   U255 : BUF_X1 port map( A => n415, Z => n321);
   U256 : BUF_X1 port map( A => n416, Z => n317);
   U257 : BUF_X1 port map( A => n393, Z => n388);
   U258 : BUF_X1 port map( A => n418, Z => n311);
   U259 : BUF_X1 port map( A => n394, Z => n385);
   U260 : BUF_X1 port map( A => n395, Z => n382);
   U261 : BUF_X1 port map( A => n396, Z => n379);
   U262 : BUF_X1 port map( A => n397, Z => n376);
   U263 : BUF_X1 port map( A => n398, Z => n373);
   U264 : BUF_X1 port map( A => n399, Z => n370);
   U265 : BUF_X1 port map( A => n419, Z => n308);
   U266 : BUF_X1 port map( A => n400, Z => n367);
   U267 : BUF_X1 port map( A => n401, Z => n364);
   U268 : BUF_X1 port map( A => n402, Z => n361);
   U269 : BUF_X1 port map( A => n403, Z => n357);
   U270 : BUF_X1 port map( A => n404, Z => n354);
   U271 : BUF_X1 port map( A => n405, Z => n351);
   U272 : BUF_X1 port map( A => n406, Z => n348);
   U273 : BUF_X1 port map( A => n407, Z => n345);
   U274 : BUF_X1 port map( A => n408, Z => n342);
   U275 : BUF_X1 port map( A => n409, Z => n339);
   U276 : BUF_X1 port map( A => n410, Z => n336);
   U277 : BUF_X1 port map( A => n411, Z => n333);
   U278 : BUF_X1 port map( A => n412, Z => n330);
   U279 : BUF_X1 port map( A => n413, Z => n327);
   U280 : BUF_X1 port map( A => n414, Z => n323);
   U281 : BUF_X1 port map( A => n417, Z => n314);
   U282 : BUF_X1 port map( A => n415, Z => n320);
   U283 : BUF_X1 port map( A => n392, Z => n391);
   U284 : BUF_X1 port map( A => n426, Z => n416);
   U285 : BUF_X1 port map( A => n426, Z => n418);
   U286 : BUF_X1 port map( A => n430, Z => n395);
   U287 : BUF_X1 port map( A => n430, Z => n396);
   U288 : BUF_X1 port map( A => n430, Z => n397);
   U289 : BUF_X1 port map( A => n430, Z => n398);
   U290 : BUF_X1 port map( A => n430, Z => n399);
   U291 : BUF_X1 port map( A => n426, Z => n419);
   U292 : BUF_X1 port map( A => n429, Z => n400);
   U293 : BUF_X1 port map( A => n429, Z => n401);
   U294 : BUF_X1 port map( A => n429, Z => n402);
   U295 : BUF_X1 port map( A => n429, Z => n403);
   U296 : BUF_X1 port map( A => n429, Z => n404);
   U297 : BUF_X1 port map( A => n428, Z => n405);
   U298 : BUF_X1 port map( A => n428, Z => n406);
   U299 : BUF_X1 port map( A => n428, Z => n407);
   U300 : BUF_X1 port map( A => n428, Z => n408);
   U301 : BUF_X1 port map( A => n428, Z => n409);
   U302 : BUF_X1 port map( A => n427, Z => n410);
   U303 : BUF_X1 port map( A => n427, Z => n411);
   U304 : BUF_X1 port map( A => n427, Z => n412);
   U305 : BUF_X1 port map( A => n427, Z => n413);
   U306 : BUF_X1 port map( A => n427, Z => n414);
   U307 : BUF_X1 port map( A => n426, Z => n417);
   U308 : BUF_X1 port map( A => n426, Z => n415);
   U309 : BUF_X1 port map( A => n431, Z => n392);
   U310 : BUF_X1 port map( A => n431, Z => n393);
   U311 : BUF_X1 port map( A => n431, Z => n394);
   U312 : BUF_X1 port map( A => n424, Z => n295);
   U313 : BUF_X1 port map( A => n422, Z => n301);
   U314 : BUF_X1 port map( A => n423, Z => n298);
   U315 : BUF_X1 port map( A => n421, Z => n304);
   U316 : BUF_X1 port map( A => n420, Z => n307);
   U317 : BUF_X1 port map( A => n424, Z => n294);
   U318 : BUF_X1 port map( A => n422, Z => n300);
   U319 : BUF_X1 port map( A => n423, Z => n297);
   U320 : BUF_X1 port map( A => n421, Z => n303);
   U321 : BUF_X1 port map( A => n420, Z => n306);
   U322 : BUF_X1 port map( A => n422, Z => n299);
   U323 : BUF_X1 port map( A => n421, Z => n302);
   U324 : BUF_X1 port map( A => n423, Z => n296);
   U325 : BUF_X1 port map( A => n420, Z => n305);
   U326 : BUF_X1 port map( A => n424, Z => n293);
   U327 : BUF_X1 port map( A => n425, Z => n422);
   U328 : BUF_X1 port map( A => n425, Z => n421);
   U329 : BUF_X1 port map( A => n425, Z => n423);
   U330 : BUF_X1 port map( A => n425, Z => n420);
   U331 : BUF_X1 port map( A => n425, Z => n424);
   U332 : BUF_X1 port map( A => n432, Z => n431);
   U333 : BUF_X1 port map( A => n149_port, Z => n138_port);
   U334 : BUF_X1 port map( A => n149_port, Z => n139_port);
   U335 : BUF_X1 port map( A => n149_port, Z => n140_port);
   U336 : BUF_X1 port map( A => n148_port, Z => n141_port);
   U337 : BUF_X1 port map( A => n148_port, Z => n142_port);
   U338 : BUF_X1 port map( A => n148_port, Z => n143_port);
   U339 : BUF_X1 port map( A => n285, Z => n274);
   U340 : BUF_X1 port map( A => n285, Z => n275);
   U341 : BUF_X1 port map( A => n285, Z => n276);
   U342 : BUF_X1 port map( A => n284, Z => n277);
   U343 : BUF_X1 port map( A => n284, Z => n278);
   U344 : BUF_X1 port map( A => n284, Z => n279);
   U345 : BUF_X1 port map( A => n115, Z => n104);
   U346 : BUF_X1 port map( A => n115, Z => n105);
   U347 : BUF_X1 port map( A => n115, Z => n106);
   U348 : BUF_X1 port map( A => n114, Z => n107);
   U349 : BUF_X1 port map( A => n114, Z => n108);
   U350 : BUF_X1 port map( A => n114, Z => n109);
   U351 : BUF_X1 port map( A => n251, Z => n240);
   U352 : BUF_X1 port map( A => n251, Z => n241);
   U353 : BUF_X1 port map( A => n251, Z => n242);
   U354 : BUF_X1 port map( A => n250, Z => n243);
   U355 : BUF_X1 port map( A => n250, Z => n244);
   U356 : BUF_X1 port map( A => n250, Z => n245);
   U357 : BUF_X1 port map( A => n150_port, Z => n136_port);
   U358 : BUF_X1 port map( A => n150_port, Z => n137_port);
   U359 : BUF_X1 port map( A => n286, Z => n272);
   U360 : BUF_X1 port map( A => n286, Z => n273);
   U361 : BUF_X1 port map( A => n116, Z => n102);
   U362 : BUF_X1 port map( A => n116, Z => n103);
   U363 : BUF_X1 port map( A => n252, Z => n238);
   U364 : BUF_X1 port map( A => n252, Z => n239);
   U365 : BUF_X1 port map( A => n132_port, Z => n121);
   U366 : BUF_X1 port map( A => n132_port, Z => n122);
   U367 : BUF_X1 port map( A => n132_port, Z => n123);
   U368 : BUF_X1 port map( A => n131_port, Z => n124);
   U369 : BUF_X1 port map( A => n131_port, Z => n125);
   U370 : BUF_X1 port map( A => n131_port, Z => n126);
   U371 : BUF_X1 port map( A => n268, Z => n257);
   U372 : BUF_X1 port map( A => n268, Z => n258);
   U373 : BUF_X1 port map( A => n268, Z => n259);
   U374 : BUF_X1 port map( A => n267, Z => n260);
   U375 : BUF_X1 port map( A => n267, Z => n261);
   U376 : BUF_X1 port map( A => n267, Z => n262);
   U377 : BUF_X1 port map( A => n98, Z => n87_port);
   U378 : BUF_X1 port map( A => n98, Z => n88_port);
   U379 : BUF_X1 port map( A => n98, Z => n89_port);
   U380 : BUF_X1 port map( A => n97, Z => n90_port);
   U381 : BUF_X1 port map( A => n97, Z => n91_port);
   U382 : BUF_X1 port map( A => n97, Z => n92);
   U383 : BUF_X1 port map( A => n234, Z => n223);
   U384 : BUF_X1 port map( A => n234, Z => n224);
   U385 : BUF_X1 port map( A => n234, Z => n225);
   U386 : BUF_X1 port map( A => n233, Z => n226);
   U387 : BUF_X1 port map( A => n233, Z => n227);
   U388 : BUF_X1 port map( A => n233, Z => n228);
   U389 : BUF_X1 port map( A => n133_port, Z => n119);
   U390 : BUF_X1 port map( A => n133_port, Z => n120);
   U391 : BUF_X1 port map( A => n269, Z => n255);
   U392 : BUF_X1 port map( A => n269, Z => n256);
   U393 : BUF_X1 port map( A => n99, Z => n85_port);
   U394 : BUF_X1 port map( A => n99, Z => n86_port);
   U395 : BUF_X1 port map( A => n235, Z => n221);
   U396 : BUF_X1 port map( A => n235, Z => n222);
   U397 : BUF_X1 port map( A => n435, Z => n434);
   U398 : BUF_X1 port map( A => n151_port, Z => n150_port);
   U399 : BUF_X1 port map( A => n134_port, Z => n133_port);
   U400 : BUF_X1 port map( A => n287, Z => n286);
   U401 : BUF_X1 port map( A => n270, Z => n269);
   U402 : BUF_X1 port map( A => n117, Z => n116);
   U403 : BUF_X1 port map( A => n100, Z => n99);
   U404 : BUF_X1 port map( A => n253, Z => n252);
   U405 : BUF_X1 port map( A => n236, Z => n235);
   U406 : BUF_X1 port map( A => n81_port, Z => n70_port);
   U407 : BUF_X1 port map( A => n47, Z => n36);
   U408 : BUF_X1 port map( A => n81_port, Z => n71_port);
   U409 : BUF_X1 port map( A => n47, Z => n37);
   U410 : BUF_X1 port map( A => n81_port, Z => n72_port);
   U411 : BUF_X1 port map( A => n47, Z => n38);
   U412 : BUF_X1 port map( A => n80_port, Z => n73_port);
   U413 : BUF_X1 port map( A => n46, Z => n39);
   U414 : BUF_X1 port map( A => n80_port, Z => n74_port);
   U415 : BUF_X1 port map( A => n46, Z => n40);
   U416 : BUF_X1 port map( A => n80_port, Z => n75_port);
   U417 : BUF_X1 port map( A => n46, Z => n41);
   U418 : BUF_X1 port map( A => n217, Z => n206);
   U419 : BUF_X1 port map( A => n183, Z => n172);
   U420 : BUF_X1 port map( A => n217, Z => n207);
   U421 : BUF_X1 port map( A => n183, Z => n173);
   U422 : BUF_X1 port map( A => n217, Z => n208);
   U423 : BUF_X1 port map( A => n183, Z => n174);
   U424 : BUF_X1 port map( A => n216, Z => n209);
   U425 : BUF_X1 port map( A => n182, Z => n175);
   U426 : BUF_X1 port map( A => n216, Z => n210);
   U427 : BUF_X1 port map( A => n182, Z => n176);
   U428 : BUF_X1 port map( A => n216, Z => n211);
   U429 : BUF_X1 port map( A => n182, Z => n177);
   U430 : BUF_X1 port map( A => n147_port, Z => n144_port);
   U431 : BUF_X1 port map( A => n147_port, Z => n145_port);
   U432 : BUF_X1 port map( A => n283, Z => n280);
   U433 : BUF_X1 port map( A => n283, Z => n281);
   U434 : BUF_X1 port map( A => n113, Z => n110);
   U435 : BUF_X1 port map( A => n113, Z => n111);
   U436 : BUF_X1 port map( A => n249, Z => n246);
   U437 : BUF_X1 port map( A => n249, Z => n247);
   U438 : BUF_X1 port map( A => n292, Z => n289);
   U439 : BUF_X1 port map( A => n292, Z => n290);
   U440 : BUF_X1 port map( A => n82_port, Z => n68_port);
   U441 : BUF_X1 port map( A => n48, Z => n34);
   U442 : BUF_X1 port map( A => n82_port, Z => n69_port);
   U443 : BUF_X1 port map( A => n48, Z => n35);
   U444 : BUF_X1 port map( A => n218, Z => n204);
   U445 : BUF_X1 port map( A => n184, Z => n170);
   U446 : BUF_X1 port map( A => n218, Z => n205);
   U447 : BUF_X1 port map( A => n184, Z => n171);
   U448 : BUF_X1 port map( A => n130_port, Z => n127_port);
   U449 : BUF_X1 port map( A => n130_port, Z => n128_port);
   U450 : BUF_X1 port map( A => n266, Z => n263);
   U451 : BUF_X1 port map( A => n266, Z => n264);
   U452 : BUF_X1 port map( A => n64_port, Z => n53);
   U453 : BUF_X1 port map( A => n30, Z => n19);
   U454 : BUF_X1 port map( A => n64_port, Z => n54);
   U455 : BUF_X1 port map( A => n30, Z => n20);
   U456 : BUF_X1 port map( A => n64_port, Z => n55);
   U457 : BUF_X1 port map( A => n30, Z => n21);
   U458 : BUF_X1 port map( A => n63_port, Z => n56);
   U459 : BUF_X1 port map( A => n29, Z => n22);
   U460 : BUF_X1 port map( A => n63_port, Z => n57);
   U461 : BUF_X1 port map( A => n29, Z => n23);
   U462 : BUF_X1 port map( A => n63_port, Z => n58);
   U463 : BUF_X1 port map( A => n29, Z => n24);
   U464 : BUF_X1 port map( A => n96, Z => n93);
   U465 : BUF_X1 port map( A => n96, Z => n94);
   U466 : BUF_X1 port map( A => n200, Z => n189);
   U467 : BUF_X1 port map( A => n166, Z => n155_port);
   U468 : BUF_X1 port map( A => n200, Z => n190);
   U469 : BUF_X1 port map( A => n166, Z => n156_port);
   U470 : BUF_X1 port map( A => n200, Z => n191);
   U471 : BUF_X1 port map( A => n166, Z => n157_port);
   U472 : BUF_X1 port map( A => n199, Z => n192);
   U473 : BUF_X1 port map( A => n165, Z => n158_port);
   U474 : BUF_X1 port map( A => n199, Z => n193);
   U475 : BUF_X1 port map( A => n165, Z => n159);
   U476 : BUF_X1 port map( A => n199, Z => n194);
   U477 : BUF_X1 port map( A => n165, Z => n160);
   U478 : BUF_X1 port map( A => n232, Z => n229);
   U479 : BUF_X1 port map( A => n232, Z => n230);
   U480 : BUF_X1 port map( A => n65_port, Z => n51);
   U481 : BUF_X1 port map( A => n31, Z => n17);
   U482 : BUF_X1 port map( A => n65_port, Z => n52);
   U483 : BUF_X1 port map( A => n31, Z => n18);
   U484 : BUF_X1 port map( A => n201, Z => n187);
   U485 : BUF_X1 port map( A => n167, Z => n153_port);
   U486 : BUF_X1 port map( A => n201, Z => n188);
   U487 : BUF_X1 port map( A => n167, Z => n154_port);
   U488 : BUF_X1 port map( A => n292, Z => n291);
   U489 : BUF_X1 port map( A => n147_port, Z => n146_port);
   U490 : BUF_X1 port map( A => n283, Z => n282);
   U491 : BUF_X1 port map( A => n113, Z => n112);
   U492 : BUF_X1 port map( A => n249, Z => n248);
   U493 : BUF_X1 port map( A => n130_port, Z => n129_port);
   U494 : BUF_X1 port map( A => n266, Z => n265);
   U495 : BUF_X1 port map( A => n96, Z => n95);
   U496 : BUF_X1 port map( A => n232, Z => n231);
   U497 : BUF_X1 port map( A => n10, Z => n152_port);
   U498 : BUF_X1 port map( A => n9, Z => n135_port);
   U499 : BUF_X1 port map( A => n16, Z => n288);
   U500 : BUF_X1 port map( A => n15, Z => n271);
   U501 : BUF_X1 port map( A => n8, Z => n118);
   U502 : BUF_X1 port map( A => n3, Z => n101);
   U503 : BUF_X1 port map( A => n14, Z => n254);
   U504 : BUF_X1 port map( A => n4, Z => n237);
   U505 : INV_X1 port map( A => RESET, ZN => n292);
   U506 : BUF_X1 port map( A => n83_port, Z => n82_port);
   U507 : BUF_X1 port map( A => n66_port, Z => n65_port);
   U508 : BUF_X1 port map( A => n49, Z => n48);
   U509 : BUF_X1 port map( A => n32, Z => n31);
   U510 : BUF_X1 port map( A => n219, Z => n218);
   U511 : BUF_X1 port map( A => n202, Z => n201);
   U512 : BUF_X1 port map( A => n185, Z => n184);
   U513 : BUF_X1 port map( A => n168, Z => n167);
   U514 : BUF_X1 port map( A => n79_port, Z => n76_port);
   U515 : BUF_X1 port map( A => n45, Z => n42);
   U516 : BUF_X1 port map( A => n79_port, Z => n77_port);
   U517 : BUF_X1 port map( A => n45, Z => n43);
   U518 : BUF_X1 port map( A => n215, Z => n212);
   U519 : BUF_X1 port map( A => n181, Z => n178);
   U520 : BUF_X1 port map( A => n215, Z => n213);
   U521 : BUF_X1 port map( A => n181, Z => n179);
   U522 : BUF_X1 port map( A => n62_port, Z => n59);
   U523 : BUF_X1 port map( A => n28, Z => n25);
   U524 : BUF_X1 port map( A => n62_port, Z => n60_port);
   U525 : BUF_X1 port map( A => n28, Z => n26);
   U526 : BUF_X1 port map( A => n198, Z => n195);
   U527 : BUF_X1 port map( A => n164, Z => n161);
   U528 : BUF_X1 port map( A => n198, Z => n196);
   U529 : BUF_X1 port map( A => n164, Z => n162);
   U530 : BUF_X1 port map( A => n79_port, Z => n78_port);
   U531 : BUF_X1 port map( A => n45, Z => n44);
   U532 : BUF_X1 port map( A => n215, Z => n214);
   U533 : BUF_X1 port map( A => n181, Z => n180);
   U534 : BUF_X1 port map( A => n62_port, Z => n61_port);
   U535 : BUF_X1 port map( A => n28, Z => n27);
   U536 : BUF_X1 port map( A => n198, Z => n197);
   U537 : BUF_X1 port map( A => n164, Z => n163);
   U538 : BUF_X1 port map( A => n7, Z => n84_port);
   U539 : BUF_X1 port map( A => n6, Z => n67_port);
   U540 : BUF_X1 port map( A => n5, Z => n50);
   U541 : BUF_X1 port map( A => n1, Z => n33);
   U542 : BUF_X1 port map( A => n13, Z => n220);
   U543 : BUF_X1 port map( A => n12, Z => n203);
   U544 : BUF_X1 port map( A => n11, Z => n186);
   U545 : BUF_X1 port map( A => n2, Z => n169);
   U546 : INV_X1 port map( A => ADD_RD1(0), ZN => n1119);
   U547 : INV_X1 port map( A => ADD_RD2(0), ZN => n2827);
   U548 : INV_X1 port map( A => ADD_RD1(2), ZN => n1117);
   U549 : INV_X1 port map( A => ADD_RD2(2), ZN => n2825);
   U550 : INV_X1 port map( A => ADD_RD1(3), ZN => n1116);
   U551 : INV_X1 port map( A => ADD_RD2(3), ZN => n2824);
   U552 : INV_X1 port map( A => ADD_RD1(1), ZN => n1118);
   U553 : INV_X1 port map( A => ADD_RD2(1), ZN => n2826);
   U554 : NOR2_X1 port map( A1 => n1117, A2 => ADD_RD1(1), ZN => n436);
   U555 : NOR2_X1 port map( A1 => n1117, A2 => n1118, ZN => n437);
   U556 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n34, B1 => 
                           REGISTERS_23_0_port, B2 => n17, ZN => n443);
   U557 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n438);
   U558 : NOR2_X1 port map( A1 => n1118, A2 => ADD_RD1(2), ZN => n439);
   U559 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n68_port, B1 => 
                           REGISTERS_19_0_port, B2 => n51, ZN => n442);
   U560 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n102, B1 => 
                           REGISTERS_22_0_port, B2 => n85_port, ZN => n441);
   U561 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n136_port, B1 => 
                           REGISTERS_18_0_port, B2 => n119, ZN => n440);
   U562 : AND4_X1 port map( A1 => n443, A2 => n442, A3 => n441, A4 => n440, ZN 
                           => n460);
   U563 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n34, B1 => 
                           REGISTERS_31_0_port, B2 => n17, ZN => n447);
   U564 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n68_port, B1 => 
                           REGISTERS_27_0_port, B2 => n51, ZN => n446);
   U565 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n102, B1 => 
                           REGISTERS_30_0_port, B2 => n85_port, ZN => n445);
   U566 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n136_port, B1 => 
                           REGISTERS_26_0_port, B2 => n119, ZN => n444);
   U567 : AND4_X1 port map( A1 => n447, A2 => n446, A3 => n445, A4 => n444, ZN 
                           => n459);
   U568 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n34, B1 => 
                           REGISTERS_7_0_port, B2 => n17, ZN => n451);
   U569 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n68_port, B1 => 
                           REGISTERS_3_0_port, B2 => n51, ZN => n450);
   U570 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n102, B1 => 
                           REGISTERS_6_0_port, B2 => n85_port, ZN => n449);
   U571 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n136_port, B1 => 
                           REGISTERS_2_0_port, B2 => n119, ZN => n448);
   U572 : NAND4_X1 port map( A1 => n451, A2 => n450, A3 => n449, A4 => n448, ZN
                           => n457);
   U573 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n34, B1 => 
                           REGISTERS_15_0_port, B2 => n17, ZN => n455);
   U574 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n68_port, B1 => 
                           REGISTERS_11_0_port, B2 => n51, ZN => n454);
   U575 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n102, B1 => 
                           REGISTERS_14_0_port, B2 => n85_port, ZN => n453);
   U576 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n136_port, B1 => 
                           REGISTERS_10_0_port, B2 => n119, ZN => n452);
   U577 : NAND4_X1 port map( A1 => n455, A2 => n454, A3 => n453, A4 => n452, ZN
                           => n456);
   U578 : AOI22_X1 port map( A1 => n457, A2 => n1110, B1 => n456, B2 => n1108, 
                           ZN => n458);
   U579 : OAI221_X1 port map( B1 => n1114, B2 => n460, C1 => n1112, C2 => n459,
                           A => n458, ZN => N91);
   U580 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n34, B1 => 
                           REGISTERS_23_1_port, B2 => n17, ZN => n464);
   U581 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n68_port, B1 => 
                           REGISTERS_19_1_port, B2 => n51, ZN => n463);
   U582 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n102, B1 => 
                           REGISTERS_22_1_port, B2 => n85_port, ZN => n462);
   U583 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n136_port, B1 => 
                           REGISTERS_18_1_port, B2 => n119, ZN => n461);
   U584 : AND4_X1 port map( A1 => n464, A2 => n463, A3 => n462, A4 => n461, ZN 
                           => n481);
   U585 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n34, B1 => 
                           REGISTERS_31_1_port, B2 => n17, ZN => n468);
   U586 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n68_port, B1 => 
                           REGISTERS_27_1_port, B2 => n51, ZN => n467);
   U587 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n102, B1 => 
                           REGISTERS_30_1_port, B2 => n85_port, ZN => n466);
   U588 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n136_port, B1 => 
                           REGISTERS_26_1_port, B2 => n119, ZN => n465);
   U589 : AND4_X1 port map( A1 => n468, A2 => n467, A3 => n466, A4 => n465, ZN 
                           => n480);
   U590 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n34, B1 => 
                           REGISTERS_7_1_port, B2 => n17, ZN => n472);
   U591 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n68_port, B1 => 
                           REGISTERS_3_1_port, B2 => n51, ZN => n471);
   U592 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n102, B1 => 
                           REGISTERS_6_1_port, B2 => n85_port, ZN => n470);
   U593 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n136_port, B1 => 
                           REGISTERS_2_1_port, B2 => n119, ZN => n469);
   U594 : NAND4_X1 port map( A1 => n472, A2 => n471, A3 => n470, A4 => n469, ZN
                           => n478);
   U595 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n34, B1 => 
                           REGISTERS_15_1_port, B2 => n17, ZN => n476);
   U596 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n68_port, B1 => 
                           REGISTERS_11_1_port, B2 => n51, ZN => n475);
   U597 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n102, B1 => 
                           REGISTERS_14_1_port, B2 => n85_port, ZN => n474);
   U598 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n136_port, B1 => 
                           REGISTERS_10_1_port, B2 => n119, ZN => n473);
   U599 : NAND4_X1 port map( A1 => n476, A2 => n475, A3 => n474, A4 => n473, ZN
                           => n477);
   U600 : AOI22_X1 port map( A1 => n478, A2 => n1110, B1 => n477, B2 => n1108, 
                           ZN => n479);
   U601 : OAI221_X1 port map( B1 => n1114, B2 => n481, C1 => n1112, C2 => n480,
                           A => n479, ZN => N90);
   U602 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n34, B1 => 
                           REGISTERS_23_2_port, B2 => n17, ZN => n485);
   U603 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n68_port, B1 => 
                           REGISTERS_19_2_port, B2 => n51, ZN => n484);
   U604 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n102, B1 => 
                           REGISTERS_22_2_port, B2 => n85_port, ZN => n483);
   U605 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n136_port, B1 => 
                           REGISTERS_18_2_port, B2 => n119, ZN => n482);
   U606 : AND4_X1 port map( A1 => n485, A2 => n484, A3 => n483, A4 => n482, ZN 
                           => n502);
   U607 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n34, B1 => 
                           REGISTERS_31_2_port, B2 => n17, ZN => n489);
   U608 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n68_port, B1 => 
                           REGISTERS_27_2_port, B2 => n51, ZN => n488);
   U609 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n102, B1 => 
                           REGISTERS_30_2_port, B2 => n85_port, ZN => n487);
   U610 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n136_port, B1 => 
                           REGISTERS_26_2_port, B2 => n119, ZN => n486);
   U611 : AND4_X1 port map( A1 => n489, A2 => n488, A3 => n487, A4 => n486, ZN 
                           => n501);
   U612 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n34, B1 => 
                           REGISTERS_7_2_port, B2 => n17, ZN => n493);
   U613 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n68_port, B1 => 
                           REGISTERS_3_2_port, B2 => n51, ZN => n492);
   U614 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n102, B1 => 
                           REGISTERS_6_2_port, B2 => n85_port, ZN => n491);
   U615 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n136_port, B1 => 
                           REGISTERS_2_2_port, B2 => n119, ZN => n490);
   U616 : NAND4_X1 port map( A1 => n493, A2 => n492, A3 => n491, A4 => n490, ZN
                           => n499);
   U617 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n34, B1 => 
                           REGISTERS_15_2_port, B2 => n17, ZN => n497);
   U618 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n68_port, B1 => 
                           REGISTERS_11_2_port, B2 => n51, ZN => n496);
   U619 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n102, B1 => 
                           REGISTERS_14_2_port, B2 => n85_port, ZN => n495);
   U620 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n136_port, B1 => 
                           REGISTERS_10_2_port, B2 => n119, ZN => n494);
   U621 : NAND4_X1 port map( A1 => n497, A2 => n496, A3 => n495, A4 => n494, ZN
                           => n498);
   U622 : AOI22_X1 port map( A1 => n499, A2 => n1110, B1 => n498, B2 => n1108, 
                           ZN => n500);
   U623 : OAI221_X1 port map( B1 => n1114, B2 => n502, C1 => n1112, C2 => n501,
                           A => n500, ZN => N89);
   U624 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n35, B1 => 
                           REGISTERS_23_3_port, B2 => n18, ZN => n506);
   U625 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n69_port, B1 => 
                           REGISTERS_19_3_port, B2 => n52, ZN => n505);
   U626 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n103, B1 => 
                           REGISTERS_22_3_port, B2 => n86_port, ZN => n504);
   U627 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n137_port, B1 => 
                           REGISTERS_18_3_port, B2 => n120, ZN => n503);
   U628 : AND4_X1 port map( A1 => n506, A2 => n505, A3 => n504, A4 => n503, ZN 
                           => n523);
   U629 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n35, B1 => 
                           REGISTERS_31_3_port, B2 => n18, ZN => n510);
   U630 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n69_port, B1 => 
                           REGISTERS_27_3_port, B2 => n52, ZN => n509);
   U631 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n103, B1 => 
                           REGISTERS_30_3_port, B2 => n86_port, ZN => n508);
   U632 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n137_port, B1 => 
                           REGISTERS_26_3_port, B2 => n120, ZN => n507);
   U633 : AND4_X1 port map( A1 => n510, A2 => n509, A3 => n508, A4 => n507, ZN 
                           => n522);
   U634 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n35, B1 => 
                           REGISTERS_7_3_port, B2 => n18, ZN => n514);
   U635 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n69_port, B1 => 
                           REGISTERS_3_3_port, B2 => n52, ZN => n513);
   U636 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n103, B1 => 
                           REGISTERS_6_3_port, B2 => n86_port, ZN => n512);
   U637 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n137_port, B1 => 
                           REGISTERS_2_3_port, B2 => n120, ZN => n511);
   U638 : NAND4_X1 port map( A1 => n514, A2 => n513, A3 => n512, A4 => n511, ZN
                           => n520);
   U639 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n35, B1 => 
                           REGISTERS_15_3_port, B2 => n18, ZN => n518);
   U640 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n69_port, B1 => 
                           REGISTERS_11_3_port, B2 => n52, ZN => n517);
   U641 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n103, B1 => 
                           REGISTERS_14_3_port, B2 => n86_port, ZN => n516);
   U642 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n137_port, B1 => 
                           REGISTERS_10_3_port, B2 => n120, ZN => n515);
   U643 : NAND4_X1 port map( A1 => n518, A2 => n517, A3 => n516, A4 => n515, ZN
                           => n519);
   U644 : AOI22_X1 port map( A1 => n520, A2 => n1110, B1 => n519, B2 => n1108, 
                           ZN => n521);
   U645 : OAI221_X1 port map( B1 => n1114, B2 => n523, C1 => n1112, C2 => n522,
                           A => n521, ZN => N88);
   U646 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n35, B1 => 
                           REGISTERS_23_4_port, B2 => n18, ZN => n527);
   U647 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n69_port, B1 => 
                           REGISTERS_19_4_port, B2 => n52, ZN => n526);
   U648 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n103, B1 => 
                           REGISTERS_22_4_port, B2 => n86_port, ZN => n525);
   U649 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n137_port, B1 => 
                           REGISTERS_18_4_port, B2 => n120, ZN => n524);
   U650 : AND4_X1 port map( A1 => n527, A2 => n526, A3 => n525, A4 => n524, ZN 
                           => n544);
   U651 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n35, B1 => 
                           REGISTERS_31_4_port, B2 => n18, ZN => n531);
   U652 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n69_port, B1 => 
                           REGISTERS_27_4_port, B2 => n52, ZN => n530);
   U653 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n103, B1 => 
                           REGISTERS_30_4_port, B2 => n86_port, ZN => n529);
   U654 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n137_port, B1 => 
                           REGISTERS_26_4_port, B2 => n120, ZN => n528);
   U655 : AND4_X1 port map( A1 => n531, A2 => n530, A3 => n529, A4 => n528, ZN 
                           => n543);
   U656 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n35, B1 => 
                           REGISTERS_7_4_port, B2 => n18, ZN => n535);
   U657 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n69_port, B1 => 
                           REGISTERS_3_4_port, B2 => n52, ZN => n534);
   U658 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n103, B1 => 
                           REGISTERS_6_4_port, B2 => n86_port, ZN => n533);
   U659 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n137_port, B1 => 
                           REGISTERS_2_4_port, B2 => n120, ZN => n532);
   U660 : NAND4_X1 port map( A1 => n535, A2 => n534, A3 => n533, A4 => n532, ZN
                           => n541);
   U661 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n35, B1 => 
                           REGISTERS_15_4_port, B2 => n18, ZN => n539);
   U662 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n69_port, B1 => 
                           REGISTERS_11_4_port, B2 => n52, ZN => n538);
   U663 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n103, B1 => 
                           REGISTERS_14_4_port, B2 => n86_port, ZN => n537);
   U664 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n137_port, B1 => 
                           REGISTERS_10_4_port, B2 => n120, ZN => n536);
   U665 : NAND4_X1 port map( A1 => n539, A2 => n538, A3 => n537, A4 => n536, ZN
                           => n540);
   U666 : AOI22_X1 port map( A1 => n541, A2 => n1110, B1 => n540, B2 => n1108, 
                           ZN => n542);
   U667 : OAI221_X1 port map( B1 => n1114, B2 => n544, C1 => n1112, C2 => n543,
                           A => n542, ZN => N87);
   U668 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n35, B1 => 
                           REGISTERS_23_5_port, B2 => n18, ZN => n548);
   U669 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n69_port, B1 => 
                           REGISTERS_19_5_port, B2 => n52, ZN => n547);
   U670 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n103, B1 => 
                           REGISTERS_22_5_port, B2 => n86_port, ZN => n546);
   U671 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n137_port, B1 => 
                           REGISTERS_18_5_port, B2 => n120, ZN => n545);
   U672 : AND4_X1 port map( A1 => n548, A2 => n547, A3 => n546, A4 => n545, ZN 
                           => n565);
   U673 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n35, B1 => 
                           REGISTERS_31_5_port, B2 => n18, ZN => n552);
   U674 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n69_port, B1 => 
                           REGISTERS_27_5_port, B2 => n52, ZN => n551);
   U675 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n103, B1 => 
                           REGISTERS_30_5_port, B2 => n86_port, ZN => n550);
   U676 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n137_port, B1 => 
                           REGISTERS_26_5_port, B2 => n120, ZN => n549);
   U677 : AND4_X1 port map( A1 => n552, A2 => n551, A3 => n550, A4 => n549, ZN 
                           => n564);
   U678 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n35, B1 => 
                           REGISTERS_7_5_port, B2 => n18, ZN => n556);
   U679 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n69_port, B1 => 
                           REGISTERS_3_5_port, B2 => n52, ZN => n555);
   U680 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n103, B1 => 
                           REGISTERS_6_5_port, B2 => n86_port, ZN => n554);
   U681 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n137_port, B1 => 
                           REGISTERS_2_5_port, B2 => n120, ZN => n553);
   U682 : NAND4_X1 port map( A1 => n556, A2 => n555, A3 => n554, A4 => n553, ZN
                           => n562);
   U683 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n35, B1 => 
                           REGISTERS_15_5_port, B2 => n18, ZN => n560);
   U684 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n69_port, B1 => 
                           REGISTERS_11_5_port, B2 => n52, ZN => n559);
   U685 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n103, B1 => 
                           REGISTERS_14_5_port, B2 => n86_port, ZN => n558);
   U686 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n137_port, B1 => 
                           REGISTERS_10_5_port, B2 => n120, ZN => n557);
   U687 : NAND4_X1 port map( A1 => n560, A2 => n559, A3 => n558, A4 => n557, ZN
                           => n561);
   U688 : AOI22_X1 port map( A1 => n562, A2 => n1110, B1 => n561, B2 => n1108, 
                           ZN => n563);
   U689 : OAI221_X1 port map( B1 => n1114, B2 => n565, C1 => n1112, C2 => n564,
                           A => n563, ZN => N86);
   U690 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n36, B1 => 
                           REGISTERS_23_6_port, B2 => n19, ZN => n569);
   U691 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n70_port, B1 => 
                           REGISTERS_19_6_port, B2 => n53, ZN => n568);
   U692 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n104, B1 => 
                           REGISTERS_22_6_port, B2 => n87_port, ZN => n567);
   U693 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n138_port, B1 => 
                           REGISTERS_18_6_port, B2 => n121, ZN => n566);
   U694 : AND4_X1 port map( A1 => n569, A2 => n568, A3 => n567, A4 => n566, ZN 
                           => n586);
   U695 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n36, B1 => 
                           REGISTERS_31_6_port, B2 => n19, ZN => n573);
   U696 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n70_port, B1 => 
                           REGISTERS_27_6_port, B2 => n53, ZN => n572);
   U697 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n104, B1 => 
                           REGISTERS_30_6_port, B2 => n87_port, ZN => n571);
   U698 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n138_port, B1 => 
                           REGISTERS_26_6_port, B2 => n121, ZN => n570);
   U699 : AND4_X1 port map( A1 => n573, A2 => n572, A3 => n571, A4 => n570, ZN 
                           => n585);
   U700 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n36, B1 => 
                           REGISTERS_7_6_port, B2 => n19, ZN => n577);
   U701 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n70_port, B1 => 
                           REGISTERS_3_6_port, B2 => n53, ZN => n576);
   U702 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n104, B1 => 
                           REGISTERS_6_6_port, B2 => n87_port, ZN => n575);
   U703 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n138_port, B1 => 
                           REGISTERS_2_6_port, B2 => n121, ZN => n574);
   U704 : NAND4_X1 port map( A1 => n577, A2 => n576, A3 => n575, A4 => n574, ZN
                           => n583);
   U705 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n36, B1 => 
                           REGISTERS_15_6_port, B2 => n19, ZN => n581);
   U706 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n70_port, B1 => 
                           REGISTERS_11_6_port, B2 => n53, ZN => n580);
   U707 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n104, B1 => 
                           REGISTERS_14_6_port, B2 => n87_port, ZN => n579);
   U708 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n138_port, B1 => 
                           REGISTERS_10_6_port, B2 => n121, ZN => n578);
   U709 : NAND4_X1 port map( A1 => n581, A2 => n580, A3 => n579, A4 => n578, ZN
                           => n582);
   U710 : AOI22_X1 port map( A1 => n583, A2 => n1110, B1 => n582, B2 => n1108, 
                           ZN => n584);
   U711 : OAI221_X1 port map( B1 => n1114, B2 => n586, C1 => n1112, C2 => n585,
                           A => n584, ZN => N85);
   U712 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n36, B1 => 
                           REGISTERS_23_7_port, B2 => n19, ZN => n590);
   U713 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n70_port, B1 => 
                           REGISTERS_19_7_port, B2 => n53, ZN => n589);
   U714 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n104, B1 => 
                           REGISTERS_22_7_port, B2 => n87_port, ZN => n588);
   U715 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n138_port, B1 => 
                           REGISTERS_18_7_port, B2 => n121, ZN => n587);
   U716 : AND4_X1 port map( A1 => n590, A2 => n589, A3 => n588, A4 => n587, ZN 
                           => n607);
   U717 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n36, B1 => 
                           REGISTERS_31_7_port, B2 => n19, ZN => n594);
   U718 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n70_port, B1 => 
                           REGISTERS_27_7_port, B2 => n53, ZN => n593);
   U719 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n104, B1 => 
                           REGISTERS_30_7_port, B2 => n87_port, ZN => n592);
   U720 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n138_port, B1 => 
                           REGISTERS_26_7_port, B2 => n121, ZN => n591);
   U721 : AND4_X1 port map( A1 => n594, A2 => n593, A3 => n592, A4 => n591, ZN 
                           => n606);
   U722 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n36, B1 => 
                           REGISTERS_7_7_port, B2 => n19, ZN => n598);
   U723 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n70_port, B1 => 
                           REGISTERS_3_7_port, B2 => n53, ZN => n597);
   U724 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n104, B1 => 
                           REGISTERS_6_7_port, B2 => n87_port, ZN => n596);
   U725 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n138_port, B1 => 
                           REGISTERS_2_7_port, B2 => n121, ZN => n595);
   U726 : NAND4_X1 port map( A1 => n598, A2 => n597, A3 => n596, A4 => n595, ZN
                           => n604);
   U727 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n36, B1 => 
                           REGISTERS_15_7_port, B2 => n19, ZN => n602);
   U728 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n70_port, B1 => 
                           REGISTERS_11_7_port, B2 => n53, ZN => n601);
   U729 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n104, B1 => 
                           REGISTERS_14_7_port, B2 => n87_port, ZN => n600);
   U730 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n138_port, B1 => 
                           REGISTERS_10_7_port, B2 => n121, ZN => n599);
   U731 : NAND4_X1 port map( A1 => n602, A2 => n601, A3 => n600, A4 => n599, ZN
                           => n603);
   U732 : AOI22_X1 port map( A1 => n604, A2 => n1110, B1 => n603, B2 => n1108, 
                           ZN => n605);
   U733 : OAI221_X1 port map( B1 => n1114, B2 => n607, C1 => n1112, C2 => n606,
                           A => n605, ZN => N84);
   U734 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n36, B1 => 
                           REGISTERS_23_8_port, B2 => n19, ZN => n611);
   U735 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n70_port, B1 => 
                           REGISTERS_19_8_port, B2 => n53, ZN => n610);
   U736 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n104, B1 => 
                           REGISTERS_22_8_port, B2 => n87_port, ZN => n609);
   U737 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n138_port, B1 => 
                           REGISTERS_18_8_port, B2 => n121, ZN => n608);
   U738 : AND4_X1 port map( A1 => n611, A2 => n610, A3 => n609, A4 => n608, ZN 
                           => n628);
   U739 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n36, B1 => 
                           REGISTERS_31_8_port, B2 => n19, ZN => n615);
   U740 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n70_port, B1 => 
                           REGISTERS_27_8_port, B2 => n53, ZN => n614);
   U741 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n104, B1 => 
                           REGISTERS_30_8_port, B2 => n87_port, ZN => n613);
   U742 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n138_port, B1 => 
                           REGISTERS_26_8_port, B2 => n121, ZN => n612);
   U743 : AND4_X1 port map( A1 => n615, A2 => n614, A3 => n613, A4 => n612, ZN 
                           => n627);
   U744 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n36, B1 => 
                           REGISTERS_7_8_port, B2 => n19, ZN => n619);
   U745 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n70_port, B1 => 
                           REGISTERS_3_8_port, B2 => n53, ZN => n618);
   U746 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n104, B1 => 
                           REGISTERS_6_8_port, B2 => n87_port, ZN => n617);
   U747 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n138_port, B1 => 
                           REGISTERS_2_8_port, B2 => n121, ZN => n616);
   U748 : NAND4_X1 port map( A1 => n619, A2 => n618, A3 => n617, A4 => n616, ZN
                           => n625);
   U749 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n36, B1 => 
                           REGISTERS_15_8_port, B2 => n19, ZN => n623);
   U750 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n70_port, B1 => 
                           REGISTERS_11_8_port, B2 => n53, ZN => n622);
   U751 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n104, B1 => 
                           REGISTERS_14_8_port, B2 => n87_port, ZN => n621);
   U752 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n138_port, B1 => 
                           REGISTERS_10_8_port, B2 => n121, ZN => n620);
   U753 : NAND4_X1 port map( A1 => n623, A2 => n622, A3 => n621, A4 => n620, ZN
                           => n624);
   U754 : AOI22_X1 port map( A1 => n625, A2 => n1110, B1 => n624, B2 => n1108, 
                           ZN => n626);
   U755 : OAI221_X1 port map( B1 => n1114, B2 => n628, C1 => n1112, C2 => n627,
                           A => n626, ZN => N83);
   U756 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n37, B1 => 
                           REGISTERS_23_9_port, B2 => n20, ZN => n632);
   U757 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n71_port, B1 => 
                           REGISTERS_19_9_port, B2 => n54, ZN => n631);
   U758 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n105, B1 => 
                           REGISTERS_22_9_port, B2 => n88_port, ZN => n630);
   U759 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n139_port, B1 => 
                           REGISTERS_18_9_port, B2 => n122, ZN => n629);
   U760 : AND4_X1 port map( A1 => n632, A2 => n631, A3 => n630, A4 => n629, ZN 
                           => n649);
   U761 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n37, B1 => 
                           REGISTERS_31_9_port, B2 => n20, ZN => n636);
   U762 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n71_port, B1 => 
                           REGISTERS_27_9_port, B2 => n54, ZN => n635);
   U763 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n105, B1 => 
                           REGISTERS_30_9_port, B2 => n88_port, ZN => n634);
   U764 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n139_port, B1 => 
                           REGISTERS_26_9_port, B2 => n122, ZN => n633);
   U765 : AND4_X1 port map( A1 => n636, A2 => n635, A3 => n634, A4 => n633, ZN 
                           => n648);
   U766 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n37, B1 => 
                           REGISTERS_7_9_port, B2 => n20, ZN => n640);
   U767 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n71_port, B1 => 
                           REGISTERS_3_9_port, B2 => n54, ZN => n639);
   U768 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n105, B1 => 
                           REGISTERS_6_9_port, B2 => n88_port, ZN => n638);
   U769 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n139_port, B1 => 
                           REGISTERS_2_9_port, B2 => n122, ZN => n637);
   U770 : NAND4_X1 port map( A1 => n640, A2 => n639, A3 => n638, A4 => n637, ZN
                           => n646);
   U771 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n37, B1 => 
                           REGISTERS_15_9_port, B2 => n20, ZN => n644);
   U772 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n71_port, B1 => 
                           REGISTERS_11_9_port, B2 => n54, ZN => n643);
   U773 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n105, B1 => 
                           REGISTERS_14_9_port, B2 => n88_port, ZN => n642);
   U774 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n139_port, B1 => 
                           REGISTERS_10_9_port, B2 => n122, ZN => n641);
   U775 : NAND4_X1 port map( A1 => n644, A2 => n643, A3 => n642, A4 => n641, ZN
                           => n645);
   U776 : AOI22_X1 port map( A1 => n646, A2 => n1110, B1 => n645, B2 => n1108, 
                           ZN => n647);
   U777 : OAI221_X1 port map( B1 => n1114, B2 => n649, C1 => n1112, C2 => n648,
                           A => n647, ZN => N82);
   U778 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n37, B1 => 
                           REGISTERS_23_10_port, B2 => n20, ZN => n653);
   U779 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n71_port, B1 => 
                           REGISTERS_19_10_port, B2 => n54, ZN => n652);
   U780 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n105, B1 => 
                           REGISTERS_22_10_port, B2 => n88_port, ZN => n651);
   U781 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n139_port, B1 =>
                           REGISTERS_18_10_port, B2 => n122, ZN => n650);
   U782 : AND4_X1 port map( A1 => n653, A2 => n652, A3 => n651, A4 => n650, ZN 
                           => n670);
   U783 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n37, B1 => 
                           REGISTERS_31_10_port, B2 => n20, ZN => n657);
   U784 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n71_port, B1 => 
                           REGISTERS_27_10_port, B2 => n54, ZN => n656);
   U785 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n105, B1 => 
                           REGISTERS_30_10_port, B2 => n88_port, ZN => n655);
   U786 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n139_port, B1 =>
                           REGISTERS_26_10_port, B2 => n122, ZN => n654);
   U787 : AND4_X1 port map( A1 => n657, A2 => n656, A3 => n655, A4 => n654, ZN 
                           => n669);
   U788 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n37, B1 => 
                           REGISTERS_7_10_port, B2 => n20, ZN => n661);
   U789 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n71_port, B1 => 
                           REGISTERS_3_10_port, B2 => n54, ZN => n660);
   U790 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n105, B1 => 
                           REGISTERS_6_10_port, B2 => n88_port, ZN => n659);
   U791 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n139_port, B1 => 
                           REGISTERS_2_10_port, B2 => n122, ZN => n658);
   U792 : NAND4_X1 port map( A1 => n661, A2 => n660, A3 => n659, A4 => n658, ZN
                           => n667);
   U793 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n37, B1 => 
                           REGISTERS_15_10_port, B2 => n20, ZN => n665);
   U794 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n71_port, B1 => 
                           REGISTERS_11_10_port, B2 => n54, ZN => n664);
   U795 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n105, B1 => 
                           REGISTERS_14_10_port, B2 => n88_port, ZN => n663);
   U796 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n139_port, B1 => 
                           REGISTERS_10_10_port, B2 => n122, ZN => n662);
   U797 : NAND4_X1 port map( A1 => n665, A2 => n664, A3 => n663, A4 => n662, ZN
                           => n666);
   U798 : AOI22_X1 port map( A1 => n667, A2 => n1110, B1 => n666, B2 => n1108, 
                           ZN => n668);
   U799 : OAI221_X1 port map( B1 => n1114, B2 => n670, C1 => n1112, C2 => n669,
                           A => n668, ZN => N81);
   U800 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n37, B1 => 
                           REGISTERS_23_11_port, B2 => n20, ZN => n674);
   U801 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n71_port, B1 => 
                           REGISTERS_19_11_port, B2 => n54, ZN => n673);
   U802 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n105, B1 => 
                           REGISTERS_22_11_port, B2 => n88_port, ZN => n672);
   U803 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n139_port, B1 =>
                           REGISTERS_18_11_port, B2 => n122, ZN => n671);
   U804 : AND4_X1 port map( A1 => n674, A2 => n673, A3 => n672, A4 => n671, ZN 
                           => n691);
   U805 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n37, B1 => 
                           REGISTERS_31_11_port, B2 => n20, ZN => n678);
   U806 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n71_port, B1 => 
                           REGISTERS_27_11_port, B2 => n54, ZN => n677);
   U807 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n105, B1 => 
                           REGISTERS_30_11_port, B2 => n88_port, ZN => n676);
   U808 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n139_port, B1 =>
                           REGISTERS_26_11_port, B2 => n122, ZN => n675);
   U809 : AND4_X1 port map( A1 => n678, A2 => n677, A3 => n676, A4 => n675, ZN 
                           => n690);
   U810 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n37, B1 => 
                           REGISTERS_7_11_port, B2 => n20, ZN => n682);
   U811 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n71_port, B1 => 
                           REGISTERS_3_11_port, B2 => n54, ZN => n681);
   U812 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n105, B1 => 
                           REGISTERS_6_11_port, B2 => n88_port, ZN => n680);
   U813 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n139_port, B1 => 
                           REGISTERS_2_11_port, B2 => n122, ZN => n679);
   U814 : NAND4_X1 port map( A1 => n682, A2 => n681, A3 => n680, A4 => n679, ZN
                           => n688);
   U815 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n37, B1 => 
                           REGISTERS_15_11_port, B2 => n20, ZN => n686);
   U816 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n71_port, B1 => 
                           REGISTERS_11_11_port, B2 => n54, ZN => n685);
   U817 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n105, B1 => 
                           REGISTERS_14_11_port, B2 => n88_port, ZN => n684);
   U818 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n139_port, B1 => 
                           REGISTERS_10_11_port, B2 => n122, ZN => n683);
   U819 : NAND4_X1 port map( A1 => n686, A2 => n685, A3 => n684, A4 => n683, ZN
                           => n687);
   U820 : AOI22_X1 port map( A1 => n688, A2 => n1110, B1 => n687, B2 => n1108, 
                           ZN => n689);
   U821 : OAI221_X1 port map( B1 => n1114, B2 => n691, C1 => n1112, C2 => n690,
                           A => n689, ZN => N80);
   U822 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n38, B1 => 
                           REGISTERS_23_12_port, B2 => n21, ZN => n695);
   U823 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n72_port, B1 => 
                           REGISTERS_19_12_port, B2 => n55, ZN => n694);
   U824 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n106, B1 => 
                           REGISTERS_22_12_port, B2 => n89_port, ZN => n693);
   U825 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n140_port, B1 =>
                           REGISTERS_18_12_port, B2 => n123, ZN => n692);
   U826 : AND4_X1 port map( A1 => n695, A2 => n694, A3 => n693, A4 => n692, ZN 
                           => n712);
   U827 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n38, B1 => 
                           REGISTERS_31_12_port, B2 => n21, ZN => n699);
   U828 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n72_port, B1 => 
                           REGISTERS_27_12_port, B2 => n55, ZN => n698);
   U829 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n106, B1 => 
                           REGISTERS_30_12_port, B2 => n89_port, ZN => n697);
   U830 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n140_port, B1 =>
                           REGISTERS_26_12_port, B2 => n123, ZN => n696);
   U831 : AND4_X1 port map( A1 => n699, A2 => n698, A3 => n697, A4 => n696, ZN 
                           => n711);
   U832 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n38, B1 => 
                           REGISTERS_7_12_port, B2 => n21, ZN => n703);
   U833 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n72_port, B1 => 
                           REGISTERS_3_12_port, B2 => n55, ZN => n702);
   U834 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n106, B1 => 
                           REGISTERS_6_12_port, B2 => n89_port, ZN => n701);
   U835 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n140_port, B1 => 
                           REGISTERS_2_12_port, B2 => n123, ZN => n700);
   U836 : NAND4_X1 port map( A1 => n703, A2 => n702, A3 => n701, A4 => n700, ZN
                           => n709);
   U837 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n38, B1 => 
                           REGISTERS_15_12_port, B2 => n21, ZN => n707);
   U838 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n72_port, B1 => 
                           REGISTERS_11_12_port, B2 => n55, ZN => n706);
   U839 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n106, B1 => 
                           REGISTERS_14_12_port, B2 => n89_port, ZN => n705);
   U840 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n140_port, B1 => 
                           REGISTERS_10_12_port, B2 => n123, ZN => n704);
   U841 : NAND4_X1 port map( A1 => n707, A2 => n706, A3 => n705, A4 => n704, ZN
                           => n708);
   U842 : AOI22_X1 port map( A1 => n709, A2 => n1110, B1 => n708, B2 => n1108, 
                           ZN => n710);
   U843 : OAI221_X1 port map( B1 => n1114, B2 => n712, C1 => n1112, C2 => n711,
                           A => n710, ZN => N79);
   U844 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n38, B1 => 
                           REGISTERS_23_13_port, B2 => n21, ZN => n716);
   U845 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n72_port, B1 => 
                           REGISTERS_19_13_port, B2 => n55, ZN => n715);
   U846 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n106, B1 => 
                           REGISTERS_22_13_port, B2 => n89_port, ZN => n714);
   U847 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n140_port, B1 =>
                           REGISTERS_18_13_port, B2 => n123, ZN => n713);
   U848 : AND4_X1 port map( A1 => n716, A2 => n715, A3 => n714, A4 => n713, ZN 
                           => n733);
   U849 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n38, B1 => 
                           REGISTERS_31_13_port, B2 => n21, ZN => n720);
   U850 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n72_port, B1 => 
                           REGISTERS_27_13_port, B2 => n55, ZN => n719);
   U851 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n106, B1 => 
                           REGISTERS_30_13_port, B2 => n89_port, ZN => n718);
   U852 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n140_port, B1 =>
                           REGISTERS_26_13_port, B2 => n123, ZN => n717);
   U853 : AND4_X1 port map( A1 => n720, A2 => n719, A3 => n718, A4 => n717, ZN 
                           => n732);
   U854 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n38, B1 => 
                           REGISTERS_7_13_port, B2 => n21, ZN => n724);
   U855 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n72_port, B1 => 
                           REGISTERS_3_13_port, B2 => n55, ZN => n723);
   U856 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n106, B1 => 
                           REGISTERS_6_13_port, B2 => n89_port, ZN => n722);
   U857 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n140_port, B1 => 
                           REGISTERS_2_13_port, B2 => n123, ZN => n721);
   U858 : NAND4_X1 port map( A1 => n724, A2 => n723, A3 => n722, A4 => n721, ZN
                           => n730);
   U859 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n38, B1 => 
                           REGISTERS_15_13_port, B2 => n21, ZN => n728);
   U860 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n72_port, B1 => 
                           REGISTERS_11_13_port, B2 => n55, ZN => n727);
   U861 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n106, B1 => 
                           REGISTERS_14_13_port, B2 => n89_port, ZN => n726);
   U862 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n140_port, B1 => 
                           REGISTERS_10_13_port, B2 => n123, ZN => n725);
   U863 : NAND4_X1 port map( A1 => n728, A2 => n727, A3 => n726, A4 => n725, ZN
                           => n729);
   U864 : AOI22_X1 port map( A1 => n730, A2 => n1110, B1 => n729, B2 => n1108, 
                           ZN => n731);
   U865 : OAI221_X1 port map( B1 => n1114, B2 => n733, C1 => n1112, C2 => n732,
                           A => n731, ZN => N78);
   U866 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n38, B1 => 
                           REGISTERS_23_14_port, B2 => n21, ZN => n737);
   U867 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n72_port, B1 => 
                           REGISTERS_19_14_port, B2 => n55, ZN => n736);
   U868 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n106, B1 => 
                           REGISTERS_22_14_port, B2 => n89_port, ZN => n735);
   U869 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n140_port, B1 =>
                           REGISTERS_18_14_port, B2 => n123, ZN => n734);
   U870 : AND4_X1 port map( A1 => n737, A2 => n736, A3 => n735, A4 => n734, ZN 
                           => n754);
   U871 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n38, B1 => 
                           REGISTERS_31_14_port, B2 => n21, ZN => n741);
   U872 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n72_port, B1 => 
                           REGISTERS_27_14_port, B2 => n55, ZN => n740);
   U873 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n106, B1 => 
                           REGISTERS_30_14_port, B2 => n89_port, ZN => n739);
   U874 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n140_port, B1 =>
                           REGISTERS_26_14_port, B2 => n123, ZN => n738);
   U875 : AND4_X1 port map( A1 => n741, A2 => n740, A3 => n739, A4 => n738, ZN 
                           => n753);
   U876 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n38, B1 => 
                           REGISTERS_7_14_port, B2 => n21, ZN => n745);
   U877 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n72_port, B1 => 
                           REGISTERS_3_14_port, B2 => n55, ZN => n744);
   U878 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n106, B1 => 
                           REGISTERS_6_14_port, B2 => n89_port, ZN => n743);
   U879 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n140_port, B1 => 
                           REGISTERS_2_14_port, B2 => n123, ZN => n742);
   U880 : NAND4_X1 port map( A1 => n745, A2 => n744, A3 => n743, A4 => n742, ZN
                           => n751);
   U881 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n38, B1 => 
                           REGISTERS_15_14_port, B2 => n21, ZN => n749);
   U882 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n72_port, B1 => 
                           REGISTERS_11_14_port, B2 => n55, ZN => n748);
   U883 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n106, B1 => 
                           REGISTERS_14_14_port, B2 => n89_port, ZN => n747);
   U884 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n140_port, B1 => 
                           REGISTERS_10_14_port, B2 => n123, ZN => n746);
   U885 : NAND4_X1 port map( A1 => n749, A2 => n748, A3 => n747, A4 => n746, ZN
                           => n750);
   U886 : AOI22_X1 port map( A1 => n751, A2 => n1110, B1 => n750, B2 => n1108, 
                           ZN => n752);
   U887 : OAI221_X1 port map( B1 => n1114, B2 => n754, C1 => n1112, C2 => n753,
                           A => n752, ZN => N77);
   U888 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n39, B1 => 
                           REGISTERS_23_15_port, B2 => n22, ZN => n758);
   U889 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n73_port, B1 => 
                           REGISTERS_19_15_port, B2 => n56, ZN => n757);
   U890 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n107, B1 => 
                           REGISTERS_22_15_port, B2 => n90_port, ZN => n756);
   U891 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n141_port, B1 =>
                           REGISTERS_18_15_port, B2 => n124, ZN => n755);
   U892 : AND4_X1 port map( A1 => n758, A2 => n757, A3 => n756, A4 => n755, ZN 
                           => n775);
   U893 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n39, B1 => 
                           REGISTERS_31_15_port, B2 => n22, ZN => n762);
   U894 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n73_port, B1 => 
                           REGISTERS_27_15_port, B2 => n56, ZN => n761);
   U895 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n107, B1 => 
                           REGISTERS_30_15_port, B2 => n90_port, ZN => n760);
   U896 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n141_port, B1 =>
                           REGISTERS_26_15_port, B2 => n124, ZN => n759);
   U897 : AND4_X1 port map( A1 => n762, A2 => n761, A3 => n760, A4 => n759, ZN 
                           => n774);
   U898 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n39, B1 => 
                           REGISTERS_7_15_port, B2 => n22, ZN => n766);
   U899 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n73_port, B1 => 
                           REGISTERS_3_15_port, B2 => n56, ZN => n765);
   U900 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n107, B1 => 
                           REGISTERS_6_15_port, B2 => n90_port, ZN => n764);
   U901 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n141_port, B1 => 
                           REGISTERS_2_15_port, B2 => n124, ZN => n763);
   U902 : NAND4_X1 port map( A1 => n766, A2 => n765, A3 => n764, A4 => n763, ZN
                           => n772);
   U903 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n39, B1 => 
                           REGISTERS_15_15_port, B2 => n22, ZN => n770);
   U904 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n73_port, B1 => 
                           REGISTERS_11_15_port, B2 => n56, ZN => n769);
   U905 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n107, B1 => 
                           REGISTERS_14_15_port, B2 => n90_port, ZN => n768);
   U906 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n141_port, B1 => 
                           REGISTERS_10_15_port, B2 => n124, ZN => n767);
   U907 : NAND4_X1 port map( A1 => n770, A2 => n769, A3 => n768, A4 => n767, ZN
                           => n771);
   U908 : AOI22_X1 port map( A1 => n772, A2 => n1110, B1 => n771, B2 => n1108, 
                           ZN => n773);
   U909 : OAI221_X1 port map( B1 => n1114, B2 => n775, C1 => n1112, C2 => n774,
                           A => n773, ZN => N76);
   U910 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n39, B1 => 
                           REGISTERS_23_16_port, B2 => n22, ZN => n779);
   U911 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n73_port, B1 => 
                           REGISTERS_19_16_port, B2 => n56, ZN => n778);
   U912 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n107, B1 => 
                           REGISTERS_22_16_port, B2 => n90_port, ZN => n777);
   U913 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n141_port, B1 =>
                           REGISTERS_18_16_port, B2 => n124, ZN => n776);
   U914 : AND4_X1 port map( A1 => n779, A2 => n778, A3 => n777, A4 => n776, ZN 
                           => n796);
   U915 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n39, B1 => 
                           REGISTERS_31_16_port, B2 => n22, ZN => n783);
   U916 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n73_port, B1 => 
                           REGISTERS_27_16_port, B2 => n56, ZN => n782);
   U917 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n107, B1 => 
                           REGISTERS_30_16_port, B2 => n90_port, ZN => n781);
   U918 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n141_port, B1 =>
                           REGISTERS_26_16_port, B2 => n124, ZN => n780);
   U919 : AND4_X1 port map( A1 => n783, A2 => n782, A3 => n781, A4 => n780, ZN 
                           => n795);
   U920 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n39, B1 => 
                           REGISTERS_7_16_port, B2 => n22, ZN => n787);
   U921 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n73_port, B1 => 
                           REGISTERS_3_16_port, B2 => n56, ZN => n786);
   U922 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n107, B1 => 
                           REGISTERS_6_16_port, B2 => n90_port, ZN => n785);
   U923 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n141_port, B1 => 
                           REGISTERS_2_16_port, B2 => n124, ZN => n784);
   U924 : NAND4_X1 port map( A1 => n787, A2 => n786, A3 => n785, A4 => n784, ZN
                           => n793);
   U925 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n39, B1 => 
                           REGISTERS_15_16_port, B2 => n22, ZN => n791);
   U926 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n73_port, B1 => 
                           REGISTERS_11_16_port, B2 => n56, ZN => n790);
   U927 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n107, B1 => 
                           REGISTERS_14_16_port, B2 => n90_port, ZN => n789);
   U928 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n141_port, B1 => 
                           REGISTERS_10_16_port, B2 => n124, ZN => n788);
   U929 : NAND4_X1 port map( A1 => n791, A2 => n790, A3 => n789, A4 => n788, ZN
                           => n792);
   U930 : AOI22_X1 port map( A1 => n793, A2 => n1110, B1 => n792, B2 => n1108, 
                           ZN => n794);
   U931 : OAI221_X1 port map( B1 => n1114, B2 => n796, C1 => n1112, C2 => n795,
                           A => n794, ZN => N75);
   U932 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n39, B1 => 
                           REGISTERS_23_17_port, B2 => n22, ZN => n800);
   U933 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n73_port, B1 => 
                           REGISTERS_19_17_port, B2 => n56, ZN => n799);
   U934 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n107, B1 => 
                           REGISTERS_22_17_port, B2 => n90_port, ZN => n798);
   U935 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n141_port, B1 =>
                           REGISTERS_18_17_port, B2 => n124, ZN => n797);
   U936 : AND4_X1 port map( A1 => n800, A2 => n799, A3 => n798, A4 => n797, ZN 
                           => n817);
   U937 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n39, B1 => 
                           REGISTERS_31_17_port, B2 => n22, ZN => n804);
   U938 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n73_port, B1 => 
                           REGISTERS_27_17_port, B2 => n56, ZN => n803);
   U939 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n107, B1 => 
                           REGISTERS_30_17_port, B2 => n90_port, ZN => n802);
   U940 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n141_port, B1 =>
                           REGISTERS_26_17_port, B2 => n124, ZN => n801);
   U941 : AND4_X1 port map( A1 => n804, A2 => n803, A3 => n802, A4 => n801, ZN 
                           => n816);
   U942 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n39, B1 => 
                           REGISTERS_7_17_port, B2 => n22, ZN => n808);
   U943 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n73_port, B1 => 
                           REGISTERS_3_17_port, B2 => n56, ZN => n807);
   U944 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n107, B1 => 
                           REGISTERS_6_17_port, B2 => n90_port, ZN => n806);
   U945 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n141_port, B1 => 
                           REGISTERS_2_17_port, B2 => n124, ZN => n805);
   U946 : NAND4_X1 port map( A1 => n808, A2 => n807, A3 => n806, A4 => n805, ZN
                           => n814);
   U947 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n39, B1 => 
                           REGISTERS_15_17_port, B2 => n22, ZN => n812);
   U948 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n73_port, B1 => 
                           REGISTERS_11_17_port, B2 => n56, ZN => n811);
   U949 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n107, B1 => 
                           REGISTERS_14_17_port, B2 => n90_port, ZN => n810);
   U950 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n141_port, B1 => 
                           REGISTERS_10_17_port, B2 => n124, ZN => n809);
   U951 : NAND4_X1 port map( A1 => n812, A2 => n811, A3 => n810, A4 => n809, ZN
                           => n813);
   U952 : AOI22_X1 port map( A1 => n814, A2 => n1110, B1 => n813, B2 => n1108, 
                           ZN => n815);
   U953 : OAI221_X1 port map( B1 => n1114, B2 => n817, C1 => n1112, C2 => n816,
                           A => n815, ZN => N74);
   U954 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n40, B1 => 
                           REGISTERS_23_18_port, B2 => n23, ZN => n821);
   U955 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n74_port, B1 => 
                           REGISTERS_19_18_port, B2 => n57, ZN => n820);
   U956 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n108, B1 => 
                           REGISTERS_22_18_port, B2 => n91_port, ZN => n819);
   U957 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n142_port, B1 =>
                           REGISTERS_18_18_port, B2 => n125, ZN => n818);
   U958 : AND4_X1 port map( A1 => n821, A2 => n820, A3 => n819, A4 => n818, ZN 
                           => n838);
   U959 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n40, B1 => 
                           REGISTERS_31_18_port, B2 => n23, ZN => n825);
   U960 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n74_port, B1 => 
                           REGISTERS_27_18_port, B2 => n57, ZN => n824);
   U961 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n108, B1 => 
                           REGISTERS_30_18_port, B2 => n91_port, ZN => n823);
   U962 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n142_port, B1 =>
                           REGISTERS_26_18_port, B2 => n125, ZN => n822);
   U963 : AND4_X1 port map( A1 => n825, A2 => n824, A3 => n823, A4 => n822, ZN 
                           => n837);
   U964 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n40, B1 => 
                           REGISTERS_7_18_port, B2 => n23, ZN => n829);
   U965 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n74_port, B1 => 
                           REGISTERS_3_18_port, B2 => n57, ZN => n828);
   U966 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n108, B1 => 
                           REGISTERS_6_18_port, B2 => n91_port, ZN => n827);
   U967 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n142_port, B1 => 
                           REGISTERS_2_18_port, B2 => n125, ZN => n826);
   U968 : NAND4_X1 port map( A1 => n829, A2 => n828, A3 => n827, A4 => n826, ZN
                           => n835);
   U969 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n40, B1 => 
                           REGISTERS_15_18_port, B2 => n23, ZN => n833);
   U970 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n74_port, B1 => 
                           REGISTERS_11_18_port, B2 => n57, ZN => n832);
   U971 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n108, B1 => 
                           REGISTERS_14_18_port, B2 => n91_port, ZN => n831);
   U972 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n142_port, B1 => 
                           REGISTERS_10_18_port, B2 => n125, ZN => n830);
   U973 : NAND4_X1 port map( A1 => n833, A2 => n832, A3 => n831, A4 => n830, ZN
                           => n834);
   U974 : AOI22_X1 port map( A1 => n835, A2 => n1110, B1 => n834, B2 => n1108, 
                           ZN => n836);
   U975 : OAI221_X1 port map( B1 => n1114, B2 => n838, C1 => n1112, C2 => n837,
                           A => n836, ZN => N73);
   U976 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n40, B1 => 
                           REGISTERS_23_19_port, B2 => n23, ZN => n842);
   U977 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n74_port, B1 => 
                           REGISTERS_19_19_port, B2 => n57, ZN => n841);
   U978 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n108, B1 => 
                           REGISTERS_22_19_port, B2 => n91_port, ZN => n840);
   U979 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n142_port, B1 =>
                           REGISTERS_18_19_port, B2 => n125, ZN => n839);
   U980 : AND4_X1 port map( A1 => n842, A2 => n841, A3 => n840, A4 => n839, ZN 
                           => n859);
   U981 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n40, B1 => 
                           REGISTERS_31_19_port, B2 => n23, ZN => n846);
   U982 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n74_port, B1 => 
                           REGISTERS_27_19_port, B2 => n57, ZN => n845);
   U983 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n108, B1 => 
                           REGISTERS_30_19_port, B2 => n91_port, ZN => n844);
   U984 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n142_port, B1 =>
                           REGISTERS_26_19_port, B2 => n125, ZN => n843);
   U985 : AND4_X1 port map( A1 => n846, A2 => n845, A3 => n844, A4 => n843, ZN 
                           => n858);
   U986 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n40, B1 => 
                           REGISTERS_7_19_port, B2 => n23, ZN => n850);
   U987 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n74_port, B1 => 
                           REGISTERS_3_19_port, B2 => n57, ZN => n849);
   U988 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n108, B1 => 
                           REGISTERS_6_19_port, B2 => n91_port, ZN => n848);
   U989 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n142_port, B1 => 
                           REGISTERS_2_19_port, B2 => n125, ZN => n847);
   U990 : NAND4_X1 port map( A1 => n850, A2 => n849, A3 => n848, A4 => n847, ZN
                           => n856);
   U991 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n40, B1 => 
                           REGISTERS_15_19_port, B2 => n23, ZN => n854);
   U992 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n74_port, B1 => 
                           REGISTERS_11_19_port, B2 => n57, ZN => n853);
   U993 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n108, B1 => 
                           REGISTERS_14_19_port, B2 => n91_port, ZN => n852);
   U994 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n142_port, B1 => 
                           REGISTERS_10_19_port, B2 => n125, ZN => n851);
   U995 : NAND4_X1 port map( A1 => n854, A2 => n853, A3 => n852, A4 => n851, ZN
                           => n855);
   U996 : AOI22_X1 port map( A1 => n856, A2 => n1110, B1 => n855, B2 => n1108, 
                           ZN => n857);
   U997 : OAI221_X1 port map( B1 => n1114, B2 => n859, C1 => n1112, C2 => n858,
                           A => n857, ZN => N72);
   U998 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n40, B1 => 
                           REGISTERS_23_20_port, B2 => n23, ZN => n863);
   U999 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n74_port, B1 => 
                           REGISTERS_19_20_port, B2 => n57, ZN => n862);
   U1000 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n108, B1 => 
                           REGISTERS_22_20_port, B2 => n91_port, ZN => n861);
   U1001 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n142_port, B1 
                           => REGISTERS_18_20_port, B2 => n125, ZN => n860);
   U1002 : AND4_X1 port map( A1 => n863, A2 => n862, A3 => n861, A4 => n860, ZN
                           => n880);
   U1003 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n40, B1 => 
                           REGISTERS_31_20_port, B2 => n23, ZN => n867);
   U1004 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n74_port, B1 =>
                           REGISTERS_27_20_port, B2 => n57, ZN => n866);
   U1005 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n108, B1 => 
                           REGISTERS_30_20_port, B2 => n91_port, ZN => n865);
   U1006 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n142_port, B1 
                           => REGISTERS_26_20_port, B2 => n125, ZN => n864);
   U1007 : AND4_X1 port map( A1 => n867, A2 => n866, A3 => n865, A4 => n864, ZN
                           => n879);
   U1008 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n40, B1 => 
                           REGISTERS_7_20_port, B2 => n23, ZN => n871);
   U1009 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n74_port, B1 => 
                           REGISTERS_3_20_port, B2 => n57, ZN => n870);
   U1010 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n108, B1 => 
                           REGISTERS_6_20_port, B2 => n91_port, ZN => n869);
   U1011 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n142_port, B1 =>
                           REGISTERS_2_20_port, B2 => n125, ZN => n868);
   U1012 : NAND4_X1 port map( A1 => n871, A2 => n870, A3 => n869, A4 => n868, 
                           ZN => n877);
   U1013 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n40, B1 => 
                           REGISTERS_15_20_port, B2 => n23, ZN => n875);
   U1014 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n74_port, B1 => 
                           REGISTERS_11_20_port, B2 => n57, ZN => n874);
   U1015 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n108, B1 => 
                           REGISTERS_14_20_port, B2 => n91_port, ZN => n873);
   U1016 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n142_port, B1 =>
                           REGISTERS_10_20_port, B2 => n125, ZN => n872);
   U1017 : NAND4_X1 port map( A1 => n875, A2 => n874, A3 => n873, A4 => n872, 
                           ZN => n876);
   U1018 : AOI22_X1 port map( A1 => n877, A2 => n1110, B1 => n876, B2 => n1108,
                           ZN => n878);
   U1019 : OAI221_X1 port map( B1 => n1114, B2 => n880, C1 => n1112, C2 => n879
                           , A => n878, ZN => N71);
   U1020 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n41, B1 => 
                           REGISTERS_23_21_port, B2 => n24, ZN => n884);
   U1021 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n75_port, B1 =>
                           REGISTERS_19_21_port, B2 => n58, ZN => n883);
   U1022 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n109, B1 => 
                           REGISTERS_22_21_port, B2 => n92, ZN => n882);
   U1023 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n143_port, B1 
                           => REGISTERS_18_21_port, B2 => n126, ZN => n881);
   U1024 : AND4_X1 port map( A1 => n884, A2 => n883, A3 => n882, A4 => n881, ZN
                           => n901);
   U1025 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n41, B1 => 
                           REGISTERS_31_21_port, B2 => n24, ZN => n888);
   U1026 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n75_port, B1 =>
                           REGISTERS_27_21_port, B2 => n58, ZN => n887);
   U1027 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n109, B1 => 
                           REGISTERS_30_21_port, B2 => n92, ZN => n886);
   U1028 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n143_port, B1 
                           => REGISTERS_26_21_port, B2 => n126, ZN => n885);
   U1029 : AND4_X1 port map( A1 => n888, A2 => n887, A3 => n886, A4 => n885, ZN
                           => n900);
   U1030 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n41, B1 => 
                           REGISTERS_7_21_port, B2 => n24, ZN => n892);
   U1031 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n75_port, B1 => 
                           REGISTERS_3_21_port, B2 => n58, ZN => n891);
   U1032 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n109, B1 => 
                           REGISTERS_6_21_port, B2 => n92, ZN => n890);
   U1033 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n143_port, B1 =>
                           REGISTERS_2_21_port, B2 => n126, ZN => n889);
   U1034 : NAND4_X1 port map( A1 => n892, A2 => n891, A3 => n890, A4 => n889, 
                           ZN => n898);
   U1035 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n41, B1 => 
                           REGISTERS_15_21_port, B2 => n24, ZN => n896);
   U1036 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n75_port, B1 => 
                           REGISTERS_11_21_port, B2 => n58, ZN => n895);
   U1037 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n109, B1 => 
                           REGISTERS_14_21_port, B2 => n92, ZN => n894);
   U1038 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n143_port, B1 =>
                           REGISTERS_10_21_port, B2 => n126, ZN => n893);
   U1039 : NAND4_X1 port map( A1 => n896, A2 => n895, A3 => n894, A4 => n893, 
                           ZN => n897);
   U1040 : AOI22_X1 port map( A1 => n898, A2 => n1110, B1 => n897, B2 => n1108,
                           ZN => n899);
   U1041 : OAI221_X1 port map( B1 => n1114, B2 => n901, C1 => n1112, C2 => n900
                           , A => n899, ZN => N70);
   U1042 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n41, B1 => 
                           REGISTERS_23_22_port, B2 => n24, ZN => n905);
   U1043 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n75_port, B1 =>
                           REGISTERS_19_22_port, B2 => n58, ZN => n904);
   U1044 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n109, B1 => 
                           REGISTERS_22_22_port, B2 => n92, ZN => n903);
   U1045 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n143_port, B1 
                           => REGISTERS_18_22_port, B2 => n126, ZN => n902);
   U1046 : AND4_X1 port map( A1 => n905, A2 => n904, A3 => n903, A4 => n902, ZN
                           => n922);
   U1047 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n41, B1 => 
                           REGISTERS_31_22_port, B2 => n24, ZN => n909);
   U1048 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n75_port, B1 =>
                           REGISTERS_27_22_port, B2 => n58, ZN => n908);
   U1049 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n109, B1 => 
                           REGISTERS_30_22_port, B2 => n92, ZN => n907);
   U1050 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n143_port, B1 
                           => REGISTERS_26_22_port, B2 => n126, ZN => n906);
   U1051 : AND4_X1 port map( A1 => n909, A2 => n908, A3 => n907, A4 => n906, ZN
                           => n921);
   U1052 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n41, B1 => 
                           REGISTERS_7_22_port, B2 => n24, ZN => n913);
   U1053 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n75_port, B1 => 
                           REGISTERS_3_22_port, B2 => n58, ZN => n912);
   U1054 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n109, B1 => 
                           REGISTERS_6_22_port, B2 => n92, ZN => n911);
   U1055 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n143_port, B1 =>
                           REGISTERS_2_22_port, B2 => n126, ZN => n910);
   U1056 : NAND4_X1 port map( A1 => n913, A2 => n912, A3 => n911, A4 => n910, 
                           ZN => n919);
   U1057 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n41, B1 => 
                           REGISTERS_15_22_port, B2 => n24, ZN => n917);
   U1058 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n75_port, B1 => 
                           REGISTERS_11_22_port, B2 => n58, ZN => n916);
   U1059 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n109, B1 => 
                           REGISTERS_14_22_port, B2 => n92, ZN => n915);
   U1060 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n143_port, B1 =>
                           REGISTERS_10_22_port, B2 => n126, ZN => n914);
   U1061 : NAND4_X1 port map( A1 => n917, A2 => n916, A3 => n915, A4 => n914, 
                           ZN => n918);
   U1062 : AOI22_X1 port map( A1 => n919, A2 => n1110, B1 => n918, B2 => n1108,
                           ZN => n920);
   U1063 : OAI221_X1 port map( B1 => n1114, B2 => n922, C1 => n1112, C2 => n921
                           , A => n920, ZN => N69);
   U1064 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n41, B1 => 
                           REGISTERS_23_23_port, B2 => n24, ZN => n926);
   U1065 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n75_port, B1 =>
                           REGISTERS_19_23_port, B2 => n58, ZN => n925);
   U1066 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n109, B1 => 
                           REGISTERS_22_23_port, B2 => n92, ZN => n924);
   U1067 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n143_port, B1 
                           => REGISTERS_18_23_port, B2 => n126, ZN => n923);
   U1068 : AND4_X1 port map( A1 => n926, A2 => n925, A3 => n924, A4 => n923, ZN
                           => n943);
   U1069 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n41, B1 => 
                           REGISTERS_31_23_port, B2 => n24, ZN => n930);
   U1070 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n75_port, B1 =>
                           REGISTERS_27_23_port, B2 => n58, ZN => n929);
   U1071 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n109, B1 => 
                           REGISTERS_30_23_port, B2 => n92, ZN => n928);
   U1072 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n143_port, B1 
                           => REGISTERS_26_23_port, B2 => n126, ZN => n927);
   U1073 : AND4_X1 port map( A1 => n930, A2 => n929, A3 => n928, A4 => n927, ZN
                           => n942);
   U1074 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n41, B1 => 
                           REGISTERS_7_23_port, B2 => n24, ZN => n934);
   U1075 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n75_port, B1 => 
                           REGISTERS_3_23_port, B2 => n58, ZN => n933);
   U1076 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n109, B1 => 
                           REGISTERS_6_23_port, B2 => n92, ZN => n932);
   U1077 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n143_port, B1 =>
                           REGISTERS_2_23_port, B2 => n126, ZN => n931);
   U1078 : NAND4_X1 port map( A1 => n934, A2 => n933, A3 => n932, A4 => n931, 
                           ZN => n940);
   U1079 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n41, B1 => 
                           REGISTERS_15_23_port, B2 => n24, ZN => n938);
   U1080 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n75_port, B1 => 
                           REGISTERS_11_23_port, B2 => n58, ZN => n937);
   U1081 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n109, B1 => 
                           REGISTERS_14_23_port, B2 => n92, ZN => n936);
   U1082 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n143_port, B1 =>
                           REGISTERS_10_23_port, B2 => n126, ZN => n935);
   U1083 : NAND4_X1 port map( A1 => n938, A2 => n937, A3 => n936, A4 => n935, 
                           ZN => n939);
   U1084 : AOI22_X1 port map( A1 => n940, A2 => n1110, B1 => n939, B2 => n1108,
                           ZN => n941);
   U1085 : OAI221_X1 port map( B1 => n1114, B2 => n943, C1 => n1112, C2 => n942
                           , A => n941, ZN => N68);
   U1086 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n42, B1 => 
                           REGISTERS_23_24_port, B2 => n25, ZN => n947);
   U1087 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n76_port, B1 =>
                           REGISTERS_19_24_port, B2 => n59, ZN => n946);
   U1088 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n110, B1 => 
                           REGISTERS_22_24_port, B2 => n93, ZN => n945);
   U1089 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n144_port, B1 
                           => REGISTERS_18_24_port, B2 => n127_port, ZN => n944
                           );
   U1090 : AND4_X1 port map( A1 => n947, A2 => n946, A3 => n945, A4 => n944, ZN
                           => n964);
   U1091 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n42, B1 => 
                           REGISTERS_31_24_port, B2 => n25, ZN => n951);
   U1092 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n76_port, B1 =>
                           REGISTERS_27_24_port, B2 => n59, ZN => n950);
   U1093 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n110, B1 => 
                           REGISTERS_30_24_port, B2 => n93, ZN => n949);
   U1094 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n144_port, B1 
                           => REGISTERS_26_24_port, B2 => n127_port, ZN => n948
                           );
   U1095 : AND4_X1 port map( A1 => n951, A2 => n950, A3 => n949, A4 => n948, ZN
                           => n963);
   U1096 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n42, B1 => 
                           REGISTERS_7_24_port, B2 => n25, ZN => n955);
   U1097 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n76_port, B1 => 
                           REGISTERS_3_24_port, B2 => n59, ZN => n954);
   U1098 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n110, B1 => 
                           REGISTERS_6_24_port, B2 => n93, ZN => n953);
   U1099 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n144_port, B1 =>
                           REGISTERS_2_24_port, B2 => n127_port, ZN => n952);
   U1100 : NAND4_X1 port map( A1 => n955, A2 => n954, A3 => n953, A4 => n952, 
                           ZN => n961);
   U1101 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n42, B1 => 
                           REGISTERS_15_24_port, B2 => n25, ZN => n959);
   U1102 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n76_port, B1 => 
                           REGISTERS_11_24_port, B2 => n59, ZN => n958);
   U1103 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n110, B1 => 
                           REGISTERS_14_24_port, B2 => n93, ZN => n957);
   U1104 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n144_port, B1 =>
                           REGISTERS_10_24_port, B2 => n127_port, ZN => n956);
   U1105 : NAND4_X1 port map( A1 => n959, A2 => n958, A3 => n957, A4 => n956, 
                           ZN => n960);
   U1106 : AOI22_X1 port map( A1 => n961, A2 => n1110, B1 => n960, B2 => n1108,
                           ZN => n962);
   U1107 : OAI221_X1 port map( B1 => n1114, B2 => n964, C1 => n1112, C2 => n963
                           , A => n962, ZN => N67);
   U1108 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n42, B1 => 
                           REGISTERS_23_25_port, B2 => n25, ZN => n968);
   U1109 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n76_port, B1 =>
                           REGISTERS_19_25_port, B2 => n59, ZN => n967);
   U1110 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n110, B1 => 
                           REGISTERS_22_25_port, B2 => n93, ZN => n966);
   U1111 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n144_port, B1 
                           => REGISTERS_18_25_port, B2 => n127_port, ZN => n965
                           );
   U1112 : AND4_X1 port map( A1 => n968, A2 => n967, A3 => n966, A4 => n965, ZN
                           => n985);
   U1113 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n42, B1 => 
                           REGISTERS_31_25_port, B2 => n25, ZN => n972);
   U1114 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n76_port, B1 =>
                           REGISTERS_27_25_port, B2 => n59, ZN => n971);
   U1115 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n110, B1 => 
                           REGISTERS_30_25_port, B2 => n93, ZN => n970);
   U1116 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n144_port, B1 
                           => REGISTERS_26_25_port, B2 => n127_port, ZN => n969
                           );
   U1117 : AND4_X1 port map( A1 => n972, A2 => n971, A3 => n970, A4 => n969, ZN
                           => n984);
   U1118 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n42, B1 => 
                           REGISTERS_7_25_port, B2 => n25, ZN => n976);
   U1119 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n76_port, B1 => 
                           REGISTERS_3_25_port, B2 => n59, ZN => n975);
   U1120 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n110, B1 => 
                           REGISTERS_6_25_port, B2 => n93, ZN => n974);
   U1121 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n144_port, B1 =>
                           REGISTERS_2_25_port, B2 => n127_port, ZN => n973);
   U1122 : NAND4_X1 port map( A1 => n976, A2 => n975, A3 => n974, A4 => n973, 
                           ZN => n982);
   U1123 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n42, B1 => 
                           REGISTERS_15_25_port, B2 => n25, ZN => n980);
   U1124 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n76_port, B1 => 
                           REGISTERS_11_25_port, B2 => n59, ZN => n979);
   U1125 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n110, B1 => 
                           REGISTERS_14_25_port, B2 => n93, ZN => n978);
   U1126 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n144_port, B1 =>
                           REGISTERS_10_25_port, B2 => n127_port, ZN => n977);
   U1127 : NAND4_X1 port map( A1 => n980, A2 => n979, A3 => n978, A4 => n977, 
                           ZN => n981);
   U1128 : AOI22_X1 port map( A1 => n982, A2 => n1110, B1 => n981, B2 => n1108,
                           ZN => n983);
   U1129 : OAI221_X1 port map( B1 => n1114, B2 => n985, C1 => n1112, C2 => n984
                           , A => n983, ZN => N66);
   U1130 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n42, B1 => 
                           REGISTERS_23_26_port, B2 => n25, ZN => n989);
   U1131 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n76_port, B1 =>
                           REGISTERS_19_26_port, B2 => n59, ZN => n988);
   U1132 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n110, B1 => 
                           REGISTERS_22_26_port, B2 => n93, ZN => n987);
   U1133 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n144_port, B1 
                           => REGISTERS_18_26_port, B2 => n127_port, ZN => n986
                           );
   U1134 : AND4_X1 port map( A1 => n989, A2 => n988, A3 => n987, A4 => n986, ZN
                           => n1006);
   U1135 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n42, B1 => 
                           REGISTERS_31_26_port, B2 => n25, ZN => n993);
   U1136 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n76_port, B1 =>
                           REGISTERS_27_26_port, B2 => n59, ZN => n992);
   U1137 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n110, B1 => 
                           REGISTERS_30_26_port, B2 => n93, ZN => n991);
   U1138 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n144_port, B1 
                           => REGISTERS_26_26_port, B2 => n127_port, ZN => n990
                           );
   U1139 : AND4_X1 port map( A1 => n993, A2 => n992, A3 => n991, A4 => n990, ZN
                           => n1005);
   U1140 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n42, B1 => 
                           REGISTERS_7_26_port, B2 => n25, ZN => n997);
   U1141 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n76_port, B1 => 
                           REGISTERS_3_26_port, B2 => n59, ZN => n996);
   U1142 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n110, B1 => 
                           REGISTERS_6_26_port, B2 => n93, ZN => n995);
   U1143 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n144_port, B1 =>
                           REGISTERS_2_26_port, B2 => n127_port, ZN => n994);
   U1144 : NAND4_X1 port map( A1 => n997, A2 => n996, A3 => n995, A4 => n994, 
                           ZN => n1003);
   U1145 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n42, B1 => 
                           REGISTERS_15_26_port, B2 => n25, ZN => n1001);
   U1146 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n76_port, B1 => 
                           REGISTERS_11_26_port, B2 => n59, ZN => n1000);
   U1147 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n110, B1 => 
                           REGISTERS_14_26_port, B2 => n93, ZN => n999);
   U1148 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n144_port, B1 =>
                           REGISTERS_10_26_port, B2 => n127_port, ZN => n998);
   U1149 : NAND4_X1 port map( A1 => n1001, A2 => n1000, A3 => n999, A4 => n998,
                           ZN => n1002);
   U1150 : AOI22_X1 port map( A1 => n1003, A2 => n1110, B1 => n1002, B2 => 
                           n1108, ZN => n1004);
   U1151 : OAI221_X1 port map( B1 => n1114, B2 => n1006, C1 => n1112, C2 => 
                           n1005, A => n1004, ZN => N65);
   U1152 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n43, B1 => 
                           REGISTERS_23_27_port, B2 => n26, ZN => n1010);
   U1153 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n77_port, B1 =>
                           REGISTERS_19_27_port, B2 => n60_port, ZN => n1009);
   U1154 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n111, B1 => 
                           REGISTERS_22_27_port, B2 => n94, ZN => n1008);
   U1155 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n145_port, B1 
                           => REGISTERS_18_27_port, B2 => n128_port, ZN => 
                           n1007);
   U1156 : AND4_X1 port map( A1 => n1010, A2 => n1009, A3 => n1008, A4 => n1007
                           , ZN => n1027);
   U1157 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n43, B1 => 
                           REGISTERS_31_27_port, B2 => n26, ZN => n1014);
   U1158 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n77_port, B1 =>
                           REGISTERS_27_27_port, B2 => n60_port, ZN => n1013);
   U1159 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n111, B1 => 
                           REGISTERS_30_27_port, B2 => n94, ZN => n1012);
   U1160 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n145_port, B1 
                           => REGISTERS_26_27_port, B2 => n128_port, ZN => 
                           n1011);
   U1161 : AND4_X1 port map( A1 => n1014, A2 => n1013, A3 => n1012, A4 => n1011
                           , ZN => n1026);
   U1162 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n43, B1 => 
                           REGISTERS_7_27_port, B2 => n26, ZN => n1018);
   U1163 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n77_port, B1 => 
                           REGISTERS_3_27_port, B2 => n60_port, ZN => n1017);
   U1164 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n111, B1 => 
                           REGISTERS_6_27_port, B2 => n94, ZN => n1016);
   U1165 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n145_port, B1 =>
                           REGISTERS_2_27_port, B2 => n128_port, ZN => n1015);
   U1166 : NAND4_X1 port map( A1 => n1018, A2 => n1017, A3 => n1016, A4 => 
                           n1015, ZN => n1024);
   U1167 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n43, B1 => 
                           REGISTERS_15_27_port, B2 => n26, ZN => n1022);
   U1168 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n77_port, B1 => 
                           REGISTERS_11_27_port, B2 => n60_port, ZN => n1021);
   U1169 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n111, B1 => 
                           REGISTERS_14_27_port, B2 => n94, ZN => n1020);
   U1170 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n145_port, B1 =>
                           REGISTERS_10_27_port, B2 => n128_port, ZN => n1019);
   U1171 : NAND4_X1 port map( A1 => n1022, A2 => n1021, A3 => n1020, A4 => 
                           n1019, ZN => n1023);
   U1172 : AOI22_X1 port map( A1 => n1024, A2 => n1110, B1 => n1023, B2 => 
                           n1108, ZN => n1025);
   U1173 : OAI221_X1 port map( B1 => n1114, B2 => n1027, C1 => n1112, C2 => 
                           n1026, A => n1025, ZN => N64);
   U1174 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n43, B1 => 
                           REGISTERS_23_28_port, B2 => n26, ZN => n1031);
   U1175 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n77_port, B1 =>
                           REGISTERS_19_28_port, B2 => n60_port, ZN => n1030);
   U1176 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n111, B1 => 
                           REGISTERS_22_28_port, B2 => n94, ZN => n1029);
   U1177 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n145_port, B1 
                           => REGISTERS_18_28_port, B2 => n128_port, ZN => 
                           n1028);
   U1178 : AND4_X1 port map( A1 => n1031, A2 => n1030, A3 => n1029, A4 => n1028
                           , ZN => n1048);
   U1179 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n43, B1 => 
                           REGISTERS_31_28_port, B2 => n26, ZN => n1035);
   U1180 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n77_port, B1 =>
                           REGISTERS_27_28_port, B2 => n60_port, ZN => n1034);
   U1181 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n111, B1 => 
                           REGISTERS_30_28_port, B2 => n94, ZN => n1033);
   U1182 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n145_port, B1 
                           => REGISTERS_26_28_port, B2 => n128_port, ZN => 
                           n1032);
   U1183 : AND4_X1 port map( A1 => n1035, A2 => n1034, A3 => n1033, A4 => n1032
                           , ZN => n1047);
   U1184 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n43, B1 => 
                           REGISTERS_7_28_port, B2 => n26, ZN => n1039);
   U1185 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n77_port, B1 => 
                           REGISTERS_3_28_port, B2 => n60_port, ZN => n1038);
   U1186 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n111, B1 => 
                           REGISTERS_6_28_port, B2 => n94, ZN => n1037);
   U1187 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n145_port, B1 =>
                           REGISTERS_2_28_port, B2 => n128_port, ZN => n1036);
   U1188 : NAND4_X1 port map( A1 => n1039, A2 => n1038, A3 => n1037, A4 => 
                           n1036, ZN => n1045);
   U1189 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n43, B1 => 
                           REGISTERS_15_28_port, B2 => n26, ZN => n1043);
   U1190 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n77_port, B1 => 
                           REGISTERS_11_28_port, B2 => n60_port, ZN => n1042);
   U1191 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n111, B1 => 
                           REGISTERS_14_28_port, B2 => n94, ZN => n1041);
   U1192 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n145_port, B1 =>
                           REGISTERS_10_28_port, B2 => n128_port, ZN => n1040);
   U1193 : NAND4_X1 port map( A1 => n1043, A2 => n1042, A3 => n1041, A4 => 
                           n1040, ZN => n1044);
   U1194 : AOI22_X1 port map( A1 => n1045, A2 => n1110, B1 => n1044, B2 => 
                           n1108, ZN => n1046);
   U1195 : OAI221_X1 port map( B1 => n1114, B2 => n1048, C1 => n1112, C2 => 
                           n1047, A => n1046, ZN => N63);
   U1196 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n43, B1 => 
                           REGISTERS_23_29_port, B2 => n26, ZN => n1052);
   U1197 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n77_port, B1 =>
                           REGISTERS_19_29_port, B2 => n60_port, ZN => n1051);
   U1198 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n111, B1 => 
                           REGISTERS_22_29_port, B2 => n94, ZN => n1050);
   U1199 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n145_port, B1 
                           => REGISTERS_18_29_port, B2 => n128_port, ZN => 
                           n1049);
   U1200 : AND4_X1 port map( A1 => n1052, A2 => n1051, A3 => n1050, A4 => n1049
                           , ZN => n1069);
   U1201 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n43, B1 => 
                           REGISTERS_31_29_port, B2 => n26, ZN => n1056);
   U1202 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n77_port, B1 =>
                           REGISTERS_27_29_port, B2 => n60_port, ZN => n1055);
   U1203 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n111, B1 => 
                           REGISTERS_30_29_port, B2 => n94, ZN => n1054);
   U1204 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n145_port, B1 
                           => REGISTERS_26_29_port, B2 => n128_port, ZN => 
                           n1053);
   U1205 : AND4_X1 port map( A1 => n1056, A2 => n1055, A3 => n1054, A4 => n1053
                           , ZN => n1068);
   U1206 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n43, B1 => 
                           REGISTERS_7_29_port, B2 => n26, ZN => n1060);
   U1207 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n77_port, B1 => 
                           REGISTERS_3_29_port, B2 => n60_port, ZN => n1059);
   U1208 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n111, B1 => 
                           REGISTERS_6_29_port, B2 => n94, ZN => n1058);
   U1209 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n145_port, B1 =>
                           REGISTERS_2_29_port, B2 => n128_port, ZN => n1057);
   U1210 : NAND4_X1 port map( A1 => n1060, A2 => n1059, A3 => n1058, A4 => 
                           n1057, ZN => n1066);
   U1211 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n43, B1 => 
                           REGISTERS_15_29_port, B2 => n26, ZN => n1064);
   U1212 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n77_port, B1 => 
                           REGISTERS_11_29_port, B2 => n60_port, ZN => n1063);
   U1213 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n111, B1 => 
                           REGISTERS_14_29_port, B2 => n94, ZN => n1062);
   U1214 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n145_port, B1 =>
                           REGISTERS_10_29_port, B2 => n128_port, ZN => n1061);
   U1215 : NAND4_X1 port map( A1 => n1064, A2 => n1063, A3 => n1062, A4 => 
                           n1061, ZN => n1065);
   U1216 : AOI22_X1 port map( A1 => n1066, A2 => n1110, B1 => n1065, B2 => 
                           n1108, ZN => n1067);
   U1217 : OAI221_X1 port map( B1 => n1114, B2 => n1069, C1 => n1112, C2 => 
                           n1068, A => n1067, ZN => N62);
   U1218 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n44, B1 => 
                           REGISTERS_23_30_port, B2 => n27, ZN => n1073);
   U1219 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n78_port, B1 =>
                           REGISTERS_19_30_port, B2 => n61_port, ZN => n1072);
   U1220 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n112, B1 => 
                           REGISTERS_22_30_port, B2 => n95, ZN => n1071);
   U1221 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n146_port, B1 
                           => REGISTERS_18_30_port, B2 => n129_port, ZN => 
                           n1070);
   U1222 : AND4_X1 port map( A1 => n1073, A2 => n1072, A3 => n1071, A4 => n1070
                           , ZN => n1090);
   U1223 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n44, B1 => 
                           REGISTERS_31_30_port, B2 => n27, ZN => n1077);
   U1224 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n78_port, B1 =>
                           REGISTERS_27_30_port, B2 => n61_port, ZN => n1076);
   U1225 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n112, B1 => 
                           REGISTERS_30_30_port, B2 => n95, ZN => n1075);
   U1226 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n146_port, B1 
                           => REGISTERS_26_30_port, B2 => n129_port, ZN => 
                           n1074);
   U1227 : AND4_X1 port map( A1 => n1077, A2 => n1076, A3 => n1075, A4 => n1074
                           , ZN => n1089);
   U1228 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n44, B1 => 
                           REGISTERS_7_30_port, B2 => n27, ZN => n1081);
   U1229 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n78_port, B1 => 
                           REGISTERS_3_30_port, B2 => n61_port, ZN => n1080);
   U1230 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n112, B1 => 
                           REGISTERS_6_30_port, B2 => n95, ZN => n1079);
   U1231 : AOI22_X1 port map( A1 => REGISTERS_0_30_port, A2 => n146_port, B1 =>
                           REGISTERS_2_30_port, B2 => n129_port, ZN => n1078);
   U1232 : NAND4_X1 port map( A1 => n1081, A2 => n1080, A3 => n1079, A4 => 
                           n1078, ZN => n1087);
   U1233 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n44, B1 => 
                           REGISTERS_15_30_port, B2 => n27, ZN => n1085);
   U1234 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n78_port, B1 => 
                           REGISTERS_11_30_port, B2 => n61_port, ZN => n1084);
   U1235 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n112, B1 => 
                           REGISTERS_14_30_port, B2 => n95, ZN => n1083);
   U1236 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n146_port, B1 =>
                           REGISTERS_10_30_port, B2 => n129_port, ZN => n1082);
   U1237 : NAND4_X1 port map( A1 => n1085, A2 => n1084, A3 => n1083, A4 => 
                           n1082, ZN => n1086);
   U1238 : AOI22_X1 port map( A1 => n1087, A2 => n1110, B1 => n1086, B2 => 
                           n1108, ZN => n1088);
   U1239 : OAI221_X1 port map( B1 => n1114, B2 => n1090, C1 => n1112, C2 => 
                           n1089, A => n1088, ZN => N61);
   U1240 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n44, B1 => 
                           REGISTERS_23_31_port, B2 => n27, ZN => n1094);
   U1241 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n78_port, B1 =>
                           REGISTERS_19_31_port, B2 => n61_port, ZN => n1093);
   U1242 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n112, B1 => 
                           REGISTERS_22_31_port, B2 => n95, ZN => n1092);
   U1243 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n146_port, B1 
                           => REGISTERS_18_31_port, B2 => n129_port, ZN => 
                           n1091);
   U1244 : AND4_X1 port map( A1 => n1094, A2 => n1093, A3 => n1092, A4 => n1091
                           , ZN => n1115);
   U1245 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n44, B1 => 
                           REGISTERS_31_31_port, B2 => n27, ZN => n1098);
   U1246 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n78_port, B1 =>
                           REGISTERS_27_31_port, B2 => n61_port, ZN => n1097);
   U1247 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n112, B1 => 
                           REGISTERS_30_31_port, B2 => n95, ZN => n1096);
   U1248 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n146_port, B1 
                           => REGISTERS_26_31_port, B2 => n129_port, ZN => 
                           n1095);
   U1249 : AND4_X1 port map( A1 => n1098, A2 => n1097, A3 => n1096, A4 => n1095
                           , ZN => n1113);
   U1250 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n44, B1 => 
                           REGISTERS_7_31_port, B2 => n27, ZN => n1102);
   U1251 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n78_port, B1 => 
                           REGISTERS_3_31_port, B2 => n61_port, ZN => n1101);
   U1252 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n112, B1 => 
                           REGISTERS_6_31_port, B2 => n95, ZN => n1100);
   U1253 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n146_port, B1 =>
                           REGISTERS_2_31_port, B2 => n129_port, ZN => n1099);
   U1254 : NAND4_X1 port map( A1 => n1102, A2 => n1101, A3 => n1100, A4 => 
                           n1099, ZN => n1109);
   U1255 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n44, B1 => 
                           REGISTERS_15_31_port, B2 => n27, ZN => n1106);
   U1256 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n78_port, B1 => 
                           REGISTERS_11_31_port, B2 => n61_port, ZN => n1105);
   U1257 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n112, B1 => 
                           REGISTERS_14_31_port, B2 => n95, ZN => n1104);
   U1258 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n146_port, B1 =>
                           REGISTERS_10_31_port, B2 => n129_port, ZN => n1103);
   U1259 : NAND4_X1 port map( A1 => n1106, A2 => n1105, A3 => n1104, A4 => 
                           n1103, ZN => n1107);
   U1260 : AOI22_X1 port map( A1 => n1110, A2 => n1109, B1 => n1108, B2 => 
                           n1107, ZN => n1111);
   U1261 : OAI221_X1 port map( B1 => n1115, B2 => n1114, C1 => n1113, C2 => 
                           n1112, A => n1111, ZN => N60);
   U1262 : NOR2_X1 port map( A1 => n2825, A2 => ADD_RD2(1), ZN => n1120);
   U1263 : NOR2_X1 port map( A1 => n2825, A2 => n2826, ZN => n1121);
   U1264 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n170, B1 => 
                           REGISTERS_23_0_port, B2 => n153_port, ZN => n1127);
   U1265 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1122);
   U1266 : NOR2_X1 port map( A1 => n2826, A2 => ADD_RD2(2), ZN => n1123);
   U1267 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n204, B1 => 
                           REGISTERS_19_0_port, B2 => n187, ZN => n1126);
   U1268 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n238, B1 => 
                           REGISTERS_22_0_port, B2 => n221, ZN => n1125);
   U1269 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n272, B1 => 
                           REGISTERS_18_0_port, B2 => n255, ZN => n1124);
   U1270 : AND4_X1 port map( A1 => n1127, A2 => n1126, A3 => n1125, A4 => n1124
                           , ZN => n1144);
   U1271 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n170, B1 => 
                           REGISTERS_31_0_port, B2 => n153_port, ZN => n1131);
   U1272 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n204, B1 => 
                           REGISTERS_27_0_port, B2 => n187, ZN => n1130);
   U1273 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n238, B1 => 
                           REGISTERS_30_0_port, B2 => n221, ZN => n1129);
   U1274 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n272, B1 => 
                           REGISTERS_26_0_port, B2 => n255, ZN => n1128);
   U1275 : AND4_X1 port map( A1 => n1131, A2 => n1130, A3 => n1129, A4 => n1128
                           , ZN => n1143);
   U1276 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n170, B1 => 
                           REGISTERS_7_0_port, B2 => n153_port, ZN => n1135);
   U1277 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n204, B1 => 
                           REGISTERS_3_0_port, B2 => n187, ZN => n1134);
   U1278 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n238, B1 => 
                           REGISTERS_6_0_port, B2 => n221, ZN => n1133);
   U1279 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n272, B1 => 
                           REGISTERS_2_0_port, B2 => n255, ZN => n1132);
   U1280 : NAND4_X1 port map( A1 => n1135, A2 => n1134, A3 => n1133, A4 => 
                           n1132, ZN => n1141);
   U1281 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n170, B1 => 
                           REGISTERS_15_0_port, B2 => n153_port, ZN => n1139);
   U1282 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n204, B1 => 
                           REGISTERS_11_0_port, B2 => n187, ZN => n1138);
   U1283 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n238, B1 => 
                           REGISTERS_14_0_port, B2 => n221, ZN => n1137);
   U1284 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n272, B1 => 
                           REGISTERS_10_0_port, B2 => n255, ZN => n1136);
   U1285 : NAND4_X1 port map( A1 => n1139, A2 => n1138, A3 => n1137, A4 => 
                           n1136, ZN => n1140);
   U1286 : AOI22_X1 port map( A1 => n1141, A2 => n2818, B1 => n1140, B2 => 
                           n2816, ZN => n1142);
   U1287 : OAI221_X1 port map( B1 => n2822, B2 => n1144, C1 => n2820, C2 => 
                           n1143, A => n1142, ZN => N158);
   U1288 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n170, B1 => 
                           REGISTERS_23_1_port, B2 => n153_port, ZN => n1148);
   U1289 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n204, B1 => 
                           REGISTERS_19_1_port, B2 => n187, ZN => n1147);
   U1290 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n238, B1 => 
                           REGISTERS_22_1_port, B2 => n221, ZN => n1146);
   U1291 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n272, B1 => 
                           REGISTERS_18_1_port, B2 => n255, ZN => n1145);
   U1292 : AND4_X1 port map( A1 => n1148, A2 => n1147, A3 => n1146, A4 => n1145
                           , ZN => n1165);
   U1293 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n170, B1 => 
                           REGISTERS_31_1_port, B2 => n153_port, ZN => n1152);
   U1294 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n204, B1 => 
                           REGISTERS_27_1_port, B2 => n187, ZN => n1151);
   U1295 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n238, B1 => 
                           REGISTERS_30_1_port, B2 => n221, ZN => n1150);
   U1296 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n272, B1 => 
                           REGISTERS_26_1_port, B2 => n255, ZN => n1149);
   U1297 : AND4_X1 port map( A1 => n1152, A2 => n1151, A3 => n1150, A4 => n1149
                           , ZN => n1164);
   U1298 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n170, B1 => 
                           REGISTERS_7_1_port, B2 => n153_port, ZN => n1156);
   U1299 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n204, B1 => 
                           REGISTERS_3_1_port, B2 => n187, ZN => n1155);
   U1300 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n238, B1 => 
                           REGISTERS_6_1_port, B2 => n221, ZN => n1154);
   U1301 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n272, B1 => 
                           REGISTERS_2_1_port, B2 => n255, ZN => n1153);
   U1302 : NAND4_X1 port map( A1 => n1156, A2 => n1155, A3 => n1154, A4 => 
                           n1153, ZN => n1162);
   U1303 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n170, B1 => 
                           REGISTERS_15_1_port, B2 => n153_port, ZN => n1160);
   U1304 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n204, B1 => 
                           REGISTERS_11_1_port, B2 => n187, ZN => n1159);
   U1305 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n238, B1 => 
                           REGISTERS_14_1_port, B2 => n221, ZN => n1158);
   U1306 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n272, B1 => 
                           REGISTERS_10_1_port, B2 => n255, ZN => n1157);
   U1307 : NAND4_X1 port map( A1 => n1160, A2 => n1159, A3 => n1158, A4 => 
                           n1157, ZN => n1161);
   U1308 : AOI22_X1 port map( A1 => n1162, A2 => n2818, B1 => n1161, B2 => 
                           n2816, ZN => n1163);
   U1309 : OAI221_X1 port map( B1 => n2822, B2 => n1165, C1 => n2820, C2 => 
                           n1164, A => n1163, ZN => N157);
   U1310 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n170, B1 => 
                           REGISTERS_23_2_port, B2 => n153_port, ZN => n1169);
   U1311 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n204, B1 => 
                           REGISTERS_19_2_port, B2 => n187, ZN => n1168);
   U1312 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n238, B1 => 
                           REGISTERS_22_2_port, B2 => n221, ZN => n1167);
   U1313 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n272, B1 => 
                           REGISTERS_18_2_port, B2 => n255, ZN => n1166);
   U1314 : AND4_X1 port map( A1 => n1169, A2 => n1168, A3 => n1167, A4 => n1166
                           , ZN => n1186);
   U1315 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n170, B1 => 
                           REGISTERS_31_2_port, B2 => n153_port, ZN => n1173);
   U1316 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n204, B1 => 
                           REGISTERS_27_2_port, B2 => n187, ZN => n1172);
   U1317 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n238, B1 => 
                           REGISTERS_30_2_port, B2 => n221, ZN => n1171);
   U1318 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n272, B1 => 
                           REGISTERS_26_2_port, B2 => n255, ZN => n1170);
   U1319 : AND4_X1 port map( A1 => n1173, A2 => n1172, A3 => n1171, A4 => n1170
                           , ZN => n1185);
   U1320 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n170, B1 => 
                           REGISTERS_7_2_port, B2 => n153_port, ZN => n1177);
   U1321 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n204, B1 => 
                           REGISTERS_3_2_port, B2 => n187, ZN => n1176);
   U1322 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n238, B1 => 
                           REGISTERS_6_2_port, B2 => n221, ZN => n1175);
   U1323 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n272, B1 => 
                           REGISTERS_2_2_port, B2 => n255, ZN => n1174);
   U1324 : NAND4_X1 port map( A1 => n1177, A2 => n1176, A3 => n1175, A4 => 
                           n1174, ZN => n1183);
   U1325 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n170, B1 => 
                           REGISTERS_15_2_port, B2 => n153_port, ZN => n1181);
   U1326 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n204, B1 => 
                           REGISTERS_11_2_port, B2 => n187, ZN => n1180);
   U1327 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n238, B1 => 
                           REGISTERS_14_2_port, B2 => n221, ZN => n1179);
   U1328 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n272, B1 => 
                           REGISTERS_10_2_port, B2 => n255, ZN => n1178);
   U1329 : NAND4_X1 port map( A1 => n1181, A2 => n1180, A3 => n1179, A4 => 
                           n1178, ZN => n1182);
   U1330 : AOI22_X1 port map( A1 => n1183, A2 => n2818, B1 => n1182, B2 => 
                           n2816, ZN => n1184);
   U1331 : OAI221_X1 port map( B1 => n2822, B2 => n1186, C1 => n2820, C2 => 
                           n1185, A => n1184, ZN => N156);
   U1332 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n171, B1 => 
                           REGISTERS_23_3_port, B2 => n154_port, ZN => n1190);
   U1333 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n205, B1 => 
                           REGISTERS_19_3_port, B2 => n188, ZN => n1189);
   U1334 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n239, B1 => 
                           REGISTERS_22_3_port, B2 => n222, ZN => n1188);
   U1335 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n273, B1 => 
                           REGISTERS_18_3_port, B2 => n256, ZN => n1187);
   U1336 : AND4_X1 port map( A1 => n1190, A2 => n1189, A3 => n1188, A4 => n1187
                           , ZN => n1207);
   U1337 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n171, B1 => 
                           REGISTERS_31_3_port, B2 => n154_port, ZN => n1194);
   U1338 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n205, B1 => 
                           REGISTERS_27_3_port, B2 => n188, ZN => n1193);
   U1339 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n239, B1 => 
                           REGISTERS_30_3_port, B2 => n222, ZN => n1192);
   U1340 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n273, B1 => 
                           REGISTERS_26_3_port, B2 => n256, ZN => n1191);
   U1341 : AND4_X1 port map( A1 => n1194, A2 => n1193, A3 => n1192, A4 => n1191
                           , ZN => n1206);
   U1342 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n171, B1 => 
                           REGISTERS_7_3_port, B2 => n154_port, ZN => n1198);
   U1343 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n205, B1 => 
                           REGISTERS_3_3_port, B2 => n188, ZN => n1197);
   U1344 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n239, B1 => 
                           REGISTERS_6_3_port, B2 => n222, ZN => n1196);
   U1345 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n273, B1 => 
                           REGISTERS_2_3_port, B2 => n256, ZN => n1195);
   U1346 : NAND4_X1 port map( A1 => n1198, A2 => n1197, A3 => n1196, A4 => 
                           n1195, ZN => n1204);
   U1347 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n171, B1 => 
                           REGISTERS_15_3_port, B2 => n154_port, ZN => n1202);
   U1348 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n205, B1 => 
                           REGISTERS_11_3_port, B2 => n188, ZN => n1201);
   U1349 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n239, B1 => 
                           REGISTERS_14_3_port, B2 => n222, ZN => n1200);
   U1350 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n273, B1 => 
                           REGISTERS_10_3_port, B2 => n256, ZN => n1199);
   U1351 : NAND4_X1 port map( A1 => n1202, A2 => n1201, A3 => n1200, A4 => 
                           n1199, ZN => n1203);
   U1352 : AOI22_X1 port map( A1 => n1204, A2 => n2818, B1 => n1203, B2 => 
                           n2816, ZN => n1205);
   U1353 : OAI221_X1 port map( B1 => n2822, B2 => n1207, C1 => n2820, C2 => 
                           n1206, A => n1205, ZN => N155);
   U1354 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n171, B1 => 
                           REGISTERS_23_4_port, B2 => n154_port, ZN => n1211);
   U1355 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n205, B1 => 
                           REGISTERS_19_4_port, B2 => n188, ZN => n1210);
   U1356 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n239, B1 => 
                           REGISTERS_22_4_port, B2 => n222, ZN => n1209);
   U1357 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n273, B1 => 
                           REGISTERS_18_4_port, B2 => n256, ZN => n1208);
   U1358 : AND4_X1 port map( A1 => n1211, A2 => n1210, A3 => n1209, A4 => n1208
                           , ZN => n1228);
   U1359 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n171, B1 => 
                           REGISTERS_31_4_port, B2 => n154_port, ZN => n1215);
   U1360 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n205, B1 => 
                           REGISTERS_27_4_port, B2 => n188, ZN => n1214);
   U1361 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n239, B1 => 
                           REGISTERS_30_4_port, B2 => n222, ZN => n1213);
   U1362 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n273, B1 => 
                           REGISTERS_26_4_port, B2 => n256, ZN => n1212);
   U1363 : AND4_X1 port map( A1 => n1215, A2 => n1214, A3 => n1213, A4 => n1212
                           , ZN => n1227);
   U1364 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n171, B1 => 
                           REGISTERS_7_4_port, B2 => n154_port, ZN => n1219);
   U1365 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n205, B1 => 
                           REGISTERS_3_4_port, B2 => n188, ZN => n1218);
   U1366 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n239, B1 => 
                           REGISTERS_6_4_port, B2 => n222, ZN => n1217);
   U1367 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n273, B1 => 
                           REGISTERS_2_4_port, B2 => n256, ZN => n1216);
   U1368 : NAND4_X1 port map( A1 => n1219, A2 => n1218, A3 => n1217, A4 => 
                           n1216, ZN => n1225);
   U1369 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n171, B1 => 
                           REGISTERS_15_4_port, B2 => n154_port, ZN => n1223);
   U1370 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n205, B1 => 
                           REGISTERS_11_4_port, B2 => n188, ZN => n1222);
   U1371 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n239, B1 => 
                           REGISTERS_14_4_port, B2 => n222, ZN => n1221);
   U1372 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n273, B1 => 
                           REGISTERS_10_4_port, B2 => n256, ZN => n1220);
   U1373 : NAND4_X1 port map( A1 => n1223, A2 => n1222, A3 => n1221, A4 => 
                           n1220, ZN => n1224);
   U1374 : AOI22_X1 port map( A1 => n1225, A2 => n2818, B1 => n1224, B2 => 
                           n2816, ZN => n1226);
   U1375 : OAI221_X1 port map( B1 => n2822, B2 => n1228, C1 => n2820, C2 => 
                           n1227, A => n1226, ZN => N154);
   U1376 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n171, B1 => 
                           REGISTERS_23_5_port, B2 => n154_port, ZN => n1232);
   U1377 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n205, B1 => 
                           REGISTERS_19_5_port, B2 => n188, ZN => n1231);
   U1378 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n239, B1 => 
                           REGISTERS_22_5_port, B2 => n222, ZN => n1230);
   U1379 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n273, B1 => 
                           REGISTERS_18_5_port, B2 => n256, ZN => n1229);
   U1380 : AND4_X1 port map( A1 => n1232, A2 => n1231, A3 => n1230, A4 => n1229
                           , ZN => n1249);
   U1381 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n171, B1 => 
                           REGISTERS_31_5_port, B2 => n154_port, ZN => n1236);
   U1382 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n205, B1 => 
                           REGISTERS_27_5_port, B2 => n188, ZN => n1235);
   U1383 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n239, B1 => 
                           REGISTERS_30_5_port, B2 => n222, ZN => n1234);
   U1384 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n273, B1 => 
                           REGISTERS_26_5_port, B2 => n256, ZN => n1233);
   U1385 : AND4_X1 port map( A1 => n1236, A2 => n1235, A3 => n1234, A4 => n1233
                           , ZN => n1248);
   U1386 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n171, B1 => 
                           REGISTERS_7_5_port, B2 => n154_port, ZN => n1240);
   U1387 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n205, B1 => 
                           REGISTERS_3_5_port, B2 => n188, ZN => n1239);
   U1388 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n239, B1 => 
                           REGISTERS_6_5_port, B2 => n222, ZN => n1238);
   U1389 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n273, B1 => 
                           REGISTERS_2_5_port, B2 => n256, ZN => n1237);
   U1390 : NAND4_X1 port map( A1 => n1240, A2 => n1239, A3 => n1238, A4 => 
                           n1237, ZN => n1246);
   U1391 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n171, B1 => 
                           REGISTERS_15_5_port, B2 => n154_port, ZN => n1244);
   U1392 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n205, B1 => 
                           REGISTERS_11_5_port, B2 => n188, ZN => n1243);
   U1393 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n239, B1 => 
                           REGISTERS_14_5_port, B2 => n222, ZN => n1242);
   U1394 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n273, B1 => 
                           REGISTERS_10_5_port, B2 => n256, ZN => n1241);
   U1395 : NAND4_X1 port map( A1 => n1244, A2 => n1243, A3 => n1242, A4 => 
                           n1241, ZN => n1245);
   U1396 : AOI22_X1 port map( A1 => n1246, A2 => n2818, B1 => n1245, B2 => 
                           n2816, ZN => n1247);
   U1397 : OAI221_X1 port map( B1 => n2822, B2 => n1249, C1 => n2820, C2 => 
                           n1248, A => n1247, ZN => N153);
   U1398 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n172, B1 => 
                           REGISTERS_23_6_port, B2 => n155_port, ZN => n1253);
   U1399 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n206, B1 => 
                           REGISTERS_19_6_port, B2 => n189, ZN => n1252);
   U1400 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n240, B1 => 
                           REGISTERS_22_6_port, B2 => n223, ZN => n1251);
   U1401 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n274, B1 => 
                           REGISTERS_18_6_port, B2 => n257, ZN => n1250);
   U1402 : AND4_X1 port map( A1 => n1253, A2 => n1252, A3 => n1251, A4 => n1250
                           , ZN => n1270);
   U1403 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n172, B1 => 
                           REGISTERS_31_6_port, B2 => n155_port, ZN => n1257);
   U1404 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n206, B1 => 
                           REGISTERS_27_6_port, B2 => n189, ZN => n1256);
   U1405 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n240, B1 => 
                           REGISTERS_30_6_port, B2 => n223, ZN => n1255);
   U1406 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n274, B1 => 
                           REGISTERS_26_6_port, B2 => n257, ZN => n1254);
   U1407 : AND4_X1 port map( A1 => n1257, A2 => n1256, A3 => n1255, A4 => n1254
                           , ZN => n1269);
   U1408 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n172, B1 => 
                           REGISTERS_7_6_port, B2 => n155_port, ZN => n1261);
   U1409 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n206, B1 => 
                           REGISTERS_3_6_port, B2 => n189, ZN => n1260);
   U1410 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n240, B1 => 
                           REGISTERS_6_6_port, B2 => n223, ZN => n1259);
   U1411 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n274, B1 => 
                           REGISTERS_2_6_port, B2 => n257, ZN => n1258);
   U1412 : NAND4_X1 port map( A1 => n1261, A2 => n1260, A3 => n1259, A4 => 
                           n1258, ZN => n1267);
   U1413 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n172, B1 => 
                           REGISTERS_15_6_port, B2 => n155_port, ZN => n1265);
   U1414 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n206, B1 => 
                           REGISTERS_11_6_port, B2 => n189, ZN => n1264);
   U1415 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n240, B1 => 
                           REGISTERS_14_6_port, B2 => n223, ZN => n1263);
   U1416 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n274, B1 => 
                           REGISTERS_10_6_port, B2 => n257, ZN => n1262);
   U1417 : NAND4_X1 port map( A1 => n1265, A2 => n1264, A3 => n1263, A4 => 
                           n1262, ZN => n1266);
   U1418 : AOI22_X1 port map( A1 => n1267, A2 => n2818, B1 => n1266, B2 => 
                           n2816, ZN => n1268);
   U1419 : OAI221_X1 port map( B1 => n2822, B2 => n1270, C1 => n2820, C2 => 
                           n1269, A => n1268, ZN => N152);
   U1420 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n172, B1 => 
                           REGISTERS_23_7_port, B2 => n155_port, ZN => n1274);
   U1421 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n206, B1 => 
                           REGISTERS_19_7_port, B2 => n189, ZN => n1273);
   U1422 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n240, B1 => 
                           REGISTERS_22_7_port, B2 => n223, ZN => n1272);
   U1423 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n274, B1 => 
                           REGISTERS_18_7_port, B2 => n257, ZN => n1271);
   U1424 : AND4_X1 port map( A1 => n1274, A2 => n1273, A3 => n1272, A4 => n1271
                           , ZN => n1291);
   U1425 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n172, B1 => 
                           REGISTERS_31_7_port, B2 => n155_port, ZN => n1278);
   U1426 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n206, B1 => 
                           REGISTERS_27_7_port, B2 => n189, ZN => n1277);
   U1427 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n240, B1 => 
                           REGISTERS_30_7_port, B2 => n223, ZN => n1276);
   U1428 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n274, B1 => 
                           REGISTERS_26_7_port, B2 => n257, ZN => n1275);
   U1429 : AND4_X1 port map( A1 => n1278, A2 => n1277, A3 => n1276, A4 => n1275
                           , ZN => n1290);
   U1430 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n172, B1 => 
                           REGISTERS_7_7_port, B2 => n155_port, ZN => n1282);
   U1431 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n206, B1 => 
                           REGISTERS_3_7_port, B2 => n189, ZN => n1281);
   U1432 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n240, B1 => 
                           REGISTERS_6_7_port, B2 => n223, ZN => n1280);
   U1433 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n274, B1 => 
                           REGISTERS_2_7_port, B2 => n257, ZN => n1279);
   U1434 : NAND4_X1 port map( A1 => n1282, A2 => n1281, A3 => n1280, A4 => 
                           n1279, ZN => n1288);
   U1435 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n172, B1 => 
                           REGISTERS_15_7_port, B2 => n155_port, ZN => n1286);
   U1436 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n206, B1 => 
                           REGISTERS_11_7_port, B2 => n189, ZN => n1285);
   U1437 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n240, B1 => 
                           REGISTERS_14_7_port, B2 => n223, ZN => n1284);
   U1438 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n274, B1 => 
                           REGISTERS_10_7_port, B2 => n257, ZN => n1283);
   U1439 : NAND4_X1 port map( A1 => n1286, A2 => n1285, A3 => n1284, A4 => 
                           n1283, ZN => n1287);
   U1440 : AOI22_X1 port map( A1 => n1288, A2 => n2818, B1 => n1287, B2 => 
                           n2816, ZN => n1289);
   U1441 : OAI221_X1 port map( B1 => n2822, B2 => n1291, C1 => n2820, C2 => 
                           n1290, A => n1289, ZN => N151);
   U1442 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n172, B1 => 
                           REGISTERS_23_8_port, B2 => n155_port, ZN => n1295);
   U1443 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n206, B1 => 
                           REGISTERS_19_8_port, B2 => n189, ZN => n1294);
   U1444 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n240, B1 => 
                           REGISTERS_22_8_port, B2 => n223, ZN => n1293);
   U1445 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n274, B1 => 
                           REGISTERS_18_8_port, B2 => n257, ZN => n1292);
   U1446 : AND4_X1 port map( A1 => n1295, A2 => n1294, A3 => n1293, A4 => n1292
                           , ZN => n2336);
   U1447 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n172, B1 => 
                           REGISTERS_31_8_port, B2 => n155_port, ZN => n1299);
   U1448 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n206, B1 => 
                           REGISTERS_27_8_port, B2 => n189, ZN => n1298);
   U1449 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n240, B1 => 
                           REGISTERS_30_8_port, B2 => n223, ZN => n1297);
   U1450 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n274, B1 => 
                           REGISTERS_26_8_port, B2 => n257, ZN => n1296);
   U1451 : AND4_X1 port map( A1 => n1299, A2 => n1298, A3 => n1297, A4 => n1296
                           , ZN => n2335);
   U1452 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n172, B1 => 
                           REGISTERS_7_8_port, B2 => n155_port, ZN => n2327);
   U1453 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n206, B1 => 
                           REGISTERS_3_8_port, B2 => n189, ZN => n1302);
   U1454 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n240, B1 => 
                           REGISTERS_6_8_port, B2 => n223, ZN => n1301);
   U1455 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n274, B1 => 
                           REGISTERS_2_8_port, B2 => n257, ZN => n1300);
   U1456 : NAND4_X1 port map( A1 => n2327, A2 => n1302, A3 => n1301, A4 => 
                           n1300, ZN => n2333);
   U1457 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n172, B1 => 
                           REGISTERS_15_8_port, B2 => n155_port, ZN => n2331);
   U1458 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n206, B1 => 
                           REGISTERS_11_8_port, B2 => n189, ZN => n2330);
   U1459 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n240, B1 => 
                           REGISTERS_14_8_port, B2 => n223, ZN => n2329);
   U1460 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n274, B1 => 
                           REGISTERS_10_8_port, B2 => n257, ZN => n2328);
   U1461 : NAND4_X1 port map( A1 => n2331, A2 => n2330, A3 => n2329, A4 => 
                           n2328, ZN => n2332);
   U1462 : AOI22_X1 port map( A1 => n2333, A2 => n2818, B1 => n2332, B2 => 
                           n2816, ZN => n2334);
   U1463 : OAI221_X1 port map( B1 => n2822, B2 => n2336, C1 => n2820, C2 => 
                           n2335, A => n2334, ZN => N150);
   U1464 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n173, B1 => 
                           REGISTERS_23_9_port, B2 => n156_port, ZN => n2340);
   U1465 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n207, B1 => 
                           REGISTERS_19_9_port, B2 => n190, ZN => n2339);
   U1466 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n241, B1 => 
                           REGISTERS_22_9_port, B2 => n224, ZN => n2338);
   U1467 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n275, B1 => 
                           REGISTERS_18_9_port, B2 => n258, ZN => n2337);
   U1468 : AND4_X1 port map( A1 => n2340, A2 => n2339, A3 => n2338, A4 => n2337
                           , ZN => n2357);
   U1469 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n173, B1 => 
                           REGISTERS_31_9_port, B2 => n156_port, ZN => n2344);
   U1470 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n207, B1 => 
                           REGISTERS_27_9_port, B2 => n190, ZN => n2343);
   U1471 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n241, B1 => 
                           REGISTERS_30_9_port, B2 => n224, ZN => n2342);
   U1472 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n275, B1 => 
                           REGISTERS_26_9_port, B2 => n258, ZN => n2341);
   U1473 : AND4_X1 port map( A1 => n2344, A2 => n2343, A3 => n2342, A4 => n2341
                           , ZN => n2356);
   U1474 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n173, B1 => 
                           REGISTERS_7_9_port, B2 => n156_port, ZN => n2348);
   U1475 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n207, B1 => 
                           REGISTERS_3_9_port, B2 => n190, ZN => n2347);
   U1476 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n241, B1 => 
                           REGISTERS_6_9_port, B2 => n224, ZN => n2346);
   U1477 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n275, B1 => 
                           REGISTERS_2_9_port, B2 => n258, ZN => n2345);
   U1478 : NAND4_X1 port map( A1 => n2348, A2 => n2347, A3 => n2346, A4 => 
                           n2345, ZN => n2354);
   U1479 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n173, B1 => 
                           REGISTERS_15_9_port, B2 => n156_port, ZN => n2352);
   U1480 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n207, B1 => 
                           REGISTERS_11_9_port, B2 => n190, ZN => n2351);
   U1481 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n241, B1 => 
                           REGISTERS_14_9_port, B2 => n224, ZN => n2350);
   U1482 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n275, B1 => 
                           REGISTERS_10_9_port, B2 => n258, ZN => n2349);
   U1483 : NAND4_X1 port map( A1 => n2352, A2 => n2351, A3 => n2350, A4 => 
                           n2349, ZN => n2353);
   U1484 : AOI22_X1 port map( A1 => n2354, A2 => n2818, B1 => n2353, B2 => 
                           n2816, ZN => n2355);
   U1485 : OAI221_X1 port map( B1 => n2822, B2 => n2357, C1 => n2820, C2 => 
                           n2356, A => n2355, ZN => N149);
   U1486 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n173, B1 => 
                           REGISTERS_23_10_port, B2 => n156_port, ZN => n2361);
   U1487 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n207, B1 => 
                           REGISTERS_19_10_port, B2 => n190, ZN => n2360);
   U1488 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n241, B1 => 
                           REGISTERS_22_10_port, B2 => n224, ZN => n2359);
   U1489 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n275, B1 => 
                           REGISTERS_18_10_port, B2 => n258, ZN => n2358);
   U1490 : AND4_X1 port map( A1 => n2361, A2 => n2360, A3 => n2359, A4 => n2358
                           , ZN => n2378);
   U1491 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n173, B1 => 
                           REGISTERS_31_10_port, B2 => n156_port, ZN => n2365);
   U1492 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n207, B1 => 
                           REGISTERS_27_10_port, B2 => n190, ZN => n2364);
   U1493 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n241, B1 => 
                           REGISTERS_30_10_port, B2 => n224, ZN => n2363);
   U1494 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n275, B1 => 
                           REGISTERS_26_10_port, B2 => n258, ZN => n2362);
   U1495 : AND4_X1 port map( A1 => n2365, A2 => n2364, A3 => n2363, A4 => n2362
                           , ZN => n2377);
   U1496 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n173, B1 => 
                           REGISTERS_7_10_port, B2 => n156_port, ZN => n2369);
   U1497 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n207, B1 => 
                           REGISTERS_3_10_port, B2 => n190, ZN => n2368);
   U1498 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n241, B1 => 
                           REGISTERS_6_10_port, B2 => n224, ZN => n2367);
   U1499 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n275, B1 => 
                           REGISTERS_2_10_port, B2 => n258, ZN => n2366);
   U1500 : NAND4_X1 port map( A1 => n2369, A2 => n2368, A3 => n2367, A4 => 
                           n2366, ZN => n2375);
   U1501 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n173, B1 => 
                           REGISTERS_15_10_port, B2 => n156_port, ZN => n2373);
   U1502 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n207, B1 => 
                           REGISTERS_11_10_port, B2 => n190, ZN => n2372);
   U1503 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n241, B1 => 
                           REGISTERS_14_10_port, B2 => n224, ZN => n2371);
   U1504 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n275, B1 => 
                           REGISTERS_10_10_port, B2 => n258, ZN => n2370);
   U1505 : NAND4_X1 port map( A1 => n2373, A2 => n2372, A3 => n2371, A4 => 
                           n2370, ZN => n2374);
   U1506 : AOI22_X1 port map( A1 => n2375, A2 => n2818, B1 => n2374, B2 => 
                           n2816, ZN => n2376);
   U1507 : OAI221_X1 port map( B1 => n2822, B2 => n2378, C1 => n2820, C2 => 
                           n2377, A => n2376, ZN => N148);
   U1508 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n173, B1 => 
                           REGISTERS_23_11_port, B2 => n156_port, ZN => n2382);
   U1509 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n207, B1 => 
                           REGISTERS_19_11_port, B2 => n190, ZN => n2381);
   U1510 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n241, B1 => 
                           REGISTERS_22_11_port, B2 => n224, ZN => n2380);
   U1511 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n275, B1 => 
                           REGISTERS_18_11_port, B2 => n258, ZN => n2379);
   U1512 : AND4_X1 port map( A1 => n2382, A2 => n2381, A3 => n2380, A4 => n2379
                           , ZN => n2399);
   U1513 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n173, B1 => 
                           REGISTERS_31_11_port, B2 => n156_port, ZN => n2386);
   U1514 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n207, B1 => 
                           REGISTERS_27_11_port, B2 => n190, ZN => n2385);
   U1515 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n241, B1 => 
                           REGISTERS_30_11_port, B2 => n224, ZN => n2384);
   U1516 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n275, B1 => 
                           REGISTERS_26_11_port, B2 => n258, ZN => n2383);
   U1517 : AND4_X1 port map( A1 => n2386, A2 => n2385, A3 => n2384, A4 => n2383
                           , ZN => n2398);
   U1518 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n173, B1 => 
                           REGISTERS_7_11_port, B2 => n156_port, ZN => n2390);
   U1519 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n207, B1 => 
                           REGISTERS_3_11_port, B2 => n190, ZN => n2389);
   U1520 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n241, B1 => 
                           REGISTERS_6_11_port, B2 => n224, ZN => n2388);
   U1521 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n275, B1 => 
                           REGISTERS_2_11_port, B2 => n258, ZN => n2387);
   U1522 : NAND4_X1 port map( A1 => n2390, A2 => n2389, A3 => n2388, A4 => 
                           n2387, ZN => n2396);
   U1523 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n173, B1 => 
                           REGISTERS_15_11_port, B2 => n156_port, ZN => n2394);
   U1524 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n207, B1 => 
                           REGISTERS_11_11_port, B2 => n190, ZN => n2393);
   U1525 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n241, B1 => 
                           REGISTERS_14_11_port, B2 => n224, ZN => n2392);
   U1526 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n275, B1 => 
                           REGISTERS_10_11_port, B2 => n258, ZN => n2391);
   U1527 : NAND4_X1 port map( A1 => n2394, A2 => n2393, A3 => n2392, A4 => 
                           n2391, ZN => n2395);
   U1528 : AOI22_X1 port map( A1 => n2396, A2 => n2818, B1 => n2395, B2 => 
                           n2816, ZN => n2397);
   U1529 : OAI221_X1 port map( B1 => n2822, B2 => n2399, C1 => n2820, C2 => 
                           n2398, A => n2397, ZN => N147);
   U1530 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n174, B1 => 
                           REGISTERS_23_12_port, B2 => n157_port, ZN => n2403);
   U1531 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n208, B1 => 
                           REGISTERS_19_12_port, B2 => n191, ZN => n2402);
   U1532 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n242, B1 => 
                           REGISTERS_22_12_port, B2 => n225, ZN => n2401);
   U1533 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n276, B1 => 
                           REGISTERS_18_12_port, B2 => n259, ZN => n2400);
   U1534 : AND4_X1 port map( A1 => n2403, A2 => n2402, A3 => n2401, A4 => n2400
                           , ZN => n2420);
   U1535 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n174, B1 => 
                           REGISTERS_31_12_port, B2 => n157_port, ZN => n2407);
   U1536 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n208, B1 => 
                           REGISTERS_27_12_port, B2 => n191, ZN => n2406);
   U1537 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n242, B1 => 
                           REGISTERS_30_12_port, B2 => n225, ZN => n2405);
   U1538 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n276, B1 => 
                           REGISTERS_26_12_port, B2 => n259, ZN => n2404);
   U1539 : AND4_X1 port map( A1 => n2407, A2 => n2406, A3 => n2405, A4 => n2404
                           , ZN => n2419);
   U1540 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n174, B1 => 
                           REGISTERS_7_12_port, B2 => n157_port, ZN => n2411);
   U1541 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n208, B1 => 
                           REGISTERS_3_12_port, B2 => n191, ZN => n2410);
   U1542 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n242, B1 => 
                           REGISTERS_6_12_port, B2 => n225, ZN => n2409);
   U1543 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n276, B1 => 
                           REGISTERS_2_12_port, B2 => n259, ZN => n2408);
   U1544 : NAND4_X1 port map( A1 => n2411, A2 => n2410, A3 => n2409, A4 => 
                           n2408, ZN => n2417);
   U1545 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n174, B1 => 
                           REGISTERS_15_12_port, B2 => n157_port, ZN => n2415);
   U1546 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n208, B1 => 
                           REGISTERS_11_12_port, B2 => n191, ZN => n2414);
   U1547 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n242, B1 => 
                           REGISTERS_14_12_port, B2 => n225, ZN => n2413);
   U1548 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n276, B1 => 
                           REGISTERS_10_12_port, B2 => n259, ZN => n2412);
   U1549 : NAND4_X1 port map( A1 => n2415, A2 => n2414, A3 => n2413, A4 => 
                           n2412, ZN => n2416);
   U1550 : AOI22_X1 port map( A1 => n2417, A2 => n2818, B1 => n2416, B2 => 
                           n2816, ZN => n2418);
   U1551 : OAI221_X1 port map( B1 => n2822, B2 => n2420, C1 => n2820, C2 => 
                           n2419, A => n2418, ZN => N146);
   U1552 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n174, B1 => 
                           REGISTERS_23_13_port, B2 => n157_port, ZN => n2424);
   U1553 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n208, B1 => 
                           REGISTERS_19_13_port, B2 => n191, ZN => n2423);
   U1554 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n242, B1 => 
                           REGISTERS_22_13_port, B2 => n225, ZN => n2422);
   U1555 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n276, B1 => 
                           REGISTERS_18_13_port, B2 => n259, ZN => n2421);
   U1556 : AND4_X1 port map( A1 => n2424, A2 => n2423, A3 => n2422, A4 => n2421
                           , ZN => n2441);
   U1557 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n174, B1 => 
                           REGISTERS_31_13_port, B2 => n157_port, ZN => n2428);
   U1558 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n208, B1 => 
                           REGISTERS_27_13_port, B2 => n191, ZN => n2427);
   U1559 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n242, B1 => 
                           REGISTERS_30_13_port, B2 => n225, ZN => n2426);
   U1560 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n276, B1 => 
                           REGISTERS_26_13_port, B2 => n259, ZN => n2425);
   U1561 : AND4_X1 port map( A1 => n2428, A2 => n2427, A3 => n2426, A4 => n2425
                           , ZN => n2440);
   U1562 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n174, B1 => 
                           REGISTERS_7_13_port, B2 => n157_port, ZN => n2432);
   U1563 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n208, B1 => 
                           REGISTERS_3_13_port, B2 => n191, ZN => n2431);
   U1564 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n242, B1 => 
                           REGISTERS_6_13_port, B2 => n225, ZN => n2430);
   U1565 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n276, B1 => 
                           REGISTERS_2_13_port, B2 => n259, ZN => n2429);
   U1566 : NAND4_X1 port map( A1 => n2432, A2 => n2431, A3 => n2430, A4 => 
                           n2429, ZN => n2438);
   U1567 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n174, B1 => 
                           REGISTERS_15_13_port, B2 => n157_port, ZN => n2436);
   U1568 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n208, B1 => 
                           REGISTERS_11_13_port, B2 => n191, ZN => n2435);
   U1569 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n242, B1 => 
                           REGISTERS_14_13_port, B2 => n225, ZN => n2434);
   U1570 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n276, B1 => 
                           REGISTERS_10_13_port, B2 => n259, ZN => n2433);
   U1571 : NAND4_X1 port map( A1 => n2436, A2 => n2435, A3 => n2434, A4 => 
                           n2433, ZN => n2437);
   U1572 : AOI22_X1 port map( A1 => n2438, A2 => n2818, B1 => n2437, B2 => 
                           n2816, ZN => n2439);
   U1573 : OAI221_X1 port map( B1 => n2822, B2 => n2441, C1 => n2820, C2 => 
                           n2440, A => n2439, ZN => N145);
   U1574 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n174, B1 => 
                           REGISTERS_23_14_port, B2 => n157_port, ZN => n2445);
   U1575 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n208, B1 => 
                           REGISTERS_19_14_port, B2 => n191, ZN => n2444);
   U1576 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n242, B1 => 
                           REGISTERS_22_14_port, B2 => n225, ZN => n2443);
   U1577 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n276, B1 => 
                           REGISTERS_18_14_port, B2 => n259, ZN => n2442);
   U1578 : AND4_X1 port map( A1 => n2445, A2 => n2444, A3 => n2443, A4 => n2442
                           , ZN => n2462);
   U1579 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n174, B1 => 
                           REGISTERS_31_14_port, B2 => n157_port, ZN => n2449);
   U1580 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n208, B1 => 
                           REGISTERS_27_14_port, B2 => n191, ZN => n2448);
   U1581 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n242, B1 => 
                           REGISTERS_30_14_port, B2 => n225, ZN => n2447);
   U1582 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n276, B1 => 
                           REGISTERS_26_14_port, B2 => n259, ZN => n2446);
   U1583 : AND4_X1 port map( A1 => n2449, A2 => n2448, A3 => n2447, A4 => n2446
                           , ZN => n2461);
   U1584 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n174, B1 => 
                           REGISTERS_7_14_port, B2 => n157_port, ZN => n2453);
   U1585 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n208, B1 => 
                           REGISTERS_3_14_port, B2 => n191, ZN => n2452);
   U1586 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n242, B1 => 
                           REGISTERS_6_14_port, B2 => n225, ZN => n2451);
   U1587 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n276, B1 => 
                           REGISTERS_2_14_port, B2 => n259, ZN => n2450);
   U1588 : NAND4_X1 port map( A1 => n2453, A2 => n2452, A3 => n2451, A4 => 
                           n2450, ZN => n2459);
   U1589 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n174, B1 => 
                           REGISTERS_15_14_port, B2 => n157_port, ZN => n2457);
   U1590 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n208, B1 => 
                           REGISTERS_11_14_port, B2 => n191, ZN => n2456);
   U1591 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n242, B1 => 
                           REGISTERS_14_14_port, B2 => n225, ZN => n2455);
   U1592 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n276, B1 => 
                           REGISTERS_10_14_port, B2 => n259, ZN => n2454);
   U1593 : NAND4_X1 port map( A1 => n2457, A2 => n2456, A3 => n2455, A4 => 
                           n2454, ZN => n2458);
   U1594 : AOI22_X1 port map( A1 => n2459, A2 => n2818, B1 => n2458, B2 => 
                           n2816, ZN => n2460);
   U1595 : OAI221_X1 port map( B1 => n2822, B2 => n2462, C1 => n2820, C2 => 
                           n2461, A => n2460, ZN => N144);
   U1596 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n175, B1 => 
                           REGISTERS_23_15_port, B2 => n158_port, ZN => n2466);
   U1597 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n209, B1 => 
                           REGISTERS_19_15_port, B2 => n192, ZN => n2465);
   U1598 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n243, B1 => 
                           REGISTERS_22_15_port, B2 => n226, ZN => n2464);
   U1599 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n277, B1 => 
                           REGISTERS_18_15_port, B2 => n260, ZN => n2463);
   U1600 : AND4_X1 port map( A1 => n2466, A2 => n2465, A3 => n2464, A4 => n2463
                           , ZN => n2483);
   U1601 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n175, B1 => 
                           REGISTERS_31_15_port, B2 => n158_port, ZN => n2470);
   U1602 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n209, B1 => 
                           REGISTERS_27_15_port, B2 => n192, ZN => n2469);
   U1603 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n243, B1 => 
                           REGISTERS_30_15_port, B2 => n226, ZN => n2468);
   U1604 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n277, B1 => 
                           REGISTERS_26_15_port, B2 => n260, ZN => n2467);
   U1605 : AND4_X1 port map( A1 => n2470, A2 => n2469, A3 => n2468, A4 => n2467
                           , ZN => n2482);
   U1606 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n175, B1 => 
                           REGISTERS_7_15_port, B2 => n158_port, ZN => n2474);
   U1607 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n209, B1 => 
                           REGISTERS_3_15_port, B2 => n192, ZN => n2473);
   U1608 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n243, B1 => 
                           REGISTERS_6_15_port, B2 => n226, ZN => n2472);
   U1609 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n277, B1 => 
                           REGISTERS_2_15_port, B2 => n260, ZN => n2471);
   U1610 : NAND4_X1 port map( A1 => n2474, A2 => n2473, A3 => n2472, A4 => 
                           n2471, ZN => n2480);
   U1611 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n175, B1 => 
                           REGISTERS_15_15_port, B2 => n158_port, ZN => n2478);
   U1612 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n209, B1 => 
                           REGISTERS_11_15_port, B2 => n192, ZN => n2477);
   U1613 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n243, B1 => 
                           REGISTERS_14_15_port, B2 => n226, ZN => n2476);
   U1614 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n277, B1 => 
                           REGISTERS_10_15_port, B2 => n260, ZN => n2475);
   U1615 : NAND4_X1 port map( A1 => n2478, A2 => n2477, A3 => n2476, A4 => 
                           n2475, ZN => n2479);
   U1616 : AOI22_X1 port map( A1 => n2480, A2 => n2818, B1 => n2479, B2 => 
                           n2816, ZN => n2481);
   U1617 : OAI221_X1 port map( B1 => n2822, B2 => n2483, C1 => n2820, C2 => 
                           n2482, A => n2481, ZN => N143);
   U1618 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n175, B1 => 
                           REGISTERS_23_16_port, B2 => n158_port, ZN => n2487);
   U1619 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n209, B1 => 
                           REGISTERS_19_16_port, B2 => n192, ZN => n2486);
   U1620 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n243, B1 => 
                           REGISTERS_22_16_port, B2 => n226, ZN => n2485);
   U1621 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n277, B1 => 
                           REGISTERS_18_16_port, B2 => n260, ZN => n2484);
   U1622 : AND4_X1 port map( A1 => n2487, A2 => n2486, A3 => n2485, A4 => n2484
                           , ZN => n2504);
   U1623 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n175, B1 => 
                           REGISTERS_31_16_port, B2 => n158_port, ZN => n2491);
   U1624 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n209, B1 => 
                           REGISTERS_27_16_port, B2 => n192, ZN => n2490);
   U1625 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n243, B1 => 
                           REGISTERS_30_16_port, B2 => n226, ZN => n2489);
   U1626 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n277, B1 => 
                           REGISTERS_26_16_port, B2 => n260, ZN => n2488);
   U1627 : AND4_X1 port map( A1 => n2491, A2 => n2490, A3 => n2489, A4 => n2488
                           , ZN => n2503);
   U1628 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n175, B1 => 
                           REGISTERS_7_16_port, B2 => n158_port, ZN => n2495);
   U1629 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n209, B1 => 
                           REGISTERS_3_16_port, B2 => n192, ZN => n2494);
   U1630 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n243, B1 => 
                           REGISTERS_6_16_port, B2 => n226, ZN => n2493);
   U1631 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n277, B1 => 
                           REGISTERS_2_16_port, B2 => n260, ZN => n2492);
   U1632 : NAND4_X1 port map( A1 => n2495, A2 => n2494, A3 => n2493, A4 => 
                           n2492, ZN => n2501);
   U1633 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n175, B1 => 
                           REGISTERS_15_16_port, B2 => n158_port, ZN => n2499);
   U1634 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n209, B1 => 
                           REGISTERS_11_16_port, B2 => n192, ZN => n2498);
   U1635 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n243, B1 => 
                           REGISTERS_14_16_port, B2 => n226, ZN => n2497);
   U1636 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n277, B1 => 
                           REGISTERS_10_16_port, B2 => n260, ZN => n2496);
   U1637 : NAND4_X1 port map( A1 => n2499, A2 => n2498, A3 => n2497, A4 => 
                           n2496, ZN => n2500);
   U1638 : AOI22_X1 port map( A1 => n2501, A2 => n2818, B1 => n2500, B2 => 
                           n2816, ZN => n2502);
   U1639 : OAI221_X1 port map( B1 => n2822, B2 => n2504, C1 => n2820, C2 => 
                           n2503, A => n2502, ZN => N142);
   U1640 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n175, B1 => 
                           REGISTERS_23_17_port, B2 => n158_port, ZN => n2508);
   U1641 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n209, B1 => 
                           REGISTERS_19_17_port, B2 => n192, ZN => n2507);
   U1642 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n243, B1 => 
                           REGISTERS_22_17_port, B2 => n226, ZN => n2506);
   U1643 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n277, B1 => 
                           REGISTERS_18_17_port, B2 => n260, ZN => n2505);
   U1644 : AND4_X1 port map( A1 => n2508, A2 => n2507, A3 => n2506, A4 => n2505
                           , ZN => n2525);
   U1645 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n175, B1 => 
                           REGISTERS_31_17_port, B2 => n158_port, ZN => n2512);
   U1646 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n209, B1 => 
                           REGISTERS_27_17_port, B2 => n192, ZN => n2511);
   U1647 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n243, B1 => 
                           REGISTERS_30_17_port, B2 => n226, ZN => n2510);
   U1648 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n277, B1 => 
                           REGISTERS_26_17_port, B2 => n260, ZN => n2509);
   U1649 : AND4_X1 port map( A1 => n2512, A2 => n2511, A3 => n2510, A4 => n2509
                           , ZN => n2524);
   U1650 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n175, B1 => 
                           REGISTERS_7_17_port, B2 => n158_port, ZN => n2516);
   U1651 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n209, B1 => 
                           REGISTERS_3_17_port, B2 => n192, ZN => n2515);
   U1652 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n243, B1 => 
                           REGISTERS_6_17_port, B2 => n226, ZN => n2514);
   U1653 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n277, B1 => 
                           REGISTERS_2_17_port, B2 => n260, ZN => n2513);
   U1654 : NAND4_X1 port map( A1 => n2516, A2 => n2515, A3 => n2514, A4 => 
                           n2513, ZN => n2522);
   U1655 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n175, B1 => 
                           REGISTERS_15_17_port, B2 => n158_port, ZN => n2520);
   U1656 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n209, B1 => 
                           REGISTERS_11_17_port, B2 => n192, ZN => n2519);
   U1657 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n243, B1 => 
                           REGISTERS_14_17_port, B2 => n226, ZN => n2518);
   U1658 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n277, B1 => 
                           REGISTERS_10_17_port, B2 => n260, ZN => n2517);
   U1659 : NAND4_X1 port map( A1 => n2520, A2 => n2519, A3 => n2518, A4 => 
                           n2517, ZN => n2521);
   U1660 : AOI22_X1 port map( A1 => n2522, A2 => n2818, B1 => n2521, B2 => 
                           n2816, ZN => n2523);
   U1661 : OAI221_X1 port map( B1 => n2822, B2 => n2525, C1 => n2820, C2 => 
                           n2524, A => n2523, ZN => N141);
   U1662 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n176, B1 => 
                           REGISTERS_23_18_port, B2 => n159, ZN => n2529);
   U1663 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n210, B1 => 
                           REGISTERS_19_18_port, B2 => n193, ZN => n2528);
   U1664 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n244, B1 => 
                           REGISTERS_22_18_port, B2 => n227, ZN => n2527);
   U1665 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n278, B1 => 
                           REGISTERS_18_18_port, B2 => n261, ZN => n2526);
   U1666 : AND4_X1 port map( A1 => n2529, A2 => n2528, A3 => n2527, A4 => n2526
                           , ZN => n2546);
   U1667 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n176, B1 => 
                           REGISTERS_31_18_port, B2 => n159, ZN => n2533);
   U1668 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n210, B1 => 
                           REGISTERS_27_18_port, B2 => n193, ZN => n2532);
   U1669 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n244, B1 => 
                           REGISTERS_30_18_port, B2 => n227, ZN => n2531);
   U1670 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n278, B1 => 
                           REGISTERS_26_18_port, B2 => n261, ZN => n2530);
   U1671 : AND4_X1 port map( A1 => n2533, A2 => n2532, A3 => n2531, A4 => n2530
                           , ZN => n2545);
   U1672 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n176, B1 => 
                           REGISTERS_7_18_port, B2 => n159, ZN => n2537);
   U1673 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n210, B1 => 
                           REGISTERS_3_18_port, B2 => n193, ZN => n2536);
   U1674 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n244, B1 => 
                           REGISTERS_6_18_port, B2 => n227, ZN => n2535);
   U1675 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n278, B1 => 
                           REGISTERS_2_18_port, B2 => n261, ZN => n2534);
   U1676 : NAND4_X1 port map( A1 => n2537, A2 => n2536, A3 => n2535, A4 => 
                           n2534, ZN => n2543);
   U1677 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n176, B1 => 
                           REGISTERS_15_18_port, B2 => n159, ZN => n2541);
   U1678 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n210, B1 => 
                           REGISTERS_11_18_port, B2 => n193, ZN => n2540);
   U1679 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n244, B1 => 
                           REGISTERS_14_18_port, B2 => n227, ZN => n2539);
   U1680 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n278, B1 => 
                           REGISTERS_10_18_port, B2 => n261, ZN => n2538);
   U1681 : NAND4_X1 port map( A1 => n2541, A2 => n2540, A3 => n2539, A4 => 
                           n2538, ZN => n2542);
   U1682 : AOI22_X1 port map( A1 => n2543, A2 => n2818, B1 => n2542, B2 => 
                           n2816, ZN => n2544);
   U1683 : OAI221_X1 port map( B1 => n2822, B2 => n2546, C1 => n2820, C2 => 
                           n2545, A => n2544, ZN => N140);
   U1684 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n176, B1 => 
                           REGISTERS_23_19_port, B2 => n159, ZN => n2550);
   U1685 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n210, B1 => 
                           REGISTERS_19_19_port, B2 => n193, ZN => n2549);
   U1686 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n244, B1 => 
                           REGISTERS_22_19_port, B2 => n227, ZN => n2548);
   U1687 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n278, B1 => 
                           REGISTERS_18_19_port, B2 => n261, ZN => n2547);
   U1688 : AND4_X1 port map( A1 => n2550, A2 => n2549, A3 => n2548, A4 => n2547
                           , ZN => n2567);
   U1689 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n176, B1 => 
                           REGISTERS_31_19_port, B2 => n159, ZN => n2554);
   U1690 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n210, B1 => 
                           REGISTERS_27_19_port, B2 => n193, ZN => n2553);
   U1691 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n244, B1 => 
                           REGISTERS_30_19_port, B2 => n227, ZN => n2552);
   U1692 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n278, B1 => 
                           REGISTERS_26_19_port, B2 => n261, ZN => n2551);
   U1693 : AND4_X1 port map( A1 => n2554, A2 => n2553, A3 => n2552, A4 => n2551
                           , ZN => n2566);
   U1694 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n176, B1 => 
                           REGISTERS_7_19_port, B2 => n159, ZN => n2558);
   U1695 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n210, B1 => 
                           REGISTERS_3_19_port, B2 => n193, ZN => n2557);
   U1696 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n244, B1 => 
                           REGISTERS_6_19_port, B2 => n227, ZN => n2556);
   U1697 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n278, B1 => 
                           REGISTERS_2_19_port, B2 => n261, ZN => n2555);
   U1698 : NAND4_X1 port map( A1 => n2558, A2 => n2557, A3 => n2556, A4 => 
                           n2555, ZN => n2564);
   U1699 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n176, B1 => 
                           REGISTERS_15_19_port, B2 => n159, ZN => n2562);
   U1700 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n210, B1 => 
                           REGISTERS_11_19_port, B2 => n193, ZN => n2561);
   U1701 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n244, B1 => 
                           REGISTERS_14_19_port, B2 => n227, ZN => n2560);
   U1702 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n278, B1 => 
                           REGISTERS_10_19_port, B2 => n261, ZN => n2559);
   U1703 : NAND4_X1 port map( A1 => n2562, A2 => n2561, A3 => n2560, A4 => 
                           n2559, ZN => n2563);
   U1704 : AOI22_X1 port map( A1 => n2564, A2 => n2818, B1 => n2563, B2 => 
                           n2816, ZN => n2565);
   U1705 : OAI221_X1 port map( B1 => n2822, B2 => n2567, C1 => n2820, C2 => 
                           n2566, A => n2565, ZN => N139);
   U1706 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n176, B1 => 
                           REGISTERS_23_20_port, B2 => n159, ZN => n2571);
   U1707 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n210, B1 => 
                           REGISTERS_19_20_port, B2 => n193, ZN => n2570);
   U1708 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n244, B1 => 
                           REGISTERS_22_20_port, B2 => n227, ZN => n2569);
   U1709 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n278, B1 => 
                           REGISTERS_18_20_port, B2 => n261, ZN => n2568);
   U1710 : AND4_X1 port map( A1 => n2571, A2 => n2570, A3 => n2569, A4 => n2568
                           , ZN => n2588);
   U1711 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n176, B1 => 
                           REGISTERS_31_20_port, B2 => n159, ZN => n2575);
   U1712 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n210, B1 => 
                           REGISTERS_27_20_port, B2 => n193, ZN => n2574);
   U1713 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n244, B1 => 
                           REGISTERS_30_20_port, B2 => n227, ZN => n2573);
   U1714 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n278, B1 => 
                           REGISTERS_26_20_port, B2 => n261, ZN => n2572);
   U1715 : AND4_X1 port map( A1 => n2575, A2 => n2574, A3 => n2573, A4 => n2572
                           , ZN => n2587);
   U1716 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n176, B1 => 
                           REGISTERS_7_20_port, B2 => n159, ZN => n2579);
   U1717 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n210, B1 => 
                           REGISTERS_3_20_port, B2 => n193, ZN => n2578);
   U1718 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n244, B1 => 
                           REGISTERS_6_20_port, B2 => n227, ZN => n2577);
   U1719 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n278, B1 => 
                           REGISTERS_2_20_port, B2 => n261, ZN => n2576);
   U1720 : NAND4_X1 port map( A1 => n2579, A2 => n2578, A3 => n2577, A4 => 
                           n2576, ZN => n2585);
   U1721 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n176, B1 => 
                           REGISTERS_15_20_port, B2 => n159, ZN => n2583);
   U1722 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n210, B1 => 
                           REGISTERS_11_20_port, B2 => n193, ZN => n2582);
   U1723 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n244, B1 => 
                           REGISTERS_14_20_port, B2 => n227, ZN => n2581);
   U1724 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n278, B1 => 
                           REGISTERS_10_20_port, B2 => n261, ZN => n2580);
   U1725 : NAND4_X1 port map( A1 => n2583, A2 => n2582, A3 => n2581, A4 => 
                           n2580, ZN => n2584);
   U1726 : AOI22_X1 port map( A1 => n2585, A2 => n2818, B1 => n2584, B2 => 
                           n2816, ZN => n2586);
   U1727 : OAI221_X1 port map( B1 => n2822, B2 => n2588, C1 => n2820, C2 => 
                           n2587, A => n2586, ZN => N138);
   U1728 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n177, B1 => 
                           REGISTERS_23_21_port, B2 => n160, ZN => n2592);
   U1729 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n211, B1 => 
                           REGISTERS_19_21_port, B2 => n194, ZN => n2591);
   U1730 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n245, B1 => 
                           REGISTERS_22_21_port, B2 => n228, ZN => n2590);
   U1731 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n279, B1 => 
                           REGISTERS_18_21_port, B2 => n262, ZN => n2589);
   U1732 : AND4_X1 port map( A1 => n2592, A2 => n2591, A3 => n2590, A4 => n2589
                           , ZN => n2609);
   U1733 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n177, B1 => 
                           REGISTERS_31_21_port, B2 => n160, ZN => n2596);
   U1734 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n211, B1 => 
                           REGISTERS_27_21_port, B2 => n194, ZN => n2595);
   U1735 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n245, B1 => 
                           REGISTERS_30_21_port, B2 => n228, ZN => n2594);
   U1736 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n279, B1 => 
                           REGISTERS_26_21_port, B2 => n262, ZN => n2593);
   U1737 : AND4_X1 port map( A1 => n2596, A2 => n2595, A3 => n2594, A4 => n2593
                           , ZN => n2608);
   U1738 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n177, B1 => 
                           REGISTERS_7_21_port, B2 => n160, ZN => n2600);
   U1739 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n211, B1 => 
                           REGISTERS_3_21_port, B2 => n194, ZN => n2599);
   U1740 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n245, B1 => 
                           REGISTERS_6_21_port, B2 => n228, ZN => n2598);
   U1741 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n279, B1 => 
                           REGISTERS_2_21_port, B2 => n262, ZN => n2597);
   U1742 : NAND4_X1 port map( A1 => n2600, A2 => n2599, A3 => n2598, A4 => 
                           n2597, ZN => n2606);
   U1743 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n177, B1 => 
                           REGISTERS_15_21_port, B2 => n160, ZN => n2604);
   U1744 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n211, B1 => 
                           REGISTERS_11_21_port, B2 => n194, ZN => n2603);
   U1745 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n245, B1 => 
                           REGISTERS_14_21_port, B2 => n228, ZN => n2602);
   U1746 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n279, B1 => 
                           REGISTERS_10_21_port, B2 => n262, ZN => n2601);
   U1747 : NAND4_X1 port map( A1 => n2604, A2 => n2603, A3 => n2602, A4 => 
                           n2601, ZN => n2605);
   U1748 : AOI22_X1 port map( A1 => n2606, A2 => n2818, B1 => n2605, B2 => 
                           n2816, ZN => n2607);
   U1749 : OAI221_X1 port map( B1 => n2822, B2 => n2609, C1 => n2820, C2 => 
                           n2608, A => n2607, ZN => N137);
   U1750 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n177, B1 => 
                           REGISTERS_23_22_port, B2 => n160, ZN => n2613);
   U1751 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n211, B1 => 
                           REGISTERS_19_22_port, B2 => n194, ZN => n2612);
   U1752 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n245, B1 => 
                           REGISTERS_22_22_port, B2 => n228, ZN => n2611);
   U1753 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n279, B1 => 
                           REGISTERS_18_22_port, B2 => n262, ZN => n2610);
   U1754 : AND4_X1 port map( A1 => n2613, A2 => n2612, A3 => n2611, A4 => n2610
                           , ZN => n2630);
   U1755 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n177, B1 => 
                           REGISTERS_31_22_port, B2 => n160, ZN => n2617);
   U1756 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n211, B1 => 
                           REGISTERS_27_22_port, B2 => n194, ZN => n2616);
   U1757 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n245, B1 => 
                           REGISTERS_30_22_port, B2 => n228, ZN => n2615);
   U1758 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n279, B1 => 
                           REGISTERS_26_22_port, B2 => n262, ZN => n2614);
   U1759 : AND4_X1 port map( A1 => n2617, A2 => n2616, A3 => n2615, A4 => n2614
                           , ZN => n2629);
   U1760 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n177, B1 => 
                           REGISTERS_7_22_port, B2 => n160, ZN => n2621);
   U1761 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n211, B1 => 
                           REGISTERS_3_22_port, B2 => n194, ZN => n2620);
   U1762 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n245, B1 => 
                           REGISTERS_6_22_port, B2 => n228, ZN => n2619);
   U1763 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n279, B1 => 
                           REGISTERS_2_22_port, B2 => n262, ZN => n2618);
   U1764 : NAND4_X1 port map( A1 => n2621, A2 => n2620, A3 => n2619, A4 => 
                           n2618, ZN => n2627);
   U1765 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n177, B1 => 
                           REGISTERS_15_22_port, B2 => n160, ZN => n2625);
   U1766 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n211, B1 => 
                           REGISTERS_11_22_port, B2 => n194, ZN => n2624);
   U1767 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n245, B1 => 
                           REGISTERS_14_22_port, B2 => n228, ZN => n2623);
   U1768 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n279, B1 => 
                           REGISTERS_10_22_port, B2 => n262, ZN => n2622);
   U1769 : NAND4_X1 port map( A1 => n2625, A2 => n2624, A3 => n2623, A4 => 
                           n2622, ZN => n2626);
   U1770 : AOI22_X1 port map( A1 => n2627, A2 => n2818, B1 => n2626, B2 => 
                           n2816, ZN => n2628);
   U1771 : OAI221_X1 port map( B1 => n2822, B2 => n2630, C1 => n2820, C2 => 
                           n2629, A => n2628, ZN => N136);
   U1772 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n177, B1 => 
                           REGISTERS_23_23_port, B2 => n160, ZN => n2634);
   U1773 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n211, B1 => 
                           REGISTERS_19_23_port, B2 => n194, ZN => n2633);
   U1774 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n245, B1 => 
                           REGISTERS_22_23_port, B2 => n228, ZN => n2632);
   U1775 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n279, B1 => 
                           REGISTERS_18_23_port, B2 => n262, ZN => n2631);
   U1776 : AND4_X1 port map( A1 => n2634, A2 => n2633, A3 => n2632, A4 => n2631
                           , ZN => n2651);
   U1777 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n177, B1 => 
                           REGISTERS_31_23_port, B2 => n160, ZN => n2638);
   U1778 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n211, B1 => 
                           REGISTERS_27_23_port, B2 => n194, ZN => n2637);
   U1779 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n245, B1 => 
                           REGISTERS_30_23_port, B2 => n228, ZN => n2636);
   U1780 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n279, B1 => 
                           REGISTERS_26_23_port, B2 => n262, ZN => n2635);
   U1781 : AND4_X1 port map( A1 => n2638, A2 => n2637, A3 => n2636, A4 => n2635
                           , ZN => n2650);
   U1782 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n177, B1 => 
                           REGISTERS_7_23_port, B2 => n160, ZN => n2642);
   U1783 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n211, B1 => 
                           REGISTERS_3_23_port, B2 => n194, ZN => n2641);
   U1784 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n245, B1 => 
                           REGISTERS_6_23_port, B2 => n228, ZN => n2640);
   U1785 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n279, B1 => 
                           REGISTERS_2_23_port, B2 => n262, ZN => n2639);
   U1786 : NAND4_X1 port map( A1 => n2642, A2 => n2641, A3 => n2640, A4 => 
                           n2639, ZN => n2648);
   U1787 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n177, B1 => 
                           REGISTERS_15_23_port, B2 => n160, ZN => n2646);
   U1788 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n211, B1 => 
                           REGISTERS_11_23_port, B2 => n194, ZN => n2645);
   U1789 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n245, B1 => 
                           REGISTERS_14_23_port, B2 => n228, ZN => n2644);
   U1790 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n279, B1 => 
                           REGISTERS_10_23_port, B2 => n262, ZN => n2643);
   U1791 : NAND4_X1 port map( A1 => n2646, A2 => n2645, A3 => n2644, A4 => 
                           n2643, ZN => n2647);
   U1792 : AOI22_X1 port map( A1 => n2648, A2 => n2818, B1 => n2647, B2 => 
                           n2816, ZN => n2649);
   U1793 : OAI221_X1 port map( B1 => n2822, B2 => n2651, C1 => n2820, C2 => 
                           n2650, A => n2649, ZN => N135);
   U1794 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n178, B1 => 
                           REGISTERS_23_24_port, B2 => n161, ZN => n2655);
   U1795 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n212, B1 => 
                           REGISTERS_19_24_port, B2 => n195, ZN => n2654);
   U1796 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n246, B1 => 
                           REGISTERS_22_24_port, B2 => n229, ZN => n2653);
   U1797 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n280, B1 => 
                           REGISTERS_18_24_port, B2 => n263, ZN => n2652);
   U1798 : AND4_X1 port map( A1 => n2655, A2 => n2654, A3 => n2653, A4 => n2652
                           , ZN => n2672);
   U1799 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n178, B1 => 
                           REGISTERS_31_24_port, B2 => n161, ZN => n2659);
   U1800 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n212, B1 => 
                           REGISTERS_27_24_port, B2 => n195, ZN => n2658);
   U1801 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n246, B1 => 
                           REGISTERS_30_24_port, B2 => n229, ZN => n2657);
   U1802 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n280, B1 => 
                           REGISTERS_26_24_port, B2 => n263, ZN => n2656);
   U1803 : AND4_X1 port map( A1 => n2659, A2 => n2658, A3 => n2657, A4 => n2656
                           , ZN => n2671);
   U1804 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n178, B1 => 
                           REGISTERS_7_24_port, B2 => n161, ZN => n2663);
   U1805 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n212, B1 => 
                           REGISTERS_3_24_port, B2 => n195, ZN => n2662);
   U1806 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n246, B1 => 
                           REGISTERS_6_24_port, B2 => n229, ZN => n2661);
   U1807 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n280, B1 => 
                           REGISTERS_2_24_port, B2 => n263, ZN => n2660);
   U1808 : NAND4_X1 port map( A1 => n2663, A2 => n2662, A3 => n2661, A4 => 
                           n2660, ZN => n2669);
   U1809 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n178, B1 => 
                           REGISTERS_15_24_port, B2 => n161, ZN => n2667);
   U1810 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n212, B1 => 
                           REGISTERS_11_24_port, B2 => n195, ZN => n2666);
   U1811 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n246, B1 => 
                           REGISTERS_14_24_port, B2 => n229, ZN => n2665);
   U1812 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n280, B1 => 
                           REGISTERS_10_24_port, B2 => n263, ZN => n2664);
   U1813 : NAND4_X1 port map( A1 => n2667, A2 => n2666, A3 => n2665, A4 => 
                           n2664, ZN => n2668);
   U1814 : AOI22_X1 port map( A1 => n2669, A2 => n2818, B1 => n2668, B2 => 
                           n2816, ZN => n2670);
   U1815 : OAI221_X1 port map( B1 => n2822, B2 => n2672, C1 => n2820, C2 => 
                           n2671, A => n2670, ZN => N134);
   U1816 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n178, B1 => 
                           REGISTERS_23_25_port, B2 => n161, ZN => n2676);
   U1817 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n212, B1 => 
                           REGISTERS_19_25_port, B2 => n195, ZN => n2675);
   U1818 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n246, B1 => 
                           REGISTERS_22_25_port, B2 => n229, ZN => n2674);
   U1819 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n280, B1 => 
                           REGISTERS_18_25_port, B2 => n263, ZN => n2673);
   U1820 : AND4_X1 port map( A1 => n2676, A2 => n2675, A3 => n2674, A4 => n2673
                           , ZN => n2693);
   U1821 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n178, B1 => 
                           REGISTERS_31_25_port, B2 => n161, ZN => n2680);
   U1822 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n212, B1 => 
                           REGISTERS_27_25_port, B2 => n195, ZN => n2679);
   U1823 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n246, B1 => 
                           REGISTERS_30_25_port, B2 => n229, ZN => n2678);
   U1824 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n280, B1 => 
                           REGISTERS_26_25_port, B2 => n263, ZN => n2677);
   U1825 : AND4_X1 port map( A1 => n2680, A2 => n2679, A3 => n2678, A4 => n2677
                           , ZN => n2692);
   U1826 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n178, B1 => 
                           REGISTERS_7_25_port, B2 => n161, ZN => n2684);
   U1827 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n212, B1 => 
                           REGISTERS_3_25_port, B2 => n195, ZN => n2683);
   U1828 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n246, B1 => 
                           REGISTERS_6_25_port, B2 => n229, ZN => n2682);
   U1829 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n280, B1 => 
                           REGISTERS_2_25_port, B2 => n263, ZN => n2681);
   U1830 : NAND4_X1 port map( A1 => n2684, A2 => n2683, A3 => n2682, A4 => 
                           n2681, ZN => n2690);
   U1831 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n178, B1 => 
                           REGISTERS_15_25_port, B2 => n161, ZN => n2688);
   U1832 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n212, B1 => 
                           REGISTERS_11_25_port, B2 => n195, ZN => n2687);
   U1833 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n246, B1 => 
                           REGISTERS_14_25_port, B2 => n229, ZN => n2686);
   U1834 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n280, B1 => 
                           REGISTERS_10_25_port, B2 => n263, ZN => n2685);
   U1835 : NAND4_X1 port map( A1 => n2688, A2 => n2687, A3 => n2686, A4 => 
                           n2685, ZN => n2689);
   U1836 : AOI22_X1 port map( A1 => n2690, A2 => n2818, B1 => n2689, B2 => 
                           n2816, ZN => n2691);
   U1837 : OAI221_X1 port map( B1 => n2822, B2 => n2693, C1 => n2820, C2 => 
                           n2692, A => n2691, ZN => N133);
   U1838 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n178, B1 => 
                           REGISTERS_23_26_port, B2 => n161, ZN => n2697);
   U1839 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n212, B1 => 
                           REGISTERS_19_26_port, B2 => n195, ZN => n2696);
   U1840 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n246, B1 => 
                           REGISTERS_22_26_port, B2 => n229, ZN => n2695);
   U1841 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n280, B1 => 
                           REGISTERS_18_26_port, B2 => n263, ZN => n2694);
   U1842 : AND4_X1 port map( A1 => n2697, A2 => n2696, A3 => n2695, A4 => n2694
                           , ZN => n2714);
   U1843 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n178, B1 => 
                           REGISTERS_31_26_port, B2 => n161, ZN => n2701);
   U1844 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n212, B1 => 
                           REGISTERS_27_26_port, B2 => n195, ZN => n2700);
   U1845 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n246, B1 => 
                           REGISTERS_30_26_port, B2 => n229, ZN => n2699);
   U1846 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n280, B1 => 
                           REGISTERS_26_26_port, B2 => n263, ZN => n2698);
   U1847 : AND4_X1 port map( A1 => n2701, A2 => n2700, A3 => n2699, A4 => n2698
                           , ZN => n2713);
   U1848 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n178, B1 => 
                           REGISTERS_7_26_port, B2 => n161, ZN => n2705);
   U1849 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n212, B1 => 
                           REGISTERS_3_26_port, B2 => n195, ZN => n2704);
   U1850 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n246, B1 => 
                           REGISTERS_6_26_port, B2 => n229, ZN => n2703);
   U1851 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n280, B1 => 
                           REGISTERS_2_26_port, B2 => n263, ZN => n2702);
   U1852 : NAND4_X1 port map( A1 => n2705, A2 => n2704, A3 => n2703, A4 => 
                           n2702, ZN => n2711);
   U1853 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n178, B1 => 
                           REGISTERS_15_26_port, B2 => n161, ZN => n2709);
   U1854 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n212, B1 => 
                           REGISTERS_11_26_port, B2 => n195, ZN => n2708);
   U1855 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n246, B1 => 
                           REGISTERS_14_26_port, B2 => n229, ZN => n2707);
   U1856 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n280, B1 => 
                           REGISTERS_10_26_port, B2 => n263, ZN => n2706);
   U1857 : NAND4_X1 port map( A1 => n2709, A2 => n2708, A3 => n2707, A4 => 
                           n2706, ZN => n2710);
   U1858 : AOI22_X1 port map( A1 => n2711, A2 => n2818, B1 => n2710, B2 => 
                           n2816, ZN => n2712);
   U1859 : OAI221_X1 port map( B1 => n2822, B2 => n2714, C1 => n2820, C2 => 
                           n2713, A => n2712, ZN => N132);
   U1860 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n179, B1 => 
                           REGISTERS_23_27_port, B2 => n162, ZN => n2718);
   U1861 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n213, B1 => 
                           REGISTERS_19_27_port, B2 => n196, ZN => n2717);
   U1862 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n247, B1 => 
                           REGISTERS_22_27_port, B2 => n230, ZN => n2716);
   U1863 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n281, B1 => 
                           REGISTERS_18_27_port, B2 => n264, ZN => n2715);
   U1864 : AND4_X1 port map( A1 => n2718, A2 => n2717, A3 => n2716, A4 => n2715
                           , ZN => n2735);
   U1865 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n179, B1 => 
                           REGISTERS_31_27_port, B2 => n162, ZN => n2722);
   U1866 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n213, B1 => 
                           REGISTERS_27_27_port, B2 => n196, ZN => n2721);
   U1867 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n247, B1 => 
                           REGISTERS_30_27_port, B2 => n230, ZN => n2720);
   U1868 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n281, B1 => 
                           REGISTERS_26_27_port, B2 => n264, ZN => n2719);
   U1869 : AND4_X1 port map( A1 => n2722, A2 => n2721, A3 => n2720, A4 => n2719
                           , ZN => n2734);
   U1870 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n179, B1 => 
                           REGISTERS_7_27_port, B2 => n162, ZN => n2726);
   U1871 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n213, B1 => 
                           REGISTERS_3_27_port, B2 => n196, ZN => n2725);
   U1872 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n247, B1 => 
                           REGISTERS_6_27_port, B2 => n230, ZN => n2724);
   U1873 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n281, B1 => 
                           REGISTERS_2_27_port, B2 => n264, ZN => n2723);
   U1874 : NAND4_X1 port map( A1 => n2726, A2 => n2725, A3 => n2724, A4 => 
                           n2723, ZN => n2732);
   U1875 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n179, B1 => 
                           REGISTERS_15_27_port, B2 => n162, ZN => n2730);
   U1876 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n213, B1 => 
                           REGISTERS_11_27_port, B2 => n196, ZN => n2729);
   U1877 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n247, B1 => 
                           REGISTERS_14_27_port, B2 => n230, ZN => n2728);
   U1878 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n281, B1 => 
                           REGISTERS_10_27_port, B2 => n264, ZN => n2727);
   U1879 : NAND4_X1 port map( A1 => n2730, A2 => n2729, A3 => n2728, A4 => 
                           n2727, ZN => n2731);
   U1880 : AOI22_X1 port map( A1 => n2732, A2 => n2818, B1 => n2731, B2 => 
                           n2816, ZN => n2733);
   U1881 : OAI221_X1 port map( B1 => n2822, B2 => n2735, C1 => n2820, C2 => 
                           n2734, A => n2733, ZN => N131);
   U1882 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n179, B1 => 
                           REGISTERS_23_28_port, B2 => n162, ZN => n2739);
   U1883 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n213, B1 => 
                           REGISTERS_19_28_port, B2 => n196, ZN => n2738);
   U1884 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n247, B1 => 
                           REGISTERS_22_28_port, B2 => n230, ZN => n2737);
   U1885 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n281, B1 => 
                           REGISTERS_18_28_port, B2 => n264, ZN => n2736);
   U1886 : AND4_X1 port map( A1 => n2739, A2 => n2738, A3 => n2737, A4 => n2736
                           , ZN => n2756);
   U1887 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n179, B1 => 
                           REGISTERS_31_28_port, B2 => n162, ZN => n2743);
   U1888 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n213, B1 => 
                           REGISTERS_27_28_port, B2 => n196, ZN => n2742);
   U1889 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n247, B1 => 
                           REGISTERS_30_28_port, B2 => n230, ZN => n2741);
   U1890 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n281, B1 => 
                           REGISTERS_26_28_port, B2 => n264, ZN => n2740);
   U1891 : AND4_X1 port map( A1 => n2743, A2 => n2742, A3 => n2741, A4 => n2740
                           , ZN => n2755);
   U1892 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n179, B1 => 
                           REGISTERS_7_28_port, B2 => n162, ZN => n2747);
   U1893 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n213, B1 => 
                           REGISTERS_3_28_port, B2 => n196, ZN => n2746);
   U1894 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n247, B1 => 
                           REGISTERS_6_28_port, B2 => n230, ZN => n2745);
   U1895 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n281, B1 => 
                           REGISTERS_2_28_port, B2 => n264, ZN => n2744);
   U1896 : NAND4_X1 port map( A1 => n2747, A2 => n2746, A3 => n2745, A4 => 
                           n2744, ZN => n2753);
   U1897 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n179, B1 => 
                           REGISTERS_15_28_port, B2 => n162, ZN => n2751);
   U1898 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n213, B1 => 
                           REGISTERS_11_28_port, B2 => n196, ZN => n2750);
   U1899 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n247, B1 => 
                           REGISTERS_14_28_port, B2 => n230, ZN => n2749);
   U1900 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n281, B1 => 
                           REGISTERS_10_28_port, B2 => n264, ZN => n2748);
   U1901 : NAND4_X1 port map( A1 => n2751, A2 => n2750, A3 => n2749, A4 => 
                           n2748, ZN => n2752);
   U1902 : AOI22_X1 port map( A1 => n2753, A2 => n2818, B1 => n2752, B2 => 
                           n2816, ZN => n2754);
   U1903 : OAI221_X1 port map( B1 => n2822, B2 => n2756, C1 => n2820, C2 => 
                           n2755, A => n2754, ZN => N130);
   U1904 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n179, B1 => 
                           REGISTERS_23_29_port, B2 => n162, ZN => n2760);
   U1905 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n213, B1 => 
                           REGISTERS_19_29_port, B2 => n196, ZN => n2759);
   U1906 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n247, B1 => 
                           REGISTERS_22_29_port, B2 => n230, ZN => n2758);
   U1907 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n281, B1 => 
                           REGISTERS_18_29_port, B2 => n264, ZN => n2757);
   U1908 : AND4_X1 port map( A1 => n2760, A2 => n2759, A3 => n2758, A4 => n2757
                           , ZN => n2777);
   U1909 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n179, B1 => 
                           REGISTERS_31_29_port, B2 => n162, ZN => n2764);
   U1910 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n213, B1 => 
                           REGISTERS_27_29_port, B2 => n196, ZN => n2763);
   U1911 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n247, B1 => 
                           REGISTERS_30_29_port, B2 => n230, ZN => n2762);
   U1912 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n281, B1 => 
                           REGISTERS_26_29_port, B2 => n264, ZN => n2761);
   U1913 : AND4_X1 port map( A1 => n2764, A2 => n2763, A3 => n2762, A4 => n2761
                           , ZN => n2776);
   U1914 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n179, B1 => 
                           REGISTERS_7_29_port, B2 => n162, ZN => n2768);
   U1915 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n213, B1 => 
                           REGISTERS_3_29_port, B2 => n196, ZN => n2767);
   U1916 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n247, B1 => 
                           REGISTERS_6_29_port, B2 => n230, ZN => n2766);
   U1917 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n281, B1 => 
                           REGISTERS_2_29_port, B2 => n264, ZN => n2765);
   U1918 : NAND4_X1 port map( A1 => n2768, A2 => n2767, A3 => n2766, A4 => 
                           n2765, ZN => n2774);
   U1919 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n179, B1 => 
                           REGISTERS_15_29_port, B2 => n162, ZN => n2772);
   U1920 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n213, B1 => 
                           REGISTERS_11_29_port, B2 => n196, ZN => n2771);
   U1921 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n247, B1 => 
                           REGISTERS_14_29_port, B2 => n230, ZN => n2770);
   U1922 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n281, B1 => 
                           REGISTERS_10_29_port, B2 => n264, ZN => n2769);
   U1923 : NAND4_X1 port map( A1 => n2772, A2 => n2771, A3 => n2770, A4 => 
                           n2769, ZN => n2773);
   U1924 : AOI22_X1 port map( A1 => n2774, A2 => n2818, B1 => n2773, B2 => 
                           n2816, ZN => n2775);
   U1925 : OAI221_X1 port map( B1 => n2822, B2 => n2777, C1 => n2820, C2 => 
                           n2776, A => n2775, ZN => N129);
   U1926 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n180, B1 => 
                           REGISTERS_23_30_port, B2 => n163, ZN => n2781);
   U1927 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n214, B1 => 
                           REGISTERS_19_30_port, B2 => n197, ZN => n2780);
   U1928 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n248, B1 => 
                           REGISTERS_22_30_port, B2 => n231, ZN => n2779);
   U1929 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n282, B1 => 
                           REGISTERS_18_30_port, B2 => n265, ZN => n2778);
   U1930 : AND4_X1 port map( A1 => n2781, A2 => n2780, A3 => n2779, A4 => n2778
                           , ZN => n2798);
   U1931 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n180, B1 => 
                           REGISTERS_31_30_port, B2 => n163, ZN => n2785);
   U1932 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n214, B1 => 
                           REGISTERS_27_30_port, B2 => n197, ZN => n2784);
   U1933 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n248, B1 => 
                           REGISTERS_30_30_port, B2 => n231, ZN => n2783);
   U1934 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n282, B1 => 
                           REGISTERS_26_30_port, B2 => n265, ZN => n2782);
   U1935 : AND4_X1 port map( A1 => n2785, A2 => n2784, A3 => n2783, A4 => n2782
                           , ZN => n2797);
   U1936 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n180, B1 => 
                           REGISTERS_7_30_port, B2 => n163, ZN => n2789);
   U1937 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n214, B1 => 
                           REGISTERS_3_30_port, B2 => n197, ZN => n2788);
   U1938 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n248, B1 => 
                           REGISTERS_6_30_port, B2 => n231, ZN => n2787);
   U1939 : AOI22_X1 port map( A1 => REGISTERS_0_30_port, A2 => n282, B1 => 
                           REGISTERS_2_30_port, B2 => n265, ZN => n2786);
   U1940 : NAND4_X1 port map( A1 => n2789, A2 => n2788, A3 => n2787, A4 => 
                           n2786, ZN => n2795);
   U1941 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n180, B1 => 
                           REGISTERS_15_30_port, B2 => n163, ZN => n2793);
   U1942 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n214, B1 => 
                           REGISTERS_11_30_port, B2 => n197, ZN => n2792);
   U1943 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n248, B1 => 
                           REGISTERS_14_30_port, B2 => n231, ZN => n2791);
   U1944 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n282, B1 => 
                           REGISTERS_10_30_port, B2 => n265, ZN => n2790);
   U1945 : NAND4_X1 port map( A1 => n2793, A2 => n2792, A3 => n2791, A4 => 
                           n2790, ZN => n2794);
   U1946 : AOI22_X1 port map( A1 => n2795, A2 => n2818, B1 => n2794, B2 => 
                           n2816, ZN => n2796);
   U1947 : OAI221_X1 port map( B1 => n2822, B2 => n2798, C1 => n2820, C2 => 
                           n2797, A => n2796, ZN => N128);
   U1948 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n180, B1 => 
                           REGISTERS_23_31_port, B2 => n163, ZN => n2802);
   U1949 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n214, B1 => 
                           REGISTERS_19_31_port, B2 => n197, ZN => n2801);
   U1950 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n248, B1 => 
                           REGISTERS_22_31_port, B2 => n231, ZN => n2800);
   U1951 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n282, B1 => 
                           REGISTERS_18_31_port, B2 => n265, ZN => n2799);
   U1952 : AND4_X1 port map( A1 => n2802, A2 => n2801, A3 => n2800, A4 => n2799
                           , ZN => n2823);
   U1953 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n180, B1 => 
                           REGISTERS_31_31_port, B2 => n163, ZN => n2806);
   U1954 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n214, B1 => 
                           REGISTERS_27_31_port, B2 => n197, ZN => n2805);
   U1955 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n248, B1 => 
                           REGISTERS_30_31_port, B2 => n231, ZN => n2804);
   U1956 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n282, B1 => 
                           REGISTERS_26_31_port, B2 => n265, ZN => n2803);
   U1957 : AND4_X1 port map( A1 => n2806, A2 => n2805, A3 => n2804, A4 => n2803
                           , ZN => n2821);
   U1958 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n180, B1 => 
                           REGISTERS_7_31_port, B2 => n163, ZN => n2810);
   U1959 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n214, B1 => 
                           REGISTERS_3_31_port, B2 => n197, ZN => n2809);
   U1960 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n248, B1 => 
                           REGISTERS_6_31_port, B2 => n231, ZN => n2808);
   U1961 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n282, B1 => 
                           REGISTERS_2_31_port, B2 => n265, ZN => n2807);
   U1962 : NAND4_X1 port map( A1 => n2810, A2 => n2809, A3 => n2808, A4 => 
                           n2807, ZN => n2817);
   U1963 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n180, B1 => 
                           REGISTERS_15_31_port, B2 => n163, ZN => n2814);
   U1964 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n214, B1 => 
                           REGISTERS_11_31_port, B2 => n197, ZN => n2813);
   U1965 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n248, B1 => 
                           REGISTERS_14_31_port, B2 => n231, ZN => n2812);
   U1966 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n282, B1 => 
                           REGISTERS_10_31_port, B2 => n265, ZN => n2811);
   U1967 : NAND4_X1 port map( A1 => n2814, A2 => n2813, A3 => n2812, A4 => 
                           n2811, ZN => n2815);
   U1968 : AOI22_X1 port map( A1 => n2818, A2 => n2817, B1 => n2816, B2 => 
                           n2815, ZN => n2819);
   U1969 : OAI221_X1 port map( B1 => n2823, B2 => n2822, C1 => n2821, C2 => 
                           n2820, A => n2819, ZN => N127);
   U1970 : OAI21_X1 port map( B1 => n3043, B2 => n2828, A => n2829, ZN => n4099
                           );
   U1971 : NAND2_X1 port map( A1 => N158, A2 => n2830, ZN => n2829);
   U1972 : OAI21_X1 port map( B1 => n3044, B2 => n2828, A => n2831, ZN => n4100
                           );
   U1973 : NAND2_X1 port map( A1 => N157, A2 => n2830, ZN => n2831);
   U1974 : OAI21_X1 port map( B1 => n3045, B2 => n2828, A => n2832, ZN => n4101
                           );
   U1975 : NAND2_X1 port map( A1 => N156, A2 => n2830, ZN => n2832);
   U1976 : OAI21_X1 port map( B1 => n3046, B2 => n2828, A => n2833, ZN => n4102
                           );
   U1977 : NAND2_X1 port map( A1 => N155, A2 => n2830, ZN => n2833);
   U1978 : OAI21_X1 port map( B1 => n3047, B2 => n2828, A => n2834, ZN => n4103
                           );
   U1979 : NAND2_X1 port map( A1 => N154, A2 => n2830, ZN => n2834);
   U1980 : OAI21_X1 port map( B1 => n3048, B2 => n2828, A => n2835, ZN => n4104
                           );
   U1981 : NAND2_X1 port map( A1 => N153, A2 => n2830, ZN => n2835);
   U1982 : OAI21_X1 port map( B1 => n3049, B2 => n2828, A => n2836, ZN => n4105
                           );
   U1983 : NAND2_X1 port map( A1 => N152, A2 => n2830, ZN => n2836);
   U1984 : OAI21_X1 port map( B1 => n3050, B2 => n2828, A => n2837, ZN => n4106
                           );
   U1985 : NAND2_X1 port map( A1 => N151, A2 => n2830, ZN => n2837);
   U1986 : OAI21_X1 port map( B1 => n3051, B2 => n2828, A => n2838, ZN => n4107
                           );
   U1987 : NAND2_X1 port map( A1 => N150, A2 => n2830, ZN => n2838);
   U1988 : OAI21_X1 port map( B1 => n3052, B2 => n2828, A => n2839, ZN => n4108
                           );
   U1989 : NAND2_X1 port map( A1 => N149, A2 => n2830, ZN => n2839);
   U1990 : OAI21_X1 port map( B1 => n3053, B2 => n2828, A => n2840, ZN => n4109
                           );
   U1991 : NAND2_X1 port map( A1 => N148, A2 => n2830, ZN => n2840);
   U1992 : OAI21_X1 port map( B1 => n3054, B2 => n2828, A => n2841, ZN => n4110
                           );
   U1993 : NAND2_X1 port map( A1 => N147, A2 => n2830, ZN => n2841);
   U1994 : OAI21_X1 port map( B1 => n3055, B2 => n2828, A => n2842, ZN => n4111
                           );
   U1995 : NAND2_X1 port map( A1 => N146, A2 => n2830, ZN => n2842);
   U1996 : OAI21_X1 port map( B1 => n3056, B2 => n2828, A => n2843, ZN => n4112
                           );
   U1997 : NAND2_X1 port map( A1 => N145, A2 => n2830, ZN => n2843);
   U1998 : OAI21_X1 port map( B1 => n3057, B2 => n2828, A => n2844, ZN => n4113
                           );
   U1999 : NAND2_X1 port map( A1 => N144, A2 => n2830, ZN => n2844);
   U2000 : OAI21_X1 port map( B1 => n3058, B2 => n2828, A => n2845, ZN => n4114
                           );
   U2001 : NAND2_X1 port map( A1 => N143, A2 => n2830, ZN => n2845);
   U2002 : OAI21_X1 port map( B1 => n3059, B2 => n2828, A => n2846, ZN => n4115
                           );
   U2003 : NAND2_X1 port map( A1 => N142, A2 => n2830, ZN => n2846);
   U2004 : OAI21_X1 port map( B1 => n3060, B2 => n2828, A => n2847, ZN => n4116
                           );
   U2005 : NAND2_X1 port map( A1 => N141, A2 => n2830, ZN => n2847);
   U2006 : OAI21_X1 port map( B1 => n3061, B2 => n2828, A => n2848, ZN => n4117
                           );
   U2007 : NAND2_X1 port map( A1 => N140, A2 => n2830, ZN => n2848);
   U2008 : OAI21_X1 port map( B1 => n3062, B2 => n2828, A => n2849, ZN => n4118
                           );
   U2009 : NAND2_X1 port map( A1 => N139, A2 => n2830, ZN => n2849);
   U2010 : OAI21_X1 port map( B1 => n3063, B2 => n2828, A => n2850, ZN => n4119
                           );
   U2011 : NAND2_X1 port map( A1 => N138, A2 => n2830, ZN => n2850);
   U2012 : OAI21_X1 port map( B1 => n3064, B2 => n2828, A => n2851, ZN => n4120
                           );
   U2013 : NAND2_X1 port map( A1 => N137, A2 => n2830, ZN => n2851);
   U2014 : OAI21_X1 port map( B1 => n3065, B2 => n2828, A => n2852, ZN => n4121
                           );
   U2015 : NAND2_X1 port map( A1 => N136, A2 => n2830, ZN => n2852);
   U2016 : OAI21_X1 port map( B1 => n3066, B2 => n2828, A => n2853, ZN => n4122
                           );
   U2017 : NAND2_X1 port map( A1 => N135, A2 => n2830, ZN => n2853);
   U2018 : OAI21_X1 port map( B1 => n3067, B2 => n2828, A => n2854, ZN => n4123
                           );
   U2019 : NAND2_X1 port map( A1 => N134, A2 => n2830, ZN => n2854);
   U2020 : OAI21_X1 port map( B1 => n3068, B2 => n2828, A => n2855, ZN => n4124
                           );
   U2021 : NAND2_X1 port map( A1 => N133, A2 => n2830, ZN => n2855);
   U2022 : OAI21_X1 port map( B1 => n3069, B2 => n2828, A => n2856, ZN => n4125
                           );
   U2023 : NAND2_X1 port map( A1 => N132, A2 => n2830, ZN => n2856);
   U2024 : OAI21_X1 port map( B1 => n3070, B2 => n2828, A => n2857, ZN => n4126
                           );
   U2025 : NAND2_X1 port map( A1 => N131, A2 => n2830, ZN => n2857);
   U2026 : OAI21_X1 port map( B1 => n3071, B2 => n2828, A => n2858, ZN => n4127
                           );
   U2027 : NAND2_X1 port map( A1 => N130, A2 => n2830, ZN => n2858);
   U2028 : OAI21_X1 port map( B1 => n3072, B2 => n2828, A => n2859, ZN => n4128
                           );
   U2029 : NAND2_X1 port map( A1 => N129, A2 => n2830, ZN => n2859);
   U2030 : OAI21_X1 port map( B1 => n3073, B2 => n2828, A => n2860, ZN => n4129
                           );
   U2031 : NAND2_X1 port map( A1 => N128, A2 => n2830, ZN => n2860);
   U2032 : OAI21_X1 port map( B1 => n3074, B2 => n2828, A => n2861, ZN => n4130
                           );
   U2033 : NAND2_X1 port map( A1 => N127, A2 => n2830, ZN => n2861);
   U2034 : NAND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => n2862);
   U2035 : OAI21_X1 port map( B1 => n3011, B2 => n2863, A => n2864, ZN => n4131
                           );
   U2036 : NAND2_X1 port map( A1 => N91, A2 => n2865, ZN => n2864);
   U2037 : OAI21_X1 port map( B1 => n3012, B2 => n2863, A => n2866, ZN => n4132
                           );
   U2038 : NAND2_X1 port map( A1 => N90, A2 => n2865, ZN => n2866);
   U2039 : OAI21_X1 port map( B1 => n3013, B2 => n2863, A => n2867, ZN => n4133
                           );
   U2040 : NAND2_X1 port map( A1 => N89, A2 => n2865, ZN => n2867);
   U2041 : OAI21_X1 port map( B1 => n3014, B2 => n2863, A => n2868, ZN => n4134
                           );
   U2042 : NAND2_X1 port map( A1 => N88, A2 => n2865, ZN => n2868);
   U2043 : OAI21_X1 port map( B1 => n3015, B2 => n2863, A => n2869, ZN => n4135
                           );
   U2044 : NAND2_X1 port map( A1 => N87, A2 => n2865, ZN => n2869);
   U2045 : OAI21_X1 port map( B1 => n3016, B2 => n2863, A => n2870, ZN => n4136
                           );
   U2046 : NAND2_X1 port map( A1 => N86, A2 => n2865, ZN => n2870);
   U2047 : OAI21_X1 port map( B1 => n3017, B2 => n2863, A => n2871, ZN => n4137
                           );
   U2048 : NAND2_X1 port map( A1 => N85, A2 => n2865, ZN => n2871);
   U2049 : OAI21_X1 port map( B1 => n3018, B2 => n2863, A => n2872, ZN => n4138
                           );
   U2050 : NAND2_X1 port map( A1 => N84, A2 => n2865, ZN => n2872);
   U2051 : OAI21_X1 port map( B1 => n3019, B2 => n2863, A => n2873, ZN => n4139
                           );
   U2052 : NAND2_X1 port map( A1 => N83, A2 => n2865, ZN => n2873);
   U2053 : OAI21_X1 port map( B1 => n3020, B2 => n2863, A => n2874, ZN => n4140
                           );
   U2054 : NAND2_X1 port map( A1 => N82, A2 => n2865, ZN => n2874);
   U2055 : OAI21_X1 port map( B1 => n3021, B2 => n2863, A => n2875, ZN => n4141
                           );
   U2056 : NAND2_X1 port map( A1 => N81, A2 => n2865, ZN => n2875);
   U2057 : OAI21_X1 port map( B1 => n3022, B2 => n2863, A => n2876, ZN => n4142
                           );
   U2058 : NAND2_X1 port map( A1 => N80, A2 => n2865, ZN => n2876);
   U2059 : OAI21_X1 port map( B1 => n3023, B2 => n2863, A => n2877, ZN => n4143
                           );
   U2060 : NAND2_X1 port map( A1 => N79, A2 => n2865, ZN => n2877);
   U2061 : OAI21_X1 port map( B1 => n3024, B2 => n2863, A => n2878, ZN => n4144
                           );
   U2062 : NAND2_X1 port map( A1 => N78, A2 => n2865, ZN => n2878);
   U2063 : OAI21_X1 port map( B1 => n3025, B2 => n2863, A => n2879, ZN => n4145
                           );
   U2064 : NAND2_X1 port map( A1 => N77, A2 => n2865, ZN => n2879);
   U2065 : OAI21_X1 port map( B1 => n3026, B2 => n2863, A => n2880, ZN => n4146
                           );
   U2066 : NAND2_X1 port map( A1 => N76, A2 => n2865, ZN => n2880);
   U2067 : OAI21_X1 port map( B1 => n3027, B2 => n2863, A => n2881, ZN => n4147
                           );
   U2068 : NAND2_X1 port map( A1 => N75, A2 => n2865, ZN => n2881);
   U2069 : OAI21_X1 port map( B1 => n3028, B2 => n2863, A => n2882, ZN => n4148
                           );
   U2070 : NAND2_X1 port map( A1 => N74, A2 => n2865, ZN => n2882);
   U2071 : OAI21_X1 port map( B1 => n3029, B2 => n2863, A => n2883, ZN => n4149
                           );
   U2072 : NAND2_X1 port map( A1 => N73, A2 => n2865, ZN => n2883);
   U2073 : OAI21_X1 port map( B1 => n3030, B2 => n2863, A => n2884, ZN => n4150
                           );
   U2074 : NAND2_X1 port map( A1 => N72, A2 => n2865, ZN => n2884);
   U2075 : OAI21_X1 port map( B1 => n3031, B2 => n2863, A => n2885, ZN => n4151
                           );
   U2076 : NAND2_X1 port map( A1 => N71, A2 => n2865, ZN => n2885);
   U2077 : OAI21_X1 port map( B1 => n3032, B2 => n2863, A => n2886, ZN => n4152
                           );
   U2078 : NAND2_X1 port map( A1 => N70, A2 => n2865, ZN => n2886);
   U2079 : OAI21_X1 port map( B1 => n3033, B2 => n2863, A => n2887, ZN => n4153
                           );
   U2080 : NAND2_X1 port map( A1 => N69, A2 => n2865, ZN => n2887);
   U2081 : OAI21_X1 port map( B1 => n3034, B2 => n2863, A => n2888, ZN => n4154
                           );
   U2082 : NAND2_X1 port map( A1 => N68, A2 => n2865, ZN => n2888);
   U2083 : OAI21_X1 port map( B1 => n3035, B2 => n2863, A => n2889, ZN => n4155
                           );
   U2084 : NAND2_X1 port map( A1 => N67, A2 => n2865, ZN => n2889);
   U2085 : OAI21_X1 port map( B1 => n3036, B2 => n2863, A => n2890, ZN => n4156
                           );
   U2086 : NAND2_X1 port map( A1 => N66, A2 => n2865, ZN => n2890);
   U2087 : OAI21_X1 port map( B1 => n3037, B2 => n2863, A => n2891, ZN => n4157
                           );
   U2088 : NAND2_X1 port map( A1 => N65, A2 => n2865, ZN => n2891);
   U2089 : OAI21_X1 port map( B1 => n3038, B2 => n2863, A => n2892, ZN => n4158
                           );
   U2090 : NAND2_X1 port map( A1 => N64, A2 => n2865, ZN => n2892);
   U2091 : OAI21_X1 port map( B1 => n3039, B2 => n2863, A => n2893, ZN => n4159
                           );
   U2092 : NAND2_X1 port map( A1 => N63, A2 => n2865, ZN => n2893);
   U2093 : OAI21_X1 port map( B1 => n3040, B2 => n2863, A => n2894, ZN => n4160
                           );
   U2094 : NAND2_X1 port map( A1 => N62, A2 => n2865, ZN => n2894);
   U2095 : OAI21_X1 port map( B1 => n3041, B2 => n2863, A => n2895, ZN => n4161
                           );
   U2096 : NAND2_X1 port map( A1 => N61, A2 => n2865, ZN => n2895);
   U2097 : OAI21_X1 port map( B1 => n3042, B2 => n2863, A => n2896, ZN => n4162
                           );
   U2098 : NAND2_X1 port map( A1 => N60, A2 => n2865, ZN => n2896);
   U2099 : NAND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => n2897);
   U2100 : OAI22_X1 port map( A1 => n2898, A2 => n2899, B1 => n4098, B2 => 
                           n2900, ZN => n2326);
   U2101 : OAI22_X1 port map( A1 => n2898, A2 => n2901, B1 => n4097, B2 => 
                           n2900, ZN => n2325);
   U2102 : OAI22_X1 port map( A1 => n2898, A2 => n2902, B1 => n4096, B2 => 
                           n2900, ZN => n2324);
   U2103 : OAI22_X1 port map( A1 => n2898, A2 => n2903, B1 => n4095, B2 => 
                           n2900, ZN => n2323);
   U2104 : OAI22_X1 port map( A1 => n2898, A2 => n2904, B1 => n4094, B2 => 
                           n2900, ZN => n2322);
   U2105 : OAI22_X1 port map( A1 => n2898, A2 => n2905, B1 => n4093, B2 => 
                           n2900, ZN => n2321);
   U2106 : OAI22_X1 port map( A1 => n2898, A2 => n2906, B1 => n4092, B2 => 
                           n2900, ZN => n2320);
   U2107 : OAI22_X1 port map( A1 => n2898, A2 => n2907, B1 => n4091, B2 => 
                           n2900, ZN => n2319);
   U2108 : OAI22_X1 port map( A1 => n2898, A2 => n2908, B1 => n4090, B2 => 
                           n2900, ZN => n2318);
   U2109 : OAI22_X1 port map( A1 => n2898, A2 => n2909, B1 => n4089, B2 => 
                           n2900, ZN => n2317);
   U2110 : OAI22_X1 port map( A1 => n2898, A2 => n2910, B1 => n4088, B2 => 
                           n2900, ZN => n2316);
   U2111 : OAI22_X1 port map( A1 => n2898, A2 => n2911, B1 => n4087, B2 => 
                           n2900, ZN => n2315);
   U2112 : OAI22_X1 port map( A1 => n2898, A2 => n2912, B1 => n4086, B2 => 
                           n2900, ZN => n2314);
   U2113 : OAI22_X1 port map( A1 => n2898, A2 => n2913, B1 => n4085, B2 => 
                           n2900, ZN => n2313);
   U2114 : OAI22_X1 port map( A1 => n2898, A2 => n2914, B1 => n4084, B2 => 
                           n2900, ZN => n2312);
   U2115 : OAI22_X1 port map( A1 => n2898, A2 => n2915, B1 => n4083, B2 => 
                           n2900, ZN => n2311);
   U2116 : OAI22_X1 port map( A1 => n2898, A2 => n2916, B1 => n4082, B2 => 
                           n2900, ZN => n2310);
   U2117 : OAI22_X1 port map( A1 => n2898, A2 => n2917, B1 => n4081, B2 => 
                           n2900, ZN => n2309);
   U2118 : OAI22_X1 port map( A1 => n2898, A2 => n2918, B1 => n4080, B2 => 
                           n2900, ZN => n2308);
   U2119 : OAI22_X1 port map( A1 => n2898, A2 => n2919, B1 => n4079, B2 => 
                           n2900, ZN => n2307);
   U2120 : OAI22_X1 port map( A1 => n2898, A2 => n2920, B1 => n4078, B2 => 
                           n2900, ZN => n2306);
   U2121 : OAI22_X1 port map( A1 => n2898, A2 => n2921, B1 => n4077, B2 => 
                           n2900, ZN => n2305);
   U2122 : OAI22_X1 port map( A1 => n2898, A2 => n2922, B1 => n4076, B2 => 
                           n2900, ZN => n2304);
   U2123 : OAI22_X1 port map( A1 => n2898, A2 => n2923, B1 => n4075, B2 => 
                           n2900, ZN => n2303);
   U2124 : OAI22_X1 port map( A1 => n2898, A2 => n2924, B1 => n4074, B2 => 
                           n2900, ZN => n2302);
   U2125 : OAI22_X1 port map( A1 => n2898, A2 => n2925, B1 => n4073, B2 => 
                           n2900, ZN => n2301);
   U2126 : OAI22_X1 port map( A1 => n2898, A2 => n2926, B1 => n4072, B2 => 
                           n2900, ZN => n2300);
   U2127 : OAI22_X1 port map( A1 => n2898, A2 => n2927, B1 => n4071, B2 => 
                           n2900, ZN => n2299);
   U2128 : OAI22_X1 port map( A1 => n2898, A2 => n2928, B1 => n4070, B2 => 
                           n2900, ZN => n2298);
   U2129 : OAI22_X1 port map( A1 => n2898, A2 => n2929, B1 => n4069, B2 => 
                           n2900, ZN => n2297);
   U2130 : OAI22_X1 port map( A1 => n2898, A2 => n2930, B1 => n4068, B2 => 
                           n2900, ZN => n2296);
   U2131 : OAI22_X1 port map( A1 => n2898, A2 => n2931, B1 => n4067, B2 => 
                           n2900, ZN => n2295);
   U2132 : OAI22_X1 port map( A1 => n2899, A2 => n2934, B1 => n4066, B2 => 
                           n2935, ZN => n2294);
   U2133 : OAI22_X1 port map( A1 => n2901, A2 => n2934, B1 => n4065, B2 => 
                           n2935, ZN => n2293);
   U2134 : OAI22_X1 port map( A1 => n2902, A2 => n2934, B1 => n4064, B2 => 
                           n2935, ZN => n2292);
   U2135 : OAI22_X1 port map( A1 => n2903, A2 => n2934, B1 => n4063, B2 => 
                           n2935, ZN => n2291);
   U2136 : OAI22_X1 port map( A1 => n2904, A2 => n2934, B1 => n4062, B2 => 
                           n2935, ZN => n2290);
   U2137 : OAI22_X1 port map( A1 => n2905, A2 => n2934, B1 => n4061, B2 => 
                           n2935, ZN => n2289);
   U2138 : OAI22_X1 port map( A1 => n2906, A2 => n2934, B1 => n4060, B2 => 
                           n2935, ZN => n2288);
   U2139 : OAI22_X1 port map( A1 => n2907, A2 => n2934, B1 => n4059, B2 => 
                           n2935, ZN => n2287);
   U2140 : OAI22_X1 port map( A1 => n2908, A2 => n2934, B1 => n4058, B2 => 
                           n2935, ZN => n2286);
   U2141 : OAI22_X1 port map( A1 => n2909, A2 => n2934, B1 => n4057, B2 => 
                           n2935, ZN => n2285);
   U2142 : OAI22_X1 port map( A1 => n2910, A2 => n2934, B1 => n4056, B2 => 
                           n2935, ZN => n2284);
   U2143 : OAI22_X1 port map( A1 => n2911, A2 => n2934, B1 => n4055, B2 => 
                           n2935, ZN => n2283);
   U2144 : OAI22_X1 port map( A1 => n2912, A2 => n2934, B1 => n4054, B2 => 
                           n2935, ZN => n2282);
   U2145 : OAI22_X1 port map( A1 => n2913, A2 => n2934, B1 => n4053, B2 => 
                           n2935, ZN => n2281);
   U2146 : OAI22_X1 port map( A1 => n2914, A2 => n2934, B1 => n4052, B2 => 
                           n2935, ZN => n2280);
   U2147 : OAI22_X1 port map( A1 => n2915, A2 => n2934, B1 => n4051, B2 => 
                           n2935, ZN => n2279);
   U2148 : OAI22_X1 port map( A1 => n2916, A2 => n2934, B1 => n4050, B2 => 
                           n2935, ZN => n2278);
   U2149 : OAI22_X1 port map( A1 => n2917, A2 => n2934, B1 => n4049, B2 => 
                           n2935, ZN => n2277);
   U2150 : OAI22_X1 port map( A1 => n2918, A2 => n2934, B1 => n4048, B2 => 
                           n2935, ZN => n2276);
   U2151 : OAI22_X1 port map( A1 => n2919, A2 => n2934, B1 => n4047, B2 => 
                           n2935, ZN => n2275);
   U2152 : OAI22_X1 port map( A1 => n2920, A2 => n2934, B1 => n4046, B2 => 
                           n2935, ZN => n2274);
   U2153 : OAI22_X1 port map( A1 => n2921, A2 => n2934, B1 => n4045, B2 => 
                           n2935, ZN => n2273);
   U2154 : OAI22_X1 port map( A1 => n2922, A2 => n2934, B1 => n4044, B2 => 
                           n2935, ZN => n2272);
   U2155 : OAI22_X1 port map( A1 => n2923, A2 => n2934, B1 => n4043, B2 => 
                           n2935, ZN => n2271);
   U2156 : OAI22_X1 port map( A1 => n2924, A2 => n2934, B1 => n4042, B2 => 
                           n2935, ZN => n2270);
   U2157 : OAI22_X1 port map( A1 => n2925, A2 => n2934, B1 => n4041, B2 => 
                           n2935, ZN => n2269);
   U2158 : OAI22_X1 port map( A1 => n2926, A2 => n2934, B1 => n4040, B2 => 
                           n2935, ZN => n2268);
   U2159 : OAI22_X1 port map( A1 => n2927, A2 => n2934, B1 => n4039, B2 => 
                           n2935, ZN => n2267);
   U2160 : OAI22_X1 port map( A1 => n2928, A2 => n2934, B1 => n4038, B2 => 
                           n2935, ZN => n2266);
   U2161 : OAI22_X1 port map( A1 => n2929, A2 => n2934, B1 => n4037, B2 => 
                           n2935, ZN => n2265);
   U2162 : OAI22_X1 port map( A1 => n2930, A2 => n2934, B1 => n4036, B2 => 
                           n2935, ZN => n2264);
   U2163 : OAI22_X1 port map( A1 => n2931, A2 => n2934, B1 => n4035, B2 => 
                           n2935, ZN => n2263);
   U2164 : OAI22_X1 port map( A1 => n2899, A2 => n2937, B1 => n4034, B2 => 
                           n2938, ZN => n2262);
   U2165 : OAI22_X1 port map( A1 => n2901, A2 => n2937, B1 => n4033, B2 => 
                           n2938, ZN => n2261);
   U2166 : OAI22_X1 port map( A1 => n2902, A2 => n2937, B1 => n4032, B2 => 
                           n2938, ZN => n2260);
   U2167 : OAI22_X1 port map( A1 => n2903, A2 => n2937, B1 => n4031, B2 => 
                           n2938, ZN => n2259);
   U2168 : OAI22_X1 port map( A1 => n2904, A2 => n2937, B1 => n4030, B2 => 
                           n2938, ZN => n2258);
   U2169 : OAI22_X1 port map( A1 => n2905, A2 => n2937, B1 => n4029, B2 => 
                           n2938, ZN => n2257);
   U2170 : OAI22_X1 port map( A1 => n2906, A2 => n2937, B1 => n4028, B2 => 
                           n2938, ZN => n2256);
   U2171 : OAI22_X1 port map( A1 => n2907, A2 => n2937, B1 => n4027, B2 => 
                           n2938, ZN => n2255);
   U2172 : OAI22_X1 port map( A1 => n2908, A2 => n2937, B1 => n4026, B2 => 
                           n2938, ZN => n2254);
   U2173 : OAI22_X1 port map( A1 => n2909, A2 => n2937, B1 => n4025, B2 => 
                           n2938, ZN => n2253);
   U2174 : OAI22_X1 port map( A1 => n2910, A2 => n2937, B1 => n4024, B2 => 
                           n2938, ZN => n2252);
   U2175 : OAI22_X1 port map( A1 => n2911, A2 => n2937, B1 => n4023, B2 => 
                           n2938, ZN => n2251);
   U2176 : OAI22_X1 port map( A1 => n2912, A2 => n2937, B1 => n4022, B2 => 
                           n2938, ZN => n2250);
   U2177 : OAI22_X1 port map( A1 => n2913, A2 => n2937, B1 => n4021, B2 => 
                           n2938, ZN => n2249);
   U2178 : OAI22_X1 port map( A1 => n2914, A2 => n2937, B1 => n4020, B2 => 
                           n2938, ZN => n2248);
   U2179 : OAI22_X1 port map( A1 => n2915, A2 => n2937, B1 => n4019, B2 => 
                           n2938, ZN => n2247);
   U2180 : OAI22_X1 port map( A1 => n2916, A2 => n2937, B1 => n4018, B2 => 
                           n2938, ZN => n2246);
   U2181 : OAI22_X1 port map( A1 => n2917, A2 => n2937, B1 => n4017, B2 => 
                           n2938, ZN => n2245);
   U2182 : OAI22_X1 port map( A1 => n2918, A2 => n2937, B1 => n4016, B2 => 
                           n2938, ZN => n2244);
   U2183 : OAI22_X1 port map( A1 => n2919, A2 => n2937, B1 => n4015, B2 => 
                           n2938, ZN => n2243);
   U2184 : OAI22_X1 port map( A1 => n2920, A2 => n2937, B1 => n4014, B2 => 
                           n2938, ZN => n2242);
   U2185 : OAI22_X1 port map( A1 => n2921, A2 => n2937, B1 => n4013, B2 => 
                           n2938, ZN => n2241);
   U2186 : OAI22_X1 port map( A1 => n2922, A2 => n2937, B1 => n4012, B2 => 
                           n2938, ZN => n2240);
   U2187 : OAI22_X1 port map( A1 => n2923, A2 => n2937, B1 => n4011, B2 => 
                           n2938, ZN => n2239);
   U2188 : OAI22_X1 port map( A1 => n2924, A2 => n2937, B1 => n4010, B2 => 
                           n2938, ZN => n2238);
   U2189 : OAI22_X1 port map( A1 => n2925, A2 => n2937, B1 => n4009, B2 => 
                           n2938, ZN => n2237);
   U2190 : OAI22_X1 port map( A1 => n2926, A2 => n2937, B1 => n4008, B2 => 
                           n2938, ZN => n2236);
   U2191 : OAI22_X1 port map( A1 => n2927, A2 => n2937, B1 => n4007, B2 => 
                           n2938, ZN => n2235);
   U2192 : OAI22_X1 port map( A1 => n2928, A2 => n2937, B1 => n4006, B2 => 
                           n2938, ZN => n2234);
   U2193 : OAI22_X1 port map( A1 => n2929, A2 => n2937, B1 => n4005, B2 => 
                           n2938, ZN => n2233);
   U2194 : OAI22_X1 port map( A1 => n2930, A2 => n2937, B1 => n4004, B2 => 
                           n2938, ZN => n2232);
   U2195 : OAI22_X1 port map( A1 => n2931, A2 => n2937, B1 => n4003, B2 => 
                           n2938, ZN => n2231);
   U2196 : OAI22_X1 port map( A1 => n2899, A2 => n2940, B1 => n4002, B2 => 
                           n2941, ZN => n2230);
   U2197 : OAI22_X1 port map( A1 => n2901, A2 => n2940, B1 => n4001, B2 => 
                           n2941, ZN => n2229);
   U2198 : OAI22_X1 port map( A1 => n2902, A2 => n2940, B1 => n4000, B2 => 
                           n2941, ZN => n2228);
   U2199 : OAI22_X1 port map( A1 => n2903, A2 => n2940, B1 => n3999, B2 => 
                           n2941, ZN => n2227);
   U2200 : OAI22_X1 port map( A1 => n2904, A2 => n2940, B1 => n3998, B2 => 
                           n2941, ZN => n2226);
   U2201 : OAI22_X1 port map( A1 => n2905, A2 => n2940, B1 => n3997, B2 => 
                           n2941, ZN => n2225);
   U2202 : OAI22_X1 port map( A1 => n2906, A2 => n2940, B1 => n3996, B2 => 
                           n2941, ZN => n2224);
   U2203 : OAI22_X1 port map( A1 => n2907, A2 => n2940, B1 => n3995, B2 => 
                           n2941, ZN => n2223);
   U2204 : OAI22_X1 port map( A1 => n2908, A2 => n2940, B1 => n3994, B2 => 
                           n2941, ZN => n2222);
   U2205 : OAI22_X1 port map( A1 => n2909, A2 => n2940, B1 => n3993, B2 => 
                           n2941, ZN => n2221);
   U2206 : OAI22_X1 port map( A1 => n2910, A2 => n2940, B1 => n3992, B2 => 
                           n2941, ZN => n2220);
   U2207 : OAI22_X1 port map( A1 => n2911, A2 => n2940, B1 => n3991, B2 => 
                           n2941, ZN => n2219);
   U2208 : OAI22_X1 port map( A1 => n2912, A2 => n2940, B1 => n3990, B2 => 
                           n2941, ZN => n2218);
   U2209 : OAI22_X1 port map( A1 => n2913, A2 => n2940, B1 => n3989, B2 => 
                           n2941, ZN => n2217);
   U2210 : OAI22_X1 port map( A1 => n2914, A2 => n2940, B1 => n3988, B2 => 
                           n2941, ZN => n2216);
   U2211 : OAI22_X1 port map( A1 => n2915, A2 => n2940, B1 => n3987, B2 => 
                           n2941, ZN => n2215);
   U2212 : OAI22_X1 port map( A1 => n2916, A2 => n2940, B1 => n3986, B2 => 
                           n2941, ZN => n2214);
   U2213 : OAI22_X1 port map( A1 => n2917, A2 => n2940, B1 => n3985, B2 => 
                           n2941, ZN => n2213);
   U2214 : OAI22_X1 port map( A1 => n2918, A2 => n2940, B1 => n3984, B2 => 
                           n2941, ZN => n2212);
   U2215 : OAI22_X1 port map( A1 => n2919, A2 => n2940, B1 => n3983, B2 => 
                           n2941, ZN => n2211);
   U2216 : OAI22_X1 port map( A1 => n2920, A2 => n2940, B1 => n3982, B2 => 
                           n2941, ZN => n2210);
   U2217 : OAI22_X1 port map( A1 => n2921, A2 => n2940, B1 => n3981, B2 => 
                           n2941, ZN => n2209);
   U2218 : OAI22_X1 port map( A1 => n2922, A2 => n2940, B1 => n3980, B2 => 
                           n2941, ZN => n2208);
   U2219 : OAI22_X1 port map( A1 => n2923, A2 => n2940, B1 => n3979, B2 => 
                           n2941, ZN => n2207);
   U2220 : OAI22_X1 port map( A1 => n2924, A2 => n2940, B1 => n3978, B2 => 
                           n2941, ZN => n2206);
   U2221 : OAI22_X1 port map( A1 => n2925, A2 => n2940, B1 => n3977, B2 => 
                           n2941, ZN => n2205);
   U2222 : OAI22_X1 port map( A1 => n2926, A2 => n2940, B1 => n3976, B2 => 
                           n2941, ZN => n2204);
   U2223 : OAI22_X1 port map( A1 => n2927, A2 => n2940, B1 => n3975, B2 => 
                           n2941, ZN => n2203);
   U2224 : OAI22_X1 port map( A1 => n2928, A2 => n2940, B1 => n3974, B2 => 
                           n2941, ZN => n2202);
   U2225 : OAI22_X1 port map( A1 => n2929, A2 => n2940, B1 => n3973, B2 => 
                           n2941, ZN => n2201);
   U2226 : OAI22_X1 port map( A1 => n2930, A2 => n2940, B1 => n3972, B2 => 
                           n2941, ZN => n2200);
   U2227 : OAI22_X1 port map( A1 => n2931, A2 => n2940, B1 => n3971, B2 => 
                           n2941, ZN => n2199);
   U2228 : OAI22_X1 port map( A1 => n2899, A2 => n2943, B1 => n3970, B2 => 
                           n2944, ZN => n2198);
   U2229 : OAI22_X1 port map( A1 => n2901, A2 => n2943, B1 => n3969, B2 => 
                           n2944, ZN => n2197);
   U2230 : OAI22_X1 port map( A1 => n2902, A2 => n2943, B1 => n3968, B2 => 
                           n2944, ZN => n2196);
   U2231 : OAI22_X1 port map( A1 => n2903, A2 => n2943, B1 => n3967, B2 => 
                           n2944, ZN => n2195);
   U2232 : OAI22_X1 port map( A1 => n2904, A2 => n2943, B1 => n3966, B2 => 
                           n2944, ZN => n2194);
   U2233 : OAI22_X1 port map( A1 => n2905, A2 => n2943, B1 => n3965, B2 => 
                           n2944, ZN => n2193);
   U2234 : OAI22_X1 port map( A1 => n2906, A2 => n2943, B1 => n3964, B2 => 
                           n2944, ZN => n2192);
   U2235 : OAI22_X1 port map( A1 => n2907, A2 => n2943, B1 => n3963, B2 => 
                           n2944, ZN => n2191);
   U2236 : OAI22_X1 port map( A1 => n2908, A2 => n2943, B1 => n3962, B2 => 
                           n2944, ZN => n2190);
   U2237 : OAI22_X1 port map( A1 => n2909, A2 => n2943, B1 => n3961, B2 => 
                           n2944, ZN => n2189);
   U2238 : OAI22_X1 port map( A1 => n2910, A2 => n2943, B1 => n3960, B2 => 
                           n2944, ZN => n2188);
   U2239 : OAI22_X1 port map( A1 => n2911, A2 => n2943, B1 => n3959, B2 => 
                           n2944, ZN => n2187);
   U2240 : OAI22_X1 port map( A1 => n2912, A2 => n2943, B1 => n3958, B2 => 
                           n2944, ZN => n2186);
   U2241 : OAI22_X1 port map( A1 => n2913, A2 => n2943, B1 => n3957, B2 => 
                           n2944, ZN => n2185);
   U2242 : OAI22_X1 port map( A1 => n2914, A2 => n2943, B1 => n3956, B2 => 
                           n2944, ZN => n2184);
   U2243 : OAI22_X1 port map( A1 => n2915, A2 => n2943, B1 => n3955, B2 => 
                           n2944, ZN => n2183);
   U2244 : OAI22_X1 port map( A1 => n2916, A2 => n2943, B1 => n3954, B2 => 
                           n2944, ZN => n2182);
   U2245 : OAI22_X1 port map( A1 => n2917, A2 => n2943, B1 => n3953, B2 => 
                           n2944, ZN => n2181);
   U2246 : OAI22_X1 port map( A1 => n2918, A2 => n2943, B1 => n3952, B2 => 
                           n2944, ZN => n2180);
   U2247 : OAI22_X1 port map( A1 => n2919, A2 => n2943, B1 => n3951, B2 => 
                           n2944, ZN => n2179);
   U2248 : OAI22_X1 port map( A1 => n2920, A2 => n2943, B1 => n3950, B2 => 
                           n2944, ZN => n2178);
   U2249 : OAI22_X1 port map( A1 => n2921, A2 => n2943, B1 => n3949, B2 => 
                           n2944, ZN => n2177);
   U2250 : OAI22_X1 port map( A1 => n2922, A2 => n2943, B1 => n3948, B2 => 
                           n2944, ZN => n2176);
   U2251 : OAI22_X1 port map( A1 => n2923, A2 => n2943, B1 => n3947, B2 => 
                           n2944, ZN => n2175);
   U2252 : OAI22_X1 port map( A1 => n2924, A2 => n2943, B1 => n3946, B2 => 
                           n2944, ZN => n2174);
   U2253 : OAI22_X1 port map( A1 => n2925, A2 => n2943, B1 => n3945, B2 => 
                           n2944, ZN => n2173);
   U2254 : OAI22_X1 port map( A1 => n2926, A2 => n2943, B1 => n3944, B2 => 
                           n2944, ZN => n2172);
   U2255 : OAI22_X1 port map( A1 => n2927, A2 => n2943, B1 => n3943, B2 => 
                           n2944, ZN => n2171);
   U2256 : OAI22_X1 port map( A1 => n2928, A2 => n2943, B1 => n3942, B2 => 
                           n2944, ZN => n2170);
   U2257 : OAI22_X1 port map( A1 => n2929, A2 => n2943, B1 => n3941, B2 => 
                           n2944, ZN => n2169);
   U2258 : OAI22_X1 port map( A1 => n2930, A2 => n2943, B1 => n3940, B2 => 
                           n2944, ZN => n2168);
   U2259 : OAI22_X1 port map( A1 => n2931, A2 => n2943, B1 => n3939, B2 => 
                           n2944, ZN => n2167);
   U2260 : OAI22_X1 port map( A1 => n2899, A2 => n2946, B1 => n3938, B2 => 
                           n2947, ZN => n2166);
   U2261 : OAI22_X1 port map( A1 => n2901, A2 => n2946, B1 => n3937, B2 => 
                           n2947, ZN => n2165);
   U2262 : OAI22_X1 port map( A1 => n2902, A2 => n2946, B1 => n3936, B2 => 
                           n2947, ZN => n2164);
   U2263 : OAI22_X1 port map( A1 => n2903, A2 => n2946, B1 => n3935, B2 => 
                           n2947, ZN => n2163);
   U2264 : OAI22_X1 port map( A1 => n2904, A2 => n2946, B1 => n3934, B2 => 
                           n2947, ZN => n2162);
   U2265 : OAI22_X1 port map( A1 => n2905, A2 => n2946, B1 => n3933, B2 => 
                           n2947, ZN => n2161);
   U2266 : OAI22_X1 port map( A1 => n2906, A2 => n2946, B1 => n3932, B2 => 
                           n2947, ZN => n2160);
   U2267 : OAI22_X1 port map( A1 => n2907, A2 => n2946, B1 => n3931, B2 => 
                           n2947, ZN => n2159);
   U2268 : OAI22_X1 port map( A1 => n2908, A2 => n2946, B1 => n3930, B2 => 
                           n2947, ZN => n2158);
   U2269 : OAI22_X1 port map( A1 => n2909, A2 => n2946, B1 => n3929, B2 => 
                           n2947, ZN => n2157);
   U2270 : OAI22_X1 port map( A1 => n2910, A2 => n2946, B1 => n3928, B2 => 
                           n2947, ZN => n2156);
   U2271 : OAI22_X1 port map( A1 => n2911, A2 => n2946, B1 => n3927, B2 => 
                           n2947, ZN => n2155);
   U2272 : OAI22_X1 port map( A1 => n2912, A2 => n2946, B1 => n3926, B2 => 
                           n2947, ZN => n2154);
   U2273 : OAI22_X1 port map( A1 => n2913, A2 => n2946, B1 => n3925, B2 => 
                           n2947, ZN => n2153);
   U2274 : OAI22_X1 port map( A1 => n2914, A2 => n2946, B1 => n3924, B2 => 
                           n2947, ZN => n2152);
   U2275 : OAI22_X1 port map( A1 => n2915, A2 => n2946, B1 => n3923, B2 => 
                           n2947, ZN => n2151);
   U2276 : OAI22_X1 port map( A1 => n2916, A2 => n2946, B1 => n3922, B2 => 
                           n2947, ZN => n2150);
   U2277 : OAI22_X1 port map( A1 => n2917, A2 => n2946, B1 => n3921, B2 => 
                           n2947, ZN => n2149);
   U2278 : OAI22_X1 port map( A1 => n2918, A2 => n2946, B1 => n3920, B2 => 
                           n2947, ZN => n2148);
   U2279 : OAI22_X1 port map( A1 => n2919, A2 => n2946, B1 => n3919, B2 => 
                           n2947, ZN => n2147);
   U2280 : OAI22_X1 port map( A1 => n2920, A2 => n2946, B1 => n3918, B2 => 
                           n2947, ZN => n2146);
   U2281 : OAI22_X1 port map( A1 => n2921, A2 => n2946, B1 => n3917, B2 => 
                           n2947, ZN => n2145);
   U2282 : OAI22_X1 port map( A1 => n2922, A2 => n2946, B1 => n3916, B2 => 
                           n2947, ZN => n2144);
   U2283 : OAI22_X1 port map( A1 => n2923, A2 => n2946, B1 => n3915, B2 => 
                           n2947, ZN => n2143);
   U2284 : OAI22_X1 port map( A1 => n2924, A2 => n2946, B1 => n3914, B2 => 
                           n2947, ZN => n2142);
   U2285 : OAI22_X1 port map( A1 => n2925, A2 => n2946, B1 => n3913, B2 => 
                           n2947, ZN => n2141);
   U2286 : OAI22_X1 port map( A1 => n2926, A2 => n2946, B1 => n3912, B2 => 
                           n2947, ZN => n2140);
   U2287 : OAI22_X1 port map( A1 => n2927, A2 => n2946, B1 => n3911, B2 => 
                           n2947, ZN => n2139);
   U2288 : OAI22_X1 port map( A1 => n2928, A2 => n2946, B1 => n3910, B2 => 
                           n2947, ZN => n2138);
   U2289 : OAI22_X1 port map( A1 => n2929, A2 => n2946, B1 => n3909, B2 => 
                           n2947, ZN => n2137);
   U2290 : OAI22_X1 port map( A1 => n2930, A2 => n2946, B1 => n3908, B2 => 
                           n2947, ZN => n2136);
   U2291 : OAI22_X1 port map( A1 => n2931, A2 => n2946, B1 => n3907, B2 => 
                           n2947, ZN => n2135);
   U2292 : OAI22_X1 port map( A1 => n2899, A2 => n2949, B1 => n3906, B2 => 
                           n2950, ZN => n2134);
   U2293 : OAI22_X1 port map( A1 => n2901, A2 => n2949, B1 => n3905, B2 => 
                           n2950, ZN => n2133);
   U2294 : OAI22_X1 port map( A1 => n2902, A2 => n2949, B1 => n3904, B2 => 
                           n2950, ZN => n2132);
   U2295 : OAI22_X1 port map( A1 => n2903, A2 => n2949, B1 => n3903, B2 => 
                           n2950, ZN => n2131);
   U2296 : OAI22_X1 port map( A1 => n2904, A2 => n2949, B1 => n3902, B2 => 
                           n2950, ZN => n2130);
   U2297 : OAI22_X1 port map( A1 => n2905, A2 => n2949, B1 => n3901, B2 => 
                           n2950, ZN => n2129);
   U2298 : OAI22_X1 port map( A1 => n2906, A2 => n2949, B1 => n3900, B2 => 
                           n2950, ZN => n2128);
   U2299 : OAI22_X1 port map( A1 => n2907, A2 => n2949, B1 => n3899, B2 => 
                           n2950, ZN => n2127);
   U2300 : OAI22_X1 port map( A1 => n2908, A2 => n2949, B1 => n3898, B2 => 
                           n2950, ZN => n2126);
   U2301 : OAI22_X1 port map( A1 => n2909, A2 => n2949, B1 => n3897, B2 => 
                           n2950, ZN => n2125);
   U2302 : OAI22_X1 port map( A1 => n2910, A2 => n2949, B1 => n3896, B2 => 
                           n2950, ZN => n2124);
   U2303 : OAI22_X1 port map( A1 => n2911, A2 => n2949, B1 => n3895, B2 => 
                           n2950, ZN => n2123);
   U2304 : OAI22_X1 port map( A1 => n2912, A2 => n2949, B1 => n3894, B2 => 
                           n2950, ZN => n2122);
   U2305 : OAI22_X1 port map( A1 => n2913, A2 => n2949, B1 => n3893, B2 => 
                           n2950, ZN => n2121);
   U2306 : OAI22_X1 port map( A1 => n2914, A2 => n2949, B1 => n3892, B2 => 
                           n2950, ZN => n2120);
   U2307 : OAI22_X1 port map( A1 => n2915, A2 => n2949, B1 => n3891, B2 => 
                           n2950, ZN => n2119);
   U2308 : OAI22_X1 port map( A1 => n2916, A2 => n2949, B1 => n3890, B2 => 
                           n2950, ZN => n2118);
   U2309 : OAI22_X1 port map( A1 => n2917, A2 => n2949, B1 => n3889, B2 => 
                           n2950, ZN => n2117);
   U2310 : OAI22_X1 port map( A1 => n2918, A2 => n2949, B1 => n3888, B2 => 
                           n2950, ZN => n2116);
   U2311 : OAI22_X1 port map( A1 => n2919, A2 => n2949, B1 => n3887, B2 => 
                           n2950, ZN => n2115);
   U2312 : OAI22_X1 port map( A1 => n2920, A2 => n2949, B1 => n3886, B2 => 
                           n2950, ZN => n2114);
   U2313 : OAI22_X1 port map( A1 => n2921, A2 => n2949, B1 => n3885, B2 => 
                           n2950, ZN => n2113);
   U2314 : OAI22_X1 port map( A1 => n2922, A2 => n2949, B1 => n3884, B2 => 
                           n2950, ZN => n2112);
   U2315 : OAI22_X1 port map( A1 => n2923, A2 => n2949, B1 => n3883, B2 => 
                           n2950, ZN => n2111);
   U2316 : OAI22_X1 port map( A1 => n2924, A2 => n2949, B1 => n3882, B2 => 
                           n2950, ZN => n2110);
   U2317 : OAI22_X1 port map( A1 => n2925, A2 => n2949, B1 => n3881, B2 => 
                           n2950, ZN => n2109);
   U2318 : OAI22_X1 port map( A1 => n2926, A2 => n2949, B1 => n3880, B2 => 
                           n2950, ZN => n2108);
   U2319 : OAI22_X1 port map( A1 => n2927, A2 => n2949, B1 => n3879, B2 => 
                           n2950, ZN => n2107);
   U2320 : OAI22_X1 port map( A1 => n2928, A2 => n2949, B1 => n3878, B2 => 
                           n2950, ZN => n2106);
   U2321 : OAI22_X1 port map( A1 => n2929, A2 => n2949, B1 => n3877, B2 => 
                           n2950, ZN => n2105);
   U2322 : OAI22_X1 port map( A1 => n2930, A2 => n2949, B1 => n3876, B2 => 
                           n2950, ZN => n2104);
   U2323 : OAI22_X1 port map( A1 => n2931, A2 => n2949, B1 => n3875, B2 => 
                           n2950, ZN => n2103);
   U2324 : OAI22_X1 port map( A1 => n2899, A2 => n2952, B1 => n3874, B2 => 
                           n2953, ZN => n2102);
   U2325 : OAI22_X1 port map( A1 => n2901, A2 => n2952, B1 => n3873, B2 => 
                           n2953, ZN => n2101);
   U2326 : OAI22_X1 port map( A1 => n2902, A2 => n2952, B1 => n3872, B2 => 
                           n2953, ZN => n2100);
   U2327 : OAI22_X1 port map( A1 => n2903, A2 => n2952, B1 => n3871, B2 => 
                           n2953, ZN => n2099);
   U2328 : OAI22_X1 port map( A1 => n2904, A2 => n2952, B1 => n3870, B2 => 
                           n2953, ZN => n2098);
   U2329 : OAI22_X1 port map( A1 => n2905, A2 => n2952, B1 => n3869, B2 => 
                           n2953, ZN => n2097);
   U2330 : OAI22_X1 port map( A1 => n2906, A2 => n2952, B1 => n3868, B2 => 
                           n2953, ZN => n2096);
   U2331 : OAI22_X1 port map( A1 => n2907, A2 => n2952, B1 => n3867, B2 => 
                           n2953, ZN => n2095);
   U2332 : OAI22_X1 port map( A1 => n2908, A2 => n2952, B1 => n3866, B2 => 
                           n2953, ZN => n2094);
   U2333 : OAI22_X1 port map( A1 => n2909, A2 => n2952, B1 => n3865, B2 => 
                           n2953, ZN => n2093);
   U2334 : OAI22_X1 port map( A1 => n2910, A2 => n2952, B1 => n3864, B2 => 
                           n2953, ZN => n2092);
   U2335 : OAI22_X1 port map( A1 => n2911, A2 => n2952, B1 => n3863, B2 => 
                           n2953, ZN => n2091);
   U2336 : OAI22_X1 port map( A1 => n2912, A2 => n2952, B1 => n3862, B2 => 
                           n2953, ZN => n2090);
   U2337 : OAI22_X1 port map( A1 => n2913, A2 => n2952, B1 => n3861, B2 => 
                           n2953, ZN => n2089);
   U2338 : OAI22_X1 port map( A1 => n2914, A2 => n2952, B1 => n3860, B2 => 
                           n2953, ZN => n2088);
   U2339 : OAI22_X1 port map( A1 => n2915, A2 => n2952, B1 => n3859, B2 => 
                           n2953, ZN => n2087);
   U2340 : OAI22_X1 port map( A1 => n2916, A2 => n2952, B1 => n3858, B2 => 
                           n2953, ZN => n2086);
   U2341 : OAI22_X1 port map( A1 => n2917, A2 => n2952, B1 => n3857, B2 => 
                           n2953, ZN => n2085);
   U2342 : OAI22_X1 port map( A1 => n2918, A2 => n2952, B1 => n3856, B2 => 
                           n2953, ZN => n2084);
   U2343 : OAI22_X1 port map( A1 => n2919, A2 => n2952, B1 => n3855, B2 => 
                           n2953, ZN => n2083);
   U2344 : OAI22_X1 port map( A1 => n2920, A2 => n2952, B1 => n3854, B2 => 
                           n2953, ZN => n2082);
   U2345 : OAI22_X1 port map( A1 => n2921, A2 => n2952, B1 => n3853, B2 => 
                           n2953, ZN => n2081);
   U2346 : OAI22_X1 port map( A1 => n2922, A2 => n2952, B1 => n3852, B2 => 
                           n2953, ZN => n2080);
   U2347 : OAI22_X1 port map( A1 => n2923, A2 => n2952, B1 => n3851, B2 => 
                           n2953, ZN => n2079);
   U2348 : OAI22_X1 port map( A1 => n2924, A2 => n2952, B1 => n3850, B2 => 
                           n2953, ZN => n2078);
   U2349 : OAI22_X1 port map( A1 => n2925, A2 => n2952, B1 => n3849, B2 => 
                           n2953, ZN => n2077);
   U2350 : OAI22_X1 port map( A1 => n2926, A2 => n2952, B1 => n3848, B2 => 
                           n2953, ZN => n2076);
   U2351 : OAI22_X1 port map( A1 => n2927, A2 => n2952, B1 => n3847, B2 => 
                           n2953, ZN => n2075);
   U2352 : OAI22_X1 port map( A1 => n2928, A2 => n2952, B1 => n3846, B2 => 
                           n2953, ZN => n2074);
   U2353 : OAI22_X1 port map( A1 => n2929, A2 => n2952, B1 => n3845, B2 => 
                           n2953, ZN => n2073);
   U2354 : OAI22_X1 port map( A1 => n2930, A2 => n2952, B1 => n3844, B2 => 
                           n2953, ZN => n2072);
   U2355 : OAI22_X1 port map( A1 => n2931, A2 => n2952, B1 => n3843, B2 => 
                           n2953, ZN => n2071);
   U2356 : AND3_X1 port map( A1 => n2955, A2 => n2956, A3 => n2957, ZN => n2933
                           );
   U2357 : OAI22_X1 port map( A1 => n2899, A2 => n2958, B1 => n3842, B2 => 
                           n2959, ZN => n2070);
   U2358 : OAI22_X1 port map( A1 => n2901, A2 => n2958, B1 => n3841, B2 => 
                           n2959, ZN => n2069);
   U2359 : OAI22_X1 port map( A1 => n2902, A2 => n2958, B1 => n3840, B2 => 
                           n2959, ZN => n2068);
   U2360 : OAI22_X1 port map( A1 => n2903, A2 => n2958, B1 => n3839, B2 => 
                           n2959, ZN => n2067);
   U2361 : OAI22_X1 port map( A1 => n2904, A2 => n2958, B1 => n3838, B2 => 
                           n2959, ZN => n2066);
   U2362 : OAI22_X1 port map( A1 => n2905, A2 => n2958, B1 => n3837, B2 => 
                           n2959, ZN => n2065);
   U2363 : OAI22_X1 port map( A1 => n2906, A2 => n2958, B1 => n3836, B2 => 
                           n2959, ZN => n2064);
   U2364 : OAI22_X1 port map( A1 => n2907, A2 => n2958, B1 => n3835, B2 => 
                           n2959, ZN => n2063);
   U2365 : OAI22_X1 port map( A1 => n2908, A2 => n2958, B1 => n3834, B2 => 
                           n2959, ZN => n2062);
   U2366 : OAI22_X1 port map( A1 => n2909, A2 => n2958, B1 => n3833, B2 => 
                           n2959, ZN => n2061);
   U2367 : OAI22_X1 port map( A1 => n2910, A2 => n2958, B1 => n3832, B2 => 
                           n2959, ZN => n2060);
   U2368 : OAI22_X1 port map( A1 => n2911, A2 => n2958, B1 => n3831, B2 => 
                           n2959, ZN => n2059);
   U2369 : OAI22_X1 port map( A1 => n2912, A2 => n2958, B1 => n3830, B2 => 
                           n2959, ZN => n2058);
   U2370 : OAI22_X1 port map( A1 => n2913, A2 => n2958, B1 => n3829, B2 => 
                           n2959, ZN => n2057);
   U2371 : OAI22_X1 port map( A1 => n2914, A2 => n2958, B1 => n3828, B2 => 
                           n2959, ZN => n2056);
   U2372 : OAI22_X1 port map( A1 => n2915, A2 => n2958, B1 => n3827, B2 => 
                           n2959, ZN => n2055);
   U2373 : OAI22_X1 port map( A1 => n2916, A2 => n2958, B1 => n3826, B2 => 
                           n2959, ZN => n2054);
   U2374 : OAI22_X1 port map( A1 => n2917, A2 => n2958, B1 => n3825, B2 => 
                           n2959, ZN => n2053);
   U2375 : OAI22_X1 port map( A1 => n2918, A2 => n2958, B1 => n3824, B2 => 
                           n2959, ZN => n2052);
   U2376 : OAI22_X1 port map( A1 => n2919, A2 => n2958, B1 => n3823, B2 => 
                           n2959, ZN => n2051);
   U2377 : OAI22_X1 port map( A1 => n2920, A2 => n2958, B1 => n3822, B2 => 
                           n2959, ZN => n2050);
   U2378 : OAI22_X1 port map( A1 => n2921, A2 => n2958, B1 => n3821, B2 => 
                           n2959, ZN => n2049);
   U2379 : OAI22_X1 port map( A1 => n2922, A2 => n2958, B1 => n3820, B2 => 
                           n2959, ZN => n2048);
   U2380 : OAI22_X1 port map( A1 => n2923, A2 => n2958, B1 => n3819, B2 => 
                           n2959, ZN => n2047);
   U2381 : OAI22_X1 port map( A1 => n2924, A2 => n2958, B1 => n3818, B2 => 
                           n2959, ZN => n2046);
   U2382 : OAI22_X1 port map( A1 => n2925, A2 => n2958, B1 => n3817, B2 => 
                           n2959, ZN => n2045);
   U2383 : OAI22_X1 port map( A1 => n2926, A2 => n2958, B1 => n3816, B2 => 
                           n2959, ZN => n2044);
   U2384 : OAI22_X1 port map( A1 => n2927, A2 => n2958, B1 => n3815, B2 => 
                           n2959, ZN => n2043);
   U2385 : OAI22_X1 port map( A1 => n2928, A2 => n2958, B1 => n3814, B2 => 
                           n2959, ZN => n2042);
   U2386 : OAI22_X1 port map( A1 => n2929, A2 => n2958, B1 => n3813, B2 => 
                           n2959, ZN => n2041);
   U2387 : OAI22_X1 port map( A1 => n2930, A2 => n2958, B1 => n3812, B2 => 
                           n2959, ZN => n2040);
   U2388 : OAI22_X1 port map( A1 => n2931, A2 => n2958, B1 => n3811, B2 => 
                           n2959, ZN => n2039);
   U2389 : OAI22_X1 port map( A1 => n2899, A2 => n2961, B1 => n3810, B2 => 
                           n2962, ZN => n2038);
   U2390 : OAI22_X1 port map( A1 => n2901, A2 => n2961, B1 => n3809, B2 => 
                           n2962, ZN => n2037);
   U2391 : OAI22_X1 port map( A1 => n2902, A2 => n2961, B1 => n3808, B2 => 
                           n2962, ZN => n2036);
   U2392 : OAI22_X1 port map( A1 => n2903, A2 => n2961, B1 => n3807, B2 => 
                           n2962, ZN => n2035);
   U2393 : OAI22_X1 port map( A1 => n2904, A2 => n2961, B1 => n3806, B2 => 
                           n2962, ZN => n2034);
   U2394 : OAI22_X1 port map( A1 => n2905, A2 => n2961, B1 => n3805, B2 => 
                           n2962, ZN => n2033);
   U2395 : OAI22_X1 port map( A1 => n2906, A2 => n2961, B1 => n3804, B2 => 
                           n2962, ZN => n2032);
   U2396 : OAI22_X1 port map( A1 => n2907, A2 => n2961, B1 => n3803, B2 => 
                           n2962, ZN => n2031);
   U2397 : OAI22_X1 port map( A1 => n2908, A2 => n2961, B1 => n3802, B2 => 
                           n2962, ZN => n2030);
   U2398 : OAI22_X1 port map( A1 => n2909, A2 => n2961, B1 => n3801, B2 => 
                           n2962, ZN => n2029);
   U2399 : OAI22_X1 port map( A1 => n2910, A2 => n2961, B1 => n3800, B2 => 
                           n2962, ZN => n2028);
   U2400 : OAI22_X1 port map( A1 => n2911, A2 => n2961, B1 => n3799, B2 => 
                           n2962, ZN => n2027);
   U2401 : OAI22_X1 port map( A1 => n2912, A2 => n2961, B1 => n3798, B2 => 
                           n2962, ZN => n2026);
   U2402 : OAI22_X1 port map( A1 => n2913, A2 => n2961, B1 => n3797, B2 => 
                           n2962, ZN => n2025);
   U2403 : OAI22_X1 port map( A1 => n2914, A2 => n2961, B1 => n3796, B2 => 
                           n2962, ZN => n2024);
   U2404 : OAI22_X1 port map( A1 => n2915, A2 => n2961, B1 => n3795, B2 => 
                           n2962, ZN => n2023);
   U2405 : OAI22_X1 port map( A1 => n2916, A2 => n2961, B1 => n3794, B2 => 
                           n2962, ZN => n2022);
   U2406 : OAI22_X1 port map( A1 => n2917, A2 => n2961, B1 => n3793, B2 => 
                           n2962, ZN => n2021);
   U2407 : OAI22_X1 port map( A1 => n2918, A2 => n2961, B1 => n3792, B2 => 
                           n2962, ZN => n2020);
   U2408 : OAI22_X1 port map( A1 => n2919, A2 => n2961, B1 => n3791, B2 => 
                           n2962, ZN => n2019);
   U2409 : OAI22_X1 port map( A1 => n2920, A2 => n2961, B1 => n3790, B2 => 
                           n2962, ZN => n2018);
   U2410 : OAI22_X1 port map( A1 => n2921, A2 => n2961, B1 => n3789, B2 => 
                           n2962, ZN => n2017);
   U2411 : OAI22_X1 port map( A1 => n2922, A2 => n2961, B1 => n3788, B2 => 
                           n2962, ZN => n2016);
   U2412 : OAI22_X1 port map( A1 => n2923, A2 => n2961, B1 => n3787, B2 => 
                           n2962, ZN => n2015);
   U2413 : OAI22_X1 port map( A1 => n2924, A2 => n2961, B1 => n3786, B2 => 
                           n2962, ZN => n2014);
   U2414 : OAI22_X1 port map( A1 => n2925, A2 => n2961, B1 => n3785, B2 => 
                           n2962, ZN => n2013);
   U2415 : OAI22_X1 port map( A1 => n2926, A2 => n2961, B1 => n3784, B2 => 
                           n2962, ZN => n2012);
   U2416 : OAI22_X1 port map( A1 => n2927, A2 => n2961, B1 => n3783, B2 => 
                           n2962, ZN => n2011);
   U2417 : OAI22_X1 port map( A1 => n2928, A2 => n2961, B1 => n3782, B2 => 
                           n2962, ZN => n2010);
   U2418 : OAI22_X1 port map( A1 => n2929, A2 => n2961, B1 => n3781, B2 => 
                           n2962, ZN => n2009);
   U2419 : OAI22_X1 port map( A1 => n2930, A2 => n2961, B1 => n3780, B2 => 
                           n2962, ZN => n2008);
   U2420 : OAI22_X1 port map( A1 => n2931, A2 => n2961, B1 => n3779, B2 => 
                           n2962, ZN => n2007);
   U2421 : OAI22_X1 port map( A1 => n2899, A2 => n2963, B1 => n3778, B2 => 
                           n2964, ZN => n2006);
   U2422 : OAI22_X1 port map( A1 => n2901, A2 => n2963, B1 => n3777, B2 => 
                           n2964, ZN => n2005);
   U2423 : OAI22_X1 port map( A1 => n2902, A2 => n2963, B1 => n3776, B2 => 
                           n2964, ZN => n2004);
   U2424 : OAI22_X1 port map( A1 => n2903, A2 => n2963, B1 => n3775, B2 => 
                           n2964, ZN => n2003);
   U2425 : OAI22_X1 port map( A1 => n2904, A2 => n2963, B1 => n3774, B2 => 
                           n2964, ZN => n2002);
   U2426 : OAI22_X1 port map( A1 => n2905, A2 => n2963, B1 => n3773, B2 => 
                           n2964, ZN => n2001);
   U2427 : OAI22_X1 port map( A1 => n2906, A2 => n2963, B1 => n3772, B2 => 
                           n2964, ZN => n2000);
   U2428 : OAI22_X1 port map( A1 => n2907, A2 => n2963, B1 => n3771, B2 => 
                           n2964, ZN => n1999);
   U2429 : OAI22_X1 port map( A1 => n2908, A2 => n2963, B1 => n3770, B2 => 
                           n2964, ZN => n1998);
   U2430 : OAI22_X1 port map( A1 => n2909, A2 => n2963, B1 => n3769, B2 => 
                           n2964, ZN => n1997);
   U2431 : OAI22_X1 port map( A1 => n2910, A2 => n2963, B1 => n3768, B2 => 
                           n2964, ZN => n1996);
   U2432 : OAI22_X1 port map( A1 => n2911, A2 => n2963, B1 => n3767, B2 => 
                           n2964, ZN => n1995);
   U2433 : OAI22_X1 port map( A1 => n2912, A2 => n2963, B1 => n3766, B2 => 
                           n2964, ZN => n1994);
   U2434 : OAI22_X1 port map( A1 => n2913, A2 => n2963, B1 => n3765, B2 => 
                           n2964, ZN => n1993);
   U2435 : OAI22_X1 port map( A1 => n2914, A2 => n2963, B1 => n3764, B2 => 
                           n2964, ZN => n1992);
   U2436 : OAI22_X1 port map( A1 => n2915, A2 => n2963, B1 => n3763, B2 => 
                           n2964, ZN => n1991);
   U2437 : OAI22_X1 port map( A1 => n2916, A2 => n2963, B1 => n3762, B2 => 
                           n2964, ZN => n1990);
   U2438 : OAI22_X1 port map( A1 => n2917, A2 => n2963, B1 => n3761, B2 => 
                           n2964, ZN => n1989);
   U2439 : OAI22_X1 port map( A1 => n2918, A2 => n2963, B1 => n3760, B2 => 
                           n2964, ZN => n1988);
   U2440 : OAI22_X1 port map( A1 => n2919, A2 => n2963, B1 => n3759, B2 => 
                           n2964, ZN => n1987);
   U2441 : OAI22_X1 port map( A1 => n2920, A2 => n2963, B1 => n3758, B2 => 
                           n2964, ZN => n1986);
   U2442 : OAI22_X1 port map( A1 => n2921, A2 => n2963, B1 => n3757, B2 => 
                           n2964, ZN => n1985);
   U2443 : OAI22_X1 port map( A1 => n2922, A2 => n2963, B1 => n3756, B2 => 
                           n2964, ZN => n1984);
   U2444 : OAI22_X1 port map( A1 => n2923, A2 => n2963, B1 => n3755, B2 => 
                           n2964, ZN => n1983);
   U2445 : OAI22_X1 port map( A1 => n2924, A2 => n2963, B1 => n3754, B2 => 
                           n2964, ZN => n1982);
   U2446 : OAI22_X1 port map( A1 => n2925, A2 => n2963, B1 => n3753, B2 => 
                           n2964, ZN => n1981);
   U2447 : OAI22_X1 port map( A1 => n2926, A2 => n2963, B1 => n3752, B2 => 
                           n2964, ZN => n1980);
   U2448 : OAI22_X1 port map( A1 => n2927, A2 => n2963, B1 => n3751, B2 => 
                           n2964, ZN => n1979);
   U2449 : OAI22_X1 port map( A1 => n2928, A2 => n2963, B1 => n3750, B2 => 
                           n2964, ZN => n1978);
   U2450 : OAI22_X1 port map( A1 => n2929, A2 => n2963, B1 => n3749, B2 => 
                           n2964, ZN => n1977);
   U2451 : OAI22_X1 port map( A1 => n2930, A2 => n2963, B1 => n3748, B2 => 
                           n2964, ZN => n1976);
   U2452 : OAI22_X1 port map( A1 => n2931, A2 => n2963, B1 => n3747, B2 => 
                           n2964, ZN => n1975);
   U2453 : OAI22_X1 port map( A1 => n2899, A2 => n2965, B1 => n3746, B2 => 
                           n2966, ZN => n1974);
   U2454 : OAI22_X1 port map( A1 => n2901, A2 => n2965, B1 => n3745, B2 => 
                           n2966, ZN => n1973);
   U2455 : OAI22_X1 port map( A1 => n2902, A2 => n2965, B1 => n3744, B2 => 
                           n2966, ZN => n1972);
   U2456 : OAI22_X1 port map( A1 => n2903, A2 => n2965, B1 => n3743, B2 => 
                           n2966, ZN => n1971);
   U2457 : OAI22_X1 port map( A1 => n2904, A2 => n2965, B1 => n3742, B2 => 
                           n2966, ZN => n1970);
   U2458 : OAI22_X1 port map( A1 => n2905, A2 => n2965, B1 => n3741, B2 => 
                           n2966, ZN => n1969);
   U2459 : OAI22_X1 port map( A1 => n2906, A2 => n2965, B1 => n3740, B2 => 
                           n2966, ZN => n1968);
   U2460 : OAI22_X1 port map( A1 => n2907, A2 => n2965, B1 => n3739, B2 => 
                           n2966, ZN => n1967);
   U2461 : OAI22_X1 port map( A1 => n2908, A2 => n2965, B1 => n3738, B2 => 
                           n2966, ZN => n1966);
   U2462 : OAI22_X1 port map( A1 => n2909, A2 => n2965, B1 => n3737, B2 => 
                           n2966, ZN => n1965);
   U2463 : OAI22_X1 port map( A1 => n2910, A2 => n2965, B1 => n3736, B2 => 
                           n2966, ZN => n1964);
   U2464 : OAI22_X1 port map( A1 => n2911, A2 => n2965, B1 => n3735, B2 => 
                           n2966, ZN => n1963);
   U2465 : OAI22_X1 port map( A1 => n2912, A2 => n2965, B1 => n3734, B2 => 
                           n2966, ZN => n1962);
   U2466 : OAI22_X1 port map( A1 => n2913, A2 => n2965, B1 => n3733, B2 => 
                           n2966, ZN => n1961);
   U2467 : OAI22_X1 port map( A1 => n2914, A2 => n2965, B1 => n3732, B2 => 
                           n2966, ZN => n1960);
   U2468 : OAI22_X1 port map( A1 => n2915, A2 => n2965, B1 => n3731, B2 => 
                           n2966, ZN => n1959);
   U2469 : OAI22_X1 port map( A1 => n2916, A2 => n2965, B1 => n3730, B2 => 
                           n2966, ZN => n1958);
   U2470 : OAI22_X1 port map( A1 => n2917, A2 => n2965, B1 => n3729, B2 => 
                           n2966, ZN => n1957);
   U2471 : OAI22_X1 port map( A1 => n2918, A2 => n2965, B1 => n3728, B2 => 
                           n2966, ZN => n1956);
   U2472 : OAI22_X1 port map( A1 => n2919, A2 => n2965, B1 => n3727, B2 => 
                           n2966, ZN => n1955);
   U2473 : OAI22_X1 port map( A1 => n2920, A2 => n2965, B1 => n3726, B2 => 
                           n2966, ZN => n1954);
   U2474 : OAI22_X1 port map( A1 => n2921, A2 => n2965, B1 => n3725, B2 => 
                           n2966, ZN => n1953);
   U2475 : OAI22_X1 port map( A1 => n2922, A2 => n2965, B1 => n3724, B2 => 
                           n2966, ZN => n1952);
   U2476 : OAI22_X1 port map( A1 => n2923, A2 => n2965, B1 => n3723, B2 => 
                           n2966, ZN => n1951);
   U2477 : OAI22_X1 port map( A1 => n2924, A2 => n2965, B1 => n3722, B2 => 
                           n2966, ZN => n1950);
   U2478 : OAI22_X1 port map( A1 => n2925, A2 => n2965, B1 => n3721, B2 => 
                           n2966, ZN => n1949);
   U2479 : OAI22_X1 port map( A1 => n2926, A2 => n2965, B1 => n3720, B2 => 
                           n2966, ZN => n1948);
   U2480 : OAI22_X1 port map( A1 => n2927, A2 => n2965, B1 => n3719, B2 => 
                           n2966, ZN => n1947);
   U2481 : OAI22_X1 port map( A1 => n2928, A2 => n2965, B1 => n3718, B2 => 
                           n2966, ZN => n1946);
   U2482 : OAI22_X1 port map( A1 => n2929, A2 => n2965, B1 => n3717, B2 => 
                           n2966, ZN => n1945);
   U2483 : OAI22_X1 port map( A1 => n2930, A2 => n2965, B1 => n3716, B2 => 
                           n2966, ZN => n1944);
   U2484 : OAI22_X1 port map( A1 => n2931, A2 => n2965, B1 => n3715, B2 => 
                           n2966, ZN => n1943);
   U2485 : OAI22_X1 port map( A1 => n2899, A2 => n2967, B1 => n3714, B2 => 
                           n2968, ZN => n1942);
   U2486 : OAI22_X1 port map( A1 => n2901, A2 => n2967, B1 => n3713, B2 => 
                           n2968, ZN => n1941);
   U2487 : OAI22_X1 port map( A1 => n2902, A2 => n2967, B1 => n3712, B2 => 
                           n2968, ZN => n1940);
   U2488 : OAI22_X1 port map( A1 => n2903, A2 => n2967, B1 => n3711, B2 => 
                           n2968, ZN => n1939);
   U2489 : OAI22_X1 port map( A1 => n2904, A2 => n2967, B1 => n3710, B2 => 
                           n2968, ZN => n1938);
   U2490 : OAI22_X1 port map( A1 => n2905, A2 => n2967, B1 => n3709, B2 => 
                           n2968, ZN => n1937);
   U2491 : OAI22_X1 port map( A1 => n2906, A2 => n2967, B1 => n3708, B2 => 
                           n2968, ZN => n1936);
   U2492 : OAI22_X1 port map( A1 => n2907, A2 => n2967, B1 => n3707, B2 => 
                           n2968, ZN => n1935);
   U2493 : OAI22_X1 port map( A1 => n2908, A2 => n2967, B1 => n3706, B2 => 
                           n2968, ZN => n1934);
   U2494 : OAI22_X1 port map( A1 => n2909, A2 => n2967, B1 => n3705, B2 => 
                           n2968, ZN => n1933);
   U2495 : OAI22_X1 port map( A1 => n2910, A2 => n2967, B1 => n3704, B2 => 
                           n2968, ZN => n1932);
   U2496 : OAI22_X1 port map( A1 => n2911, A2 => n2967, B1 => n3703, B2 => 
                           n2968, ZN => n1931);
   U2497 : OAI22_X1 port map( A1 => n2912, A2 => n2967, B1 => n3702, B2 => 
                           n2968, ZN => n1930);
   U2498 : OAI22_X1 port map( A1 => n2913, A2 => n2967, B1 => n3701, B2 => 
                           n2968, ZN => n1929);
   U2499 : OAI22_X1 port map( A1 => n2914, A2 => n2967, B1 => n3700, B2 => 
                           n2968, ZN => n1928);
   U2500 : OAI22_X1 port map( A1 => n2915, A2 => n2967, B1 => n3699, B2 => 
                           n2968, ZN => n1927);
   U2501 : OAI22_X1 port map( A1 => n2916, A2 => n2967, B1 => n3698, B2 => 
                           n2968, ZN => n1926);
   U2502 : OAI22_X1 port map( A1 => n2917, A2 => n2967, B1 => n3697, B2 => 
                           n2968, ZN => n1925);
   U2503 : OAI22_X1 port map( A1 => n2918, A2 => n2967, B1 => n3696, B2 => 
                           n2968, ZN => n1924);
   U2504 : OAI22_X1 port map( A1 => n2919, A2 => n2967, B1 => n3695, B2 => 
                           n2968, ZN => n1923);
   U2505 : OAI22_X1 port map( A1 => n2920, A2 => n2967, B1 => n3694, B2 => 
                           n2968, ZN => n1922);
   U2506 : OAI22_X1 port map( A1 => n2921, A2 => n2967, B1 => n3693, B2 => 
                           n2968, ZN => n1921);
   U2507 : OAI22_X1 port map( A1 => n2922, A2 => n2967, B1 => n3692, B2 => 
                           n2968, ZN => n1920);
   U2508 : OAI22_X1 port map( A1 => n2923, A2 => n2967, B1 => n3691, B2 => 
                           n2968, ZN => n1919);
   U2509 : OAI22_X1 port map( A1 => n2924, A2 => n2967, B1 => n3690, B2 => 
                           n2968, ZN => n1918);
   U2510 : OAI22_X1 port map( A1 => n2925, A2 => n2967, B1 => n3689, B2 => 
                           n2968, ZN => n1917);
   U2511 : OAI22_X1 port map( A1 => n2926, A2 => n2967, B1 => n3688, B2 => 
                           n2968, ZN => n1916);
   U2512 : OAI22_X1 port map( A1 => n2927, A2 => n2967, B1 => n3687, B2 => 
                           n2968, ZN => n1915);
   U2513 : OAI22_X1 port map( A1 => n2928, A2 => n2967, B1 => n3686, B2 => 
                           n2968, ZN => n1914);
   U2514 : OAI22_X1 port map( A1 => n2929, A2 => n2967, B1 => n3685, B2 => 
                           n2968, ZN => n1913);
   U2515 : OAI22_X1 port map( A1 => n2930, A2 => n2967, B1 => n3684, B2 => 
                           n2968, ZN => n1912);
   U2516 : OAI22_X1 port map( A1 => n2931, A2 => n2967, B1 => n3683, B2 => 
                           n2968, ZN => n1911);
   U2517 : OAI22_X1 port map( A1 => n2899, A2 => n2969, B1 => n3682, B2 => 
                           n2970, ZN => n1910);
   U2518 : OAI22_X1 port map( A1 => n2901, A2 => n2969, B1 => n3681, B2 => 
                           n2970, ZN => n1909);
   U2519 : OAI22_X1 port map( A1 => n2902, A2 => n2969, B1 => n3680, B2 => 
                           n2970, ZN => n1908);
   U2520 : OAI22_X1 port map( A1 => n2903, A2 => n2969, B1 => n3679, B2 => 
                           n2970, ZN => n1907);
   U2521 : OAI22_X1 port map( A1 => n2904, A2 => n2969, B1 => n3678, B2 => 
                           n2970, ZN => n1906);
   U2522 : OAI22_X1 port map( A1 => n2905, A2 => n2969, B1 => n3677, B2 => 
                           n2970, ZN => n1905);
   U2523 : OAI22_X1 port map( A1 => n2906, A2 => n2969, B1 => n3676, B2 => 
                           n2970, ZN => n1904);
   U2524 : OAI22_X1 port map( A1 => n2907, A2 => n2969, B1 => n3675, B2 => 
                           n2970, ZN => n1903);
   U2525 : OAI22_X1 port map( A1 => n2908, A2 => n2969, B1 => n3674, B2 => 
                           n2970, ZN => n1902);
   U2526 : OAI22_X1 port map( A1 => n2909, A2 => n2969, B1 => n3673, B2 => 
                           n2970, ZN => n1901);
   U2527 : OAI22_X1 port map( A1 => n2910, A2 => n2969, B1 => n3672, B2 => 
                           n2970, ZN => n1900);
   U2528 : OAI22_X1 port map( A1 => n2911, A2 => n2969, B1 => n3671, B2 => 
                           n2970, ZN => n1899);
   U2529 : OAI22_X1 port map( A1 => n2912, A2 => n2969, B1 => n3670, B2 => 
                           n2970, ZN => n1898);
   U2530 : OAI22_X1 port map( A1 => n2913, A2 => n2969, B1 => n3669, B2 => 
                           n2970, ZN => n1897);
   U2531 : OAI22_X1 port map( A1 => n2914, A2 => n2969, B1 => n3668, B2 => 
                           n2970, ZN => n1896);
   U2532 : OAI22_X1 port map( A1 => n2915, A2 => n2969, B1 => n3667, B2 => 
                           n2970, ZN => n1895);
   U2533 : OAI22_X1 port map( A1 => n2916, A2 => n2969, B1 => n3666, B2 => 
                           n2970, ZN => n1894);
   U2534 : OAI22_X1 port map( A1 => n2917, A2 => n2969, B1 => n3665, B2 => 
                           n2970, ZN => n1893);
   U2535 : OAI22_X1 port map( A1 => n2918, A2 => n2969, B1 => n3664, B2 => 
                           n2970, ZN => n1892);
   U2536 : OAI22_X1 port map( A1 => n2919, A2 => n2969, B1 => n3663, B2 => 
                           n2970, ZN => n1891);
   U2537 : OAI22_X1 port map( A1 => n2920, A2 => n2969, B1 => n3662, B2 => 
                           n2970, ZN => n1890);
   U2538 : OAI22_X1 port map( A1 => n2921, A2 => n2969, B1 => n3661, B2 => 
                           n2970, ZN => n1889);
   U2539 : OAI22_X1 port map( A1 => n2922, A2 => n2969, B1 => n3660, B2 => 
                           n2970, ZN => n1888);
   U2540 : OAI22_X1 port map( A1 => n2923, A2 => n2969, B1 => n3659, B2 => 
                           n2970, ZN => n1887);
   U2541 : OAI22_X1 port map( A1 => n2924, A2 => n2969, B1 => n3658, B2 => 
                           n2970, ZN => n1886);
   U2542 : OAI22_X1 port map( A1 => n2925, A2 => n2969, B1 => n3657, B2 => 
                           n2970, ZN => n1885);
   U2543 : OAI22_X1 port map( A1 => n2926, A2 => n2969, B1 => n3656, B2 => 
                           n2970, ZN => n1884);
   U2544 : OAI22_X1 port map( A1 => n2927, A2 => n2969, B1 => n3655, B2 => 
                           n2970, ZN => n1883);
   U2545 : OAI22_X1 port map( A1 => n2928, A2 => n2969, B1 => n3654, B2 => 
                           n2970, ZN => n1882);
   U2546 : OAI22_X1 port map( A1 => n2929, A2 => n2969, B1 => n3653, B2 => 
                           n2970, ZN => n1881);
   U2547 : OAI22_X1 port map( A1 => n2930, A2 => n2969, B1 => n3652, B2 => 
                           n2970, ZN => n1880);
   U2548 : OAI22_X1 port map( A1 => n2931, A2 => n2969, B1 => n3651, B2 => 
                           n2970, ZN => n1879);
   U2549 : OAI22_X1 port map( A1 => n2899, A2 => n2971, B1 => n3650, B2 => 
                           n2972, ZN => n1878);
   U2550 : OAI22_X1 port map( A1 => n2901, A2 => n2971, B1 => n3649, B2 => 
                           n2972, ZN => n1877);
   U2551 : OAI22_X1 port map( A1 => n2902, A2 => n2971, B1 => n3648, B2 => 
                           n2972, ZN => n1876);
   U2552 : OAI22_X1 port map( A1 => n2903, A2 => n2971, B1 => n3647, B2 => 
                           n2972, ZN => n1875);
   U2553 : OAI22_X1 port map( A1 => n2904, A2 => n2971, B1 => n3646, B2 => 
                           n2972, ZN => n1874);
   U2554 : OAI22_X1 port map( A1 => n2905, A2 => n2971, B1 => n3645, B2 => 
                           n2972, ZN => n1873);
   U2555 : OAI22_X1 port map( A1 => n2906, A2 => n2971, B1 => n3644, B2 => 
                           n2972, ZN => n1872);
   U2556 : OAI22_X1 port map( A1 => n2907, A2 => n2971, B1 => n3643, B2 => 
                           n2972, ZN => n1871);
   U2557 : OAI22_X1 port map( A1 => n2908, A2 => n2971, B1 => n3642, B2 => 
                           n2972, ZN => n1870);
   U2558 : OAI22_X1 port map( A1 => n2909, A2 => n2971, B1 => n3641, B2 => 
                           n2972, ZN => n1869);
   U2559 : OAI22_X1 port map( A1 => n2910, A2 => n2971, B1 => n3640, B2 => 
                           n2972, ZN => n1868);
   U2560 : OAI22_X1 port map( A1 => n2911, A2 => n2971, B1 => n3639, B2 => 
                           n2972, ZN => n1867);
   U2561 : OAI22_X1 port map( A1 => n2912, A2 => n2971, B1 => n3638, B2 => 
                           n2972, ZN => n1866);
   U2562 : OAI22_X1 port map( A1 => n2913, A2 => n2971, B1 => n3637, B2 => 
                           n2972, ZN => n1865);
   U2563 : OAI22_X1 port map( A1 => n2914, A2 => n2971, B1 => n3636, B2 => 
                           n2972, ZN => n1864);
   U2564 : OAI22_X1 port map( A1 => n2915, A2 => n2971, B1 => n3635, B2 => 
                           n2972, ZN => n1863);
   U2565 : OAI22_X1 port map( A1 => n2916, A2 => n2971, B1 => n3634, B2 => 
                           n2972, ZN => n1862);
   U2566 : OAI22_X1 port map( A1 => n2917, A2 => n2971, B1 => n3633, B2 => 
                           n2972, ZN => n1861);
   U2567 : OAI22_X1 port map( A1 => n2918, A2 => n2971, B1 => n3632, B2 => 
                           n2972, ZN => n1860);
   U2568 : OAI22_X1 port map( A1 => n2919, A2 => n2971, B1 => n3631, B2 => 
                           n2972, ZN => n1859);
   U2569 : OAI22_X1 port map( A1 => n2920, A2 => n2971, B1 => n3630, B2 => 
                           n2972, ZN => n1858);
   U2570 : OAI22_X1 port map( A1 => n2921, A2 => n2971, B1 => n3629, B2 => 
                           n2972, ZN => n1857);
   U2571 : OAI22_X1 port map( A1 => n2922, A2 => n2971, B1 => n3628, B2 => 
                           n2972, ZN => n1856);
   U2572 : OAI22_X1 port map( A1 => n2923, A2 => n2971, B1 => n3627, B2 => 
                           n2972, ZN => n1855);
   U2573 : OAI22_X1 port map( A1 => n2924, A2 => n2971, B1 => n3626, B2 => 
                           n2972, ZN => n1854);
   U2574 : OAI22_X1 port map( A1 => n2925, A2 => n2971, B1 => n3625, B2 => 
                           n2972, ZN => n1853);
   U2575 : OAI22_X1 port map( A1 => n2926, A2 => n2971, B1 => n3624, B2 => 
                           n2972, ZN => n1852);
   U2576 : OAI22_X1 port map( A1 => n2927, A2 => n2971, B1 => n3623, B2 => 
                           n2972, ZN => n1851);
   U2577 : OAI22_X1 port map( A1 => n2928, A2 => n2971, B1 => n3622, B2 => 
                           n2972, ZN => n1850);
   U2578 : OAI22_X1 port map( A1 => n2929, A2 => n2971, B1 => n3621, B2 => 
                           n2972, ZN => n1849);
   U2579 : OAI22_X1 port map( A1 => n2930, A2 => n2971, B1 => n3620, B2 => 
                           n2972, ZN => n1848);
   U2580 : OAI22_X1 port map( A1 => n2931, A2 => n2971, B1 => n3619, B2 => 
                           n2972, ZN => n1847);
   U2581 : OAI22_X1 port map( A1 => n2899, A2 => n2973, B1 => n3618, B2 => 
                           n2974, ZN => n1846);
   U2582 : OAI22_X1 port map( A1 => n2901, A2 => n2973, B1 => n3617, B2 => 
                           n2974, ZN => n1845);
   U2583 : OAI22_X1 port map( A1 => n2902, A2 => n2973, B1 => n3616, B2 => 
                           n2974, ZN => n1844);
   U2584 : OAI22_X1 port map( A1 => n2903, A2 => n2973, B1 => n3615, B2 => 
                           n2974, ZN => n1843);
   U2585 : OAI22_X1 port map( A1 => n2904, A2 => n2973, B1 => n3614, B2 => 
                           n2974, ZN => n1842);
   U2586 : OAI22_X1 port map( A1 => n2905, A2 => n2973, B1 => n3613, B2 => 
                           n2974, ZN => n1841);
   U2587 : OAI22_X1 port map( A1 => n2906, A2 => n2973, B1 => n3612, B2 => 
                           n2974, ZN => n1840);
   U2588 : OAI22_X1 port map( A1 => n2907, A2 => n2973, B1 => n3611, B2 => 
                           n2974, ZN => n1839);
   U2589 : OAI22_X1 port map( A1 => n2908, A2 => n2973, B1 => n3610, B2 => 
                           n2974, ZN => n1838);
   U2590 : OAI22_X1 port map( A1 => n2909, A2 => n2973, B1 => n3609, B2 => 
                           n2974, ZN => n1837);
   U2591 : OAI22_X1 port map( A1 => n2910, A2 => n2973, B1 => n3608, B2 => 
                           n2974, ZN => n1836);
   U2592 : OAI22_X1 port map( A1 => n2911, A2 => n2973, B1 => n3607, B2 => 
                           n2974, ZN => n1835);
   U2593 : OAI22_X1 port map( A1 => n2912, A2 => n2973, B1 => n3606, B2 => 
                           n2974, ZN => n1834);
   U2594 : OAI22_X1 port map( A1 => n2913, A2 => n2973, B1 => n3605, B2 => 
                           n2974, ZN => n1833);
   U2595 : OAI22_X1 port map( A1 => n2914, A2 => n2973, B1 => n3604, B2 => 
                           n2974, ZN => n1832);
   U2596 : OAI22_X1 port map( A1 => n2915, A2 => n2973, B1 => n3603, B2 => 
                           n2974, ZN => n1831);
   U2597 : OAI22_X1 port map( A1 => n2916, A2 => n2973, B1 => n3602, B2 => 
                           n2974, ZN => n1830);
   U2598 : OAI22_X1 port map( A1 => n2917, A2 => n2973, B1 => n3601, B2 => 
                           n2974, ZN => n1829);
   U2599 : OAI22_X1 port map( A1 => n2918, A2 => n2973, B1 => n3600, B2 => 
                           n2974, ZN => n1828);
   U2600 : OAI22_X1 port map( A1 => n2919, A2 => n2973, B1 => n3599, B2 => 
                           n2974, ZN => n1827);
   U2601 : OAI22_X1 port map( A1 => n2920, A2 => n2973, B1 => n3598, B2 => 
                           n2974, ZN => n1826);
   U2602 : OAI22_X1 port map( A1 => n2921, A2 => n2973, B1 => n3597, B2 => 
                           n2974, ZN => n1825);
   U2603 : OAI22_X1 port map( A1 => n2922, A2 => n2973, B1 => n3596, B2 => 
                           n2974, ZN => n1824);
   U2604 : OAI22_X1 port map( A1 => n2923, A2 => n2973, B1 => n3595, B2 => 
                           n2974, ZN => n1823);
   U2605 : OAI22_X1 port map( A1 => n2924, A2 => n2973, B1 => n3594, B2 => 
                           n2974, ZN => n1822);
   U2606 : OAI22_X1 port map( A1 => n2925, A2 => n2973, B1 => n3593, B2 => 
                           n2974, ZN => n1821);
   U2607 : OAI22_X1 port map( A1 => n2926, A2 => n2973, B1 => n3592, B2 => 
                           n2974, ZN => n1820);
   U2608 : OAI22_X1 port map( A1 => n2927, A2 => n2973, B1 => n3591, B2 => 
                           n2974, ZN => n1819);
   U2609 : OAI22_X1 port map( A1 => n2928, A2 => n2973, B1 => n3590, B2 => 
                           n2974, ZN => n1818);
   U2610 : OAI22_X1 port map( A1 => n2929, A2 => n2973, B1 => n3589, B2 => 
                           n2974, ZN => n1817);
   U2611 : OAI22_X1 port map( A1 => n2930, A2 => n2973, B1 => n3588, B2 => 
                           n2974, ZN => n1816);
   U2612 : OAI22_X1 port map( A1 => n2931, A2 => n2973, B1 => n3587, B2 => 
                           n2974, ZN => n1815);
   U2613 : AND3_X1 port map( A1 => n2957, A2 => n2956, A3 => ADD_WR(3), ZN => 
                           n2960);
   U2614 : INV_X1 port map( A => ADD_WR(4), ZN => n2956);
   U2615 : OAI22_X1 port map( A1 => n2899, A2 => n2975, B1 => n3586, B2 => 
                           n2976, ZN => n1814);
   U2616 : OAI22_X1 port map( A1 => n2901, A2 => n2975, B1 => n3585, B2 => 
                           n2976, ZN => n1813);
   U2617 : OAI22_X1 port map( A1 => n2902, A2 => n2975, B1 => n3584, B2 => 
                           n2976, ZN => n1812);
   U2618 : OAI22_X1 port map( A1 => n2903, A2 => n2975, B1 => n3583, B2 => 
                           n2976, ZN => n1811);
   U2619 : OAI22_X1 port map( A1 => n2904, A2 => n2975, B1 => n3582, B2 => 
                           n2976, ZN => n1810);
   U2620 : OAI22_X1 port map( A1 => n2905, A2 => n2975, B1 => n3581, B2 => 
                           n2976, ZN => n1809);
   U2621 : OAI22_X1 port map( A1 => n2906, A2 => n2975, B1 => n3580, B2 => 
                           n2976, ZN => n1808);
   U2622 : OAI22_X1 port map( A1 => n2907, A2 => n2975, B1 => n3579, B2 => 
                           n2976, ZN => n1807);
   U2623 : OAI22_X1 port map( A1 => n2908, A2 => n2975, B1 => n3578, B2 => 
                           n2976, ZN => n1806);
   U2624 : OAI22_X1 port map( A1 => n2909, A2 => n2975, B1 => n3577, B2 => 
                           n2976, ZN => n1805);
   U2625 : OAI22_X1 port map( A1 => n2910, A2 => n2975, B1 => n3576, B2 => 
                           n2976, ZN => n1804);
   U2626 : OAI22_X1 port map( A1 => n2911, A2 => n2975, B1 => n3575, B2 => 
                           n2976, ZN => n1803);
   U2627 : OAI22_X1 port map( A1 => n2912, A2 => n2975, B1 => n3574, B2 => 
                           n2976, ZN => n1802);
   U2628 : OAI22_X1 port map( A1 => n2913, A2 => n2975, B1 => n3573, B2 => 
                           n2976, ZN => n1801);
   U2629 : OAI22_X1 port map( A1 => n2914, A2 => n2975, B1 => n3572, B2 => 
                           n2976, ZN => n1800);
   U2630 : OAI22_X1 port map( A1 => n2915, A2 => n2975, B1 => n3571, B2 => 
                           n2976, ZN => n1799);
   U2631 : OAI22_X1 port map( A1 => n2916, A2 => n2975, B1 => n3570, B2 => 
                           n2976, ZN => n1798);
   U2632 : OAI22_X1 port map( A1 => n2917, A2 => n2975, B1 => n3569, B2 => 
                           n2976, ZN => n1797);
   U2633 : OAI22_X1 port map( A1 => n2918, A2 => n2975, B1 => n3568, B2 => 
                           n2976, ZN => n1796);
   U2634 : OAI22_X1 port map( A1 => n2919, A2 => n2975, B1 => n3567, B2 => 
                           n2976, ZN => n1795);
   U2635 : OAI22_X1 port map( A1 => n2920, A2 => n2975, B1 => n3566, B2 => 
                           n2976, ZN => n1794);
   U2636 : OAI22_X1 port map( A1 => n2921, A2 => n2975, B1 => n3565, B2 => 
                           n2976, ZN => n1793);
   U2637 : OAI22_X1 port map( A1 => n2922, A2 => n2975, B1 => n3564, B2 => 
                           n2976, ZN => n1792);
   U2638 : OAI22_X1 port map( A1 => n2923, A2 => n2975, B1 => n3563, B2 => 
                           n2976, ZN => n1791);
   U2639 : OAI22_X1 port map( A1 => n2924, A2 => n2975, B1 => n3562, B2 => 
                           n2976, ZN => n1790);
   U2640 : OAI22_X1 port map( A1 => n2925, A2 => n2975, B1 => n3561, B2 => 
                           n2976, ZN => n1789);
   U2641 : OAI22_X1 port map( A1 => n2926, A2 => n2975, B1 => n3560, B2 => 
                           n2976, ZN => n1788);
   U2642 : OAI22_X1 port map( A1 => n2927, A2 => n2975, B1 => n3559, B2 => 
                           n2976, ZN => n1787);
   U2643 : OAI22_X1 port map( A1 => n2928, A2 => n2975, B1 => n3558, B2 => 
                           n2976, ZN => n1786);
   U2644 : OAI22_X1 port map( A1 => n2929, A2 => n2975, B1 => n3557, B2 => 
                           n2976, ZN => n1785);
   U2645 : OAI22_X1 port map( A1 => n2930, A2 => n2975, B1 => n3556, B2 => 
                           n2976, ZN => n1784);
   U2646 : OAI22_X1 port map( A1 => n2931, A2 => n2975, B1 => n3555, B2 => 
                           n2976, ZN => n1783);
   U2647 : OAI22_X1 port map( A1 => n2899, A2 => n2978, B1 => n3554, B2 => 
                           n2979, ZN => n1782);
   U2648 : OAI22_X1 port map( A1 => n2901, A2 => n2978, B1 => n3553, B2 => 
                           n2979, ZN => n1781);
   U2649 : OAI22_X1 port map( A1 => n2902, A2 => n2978, B1 => n3552, B2 => 
                           n2979, ZN => n1780);
   U2650 : OAI22_X1 port map( A1 => n2903, A2 => n2978, B1 => n3551, B2 => 
                           n2979, ZN => n1779);
   U2651 : OAI22_X1 port map( A1 => n2904, A2 => n2978, B1 => n3550, B2 => 
                           n2979, ZN => n1778);
   U2652 : OAI22_X1 port map( A1 => n2905, A2 => n2978, B1 => n3549, B2 => 
                           n2979, ZN => n1777);
   U2653 : OAI22_X1 port map( A1 => n2906, A2 => n2978, B1 => n3548, B2 => 
                           n2979, ZN => n1776);
   U2654 : OAI22_X1 port map( A1 => n2907, A2 => n2978, B1 => n3547, B2 => 
                           n2979, ZN => n1775);
   U2655 : OAI22_X1 port map( A1 => n2908, A2 => n2978, B1 => n3546, B2 => 
                           n2979, ZN => n1774);
   U2656 : OAI22_X1 port map( A1 => n2909, A2 => n2978, B1 => n3545, B2 => 
                           n2979, ZN => n1773);
   U2657 : OAI22_X1 port map( A1 => n2910, A2 => n2978, B1 => n3544, B2 => 
                           n2979, ZN => n1772);
   U2658 : OAI22_X1 port map( A1 => n2911, A2 => n2978, B1 => n3543, B2 => 
                           n2979, ZN => n1771);
   U2659 : OAI22_X1 port map( A1 => n2912, A2 => n2978, B1 => n3542, B2 => 
                           n2979, ZN => n1770);
   U2660 : OAI22_X1 port map( A1 => n2913, A2 => n2978, B1 => n3541, B2 => 
                           n2979, ZN => n1769);
   U2661 : OAI22_X1 port map( A1 => n2914, A2 => n2978, B1 => n3540, B2 => 
                           n2979, ZN => n1768);
   U2662 : OAI22_X1 port map( A1 => n2915, A2 => n2978, B1 => n3539, B2 => 
                           n2979, ZN => n1767);
   U2663 : OAI22_X1 port map( A1 => n2916, A2 => n2978, B1 => n3538, B2 => 
                           n2979, ZN => n1766);
   U2664 : OAI22_X1 port map( A1 => n2917, A2 => n2978, B1 => n3537, B2 => 
                           n2979, ZN => n1765);
   U2665 : OAI22_X1 port map( A1 => n2918, A2 => n2978, B1 => n3536, B2 => 
                           n2979, ZN => n1764);
   U2666 : OAI22_X1 port map( A1 => n2919, A2 => n2978, B1 => n3535, B2 => 
                           n2979, ZN => n1763);
   U2667 : OAI22_X1 port map( A1 => n2920, A2 => n2978, B1 => n3534, B2 => 
                           n2979, ZN => n1762);
   U2668 : OAI22_X1 port map( A1 => n2921, A2 => n2978, B1 => n3533, B2 => 
                           n2979, ZN => n1761);
   U2669 : OAI22_X1 port map( A1 => n2922, A2 => n2978, B1 => n3532, B2 => 
                           n2979, ZN => n1760);
   U2670 : OAI22_X1 port map( A1 => n2923, A2 => n2978, B1 => n3531, B2 => 
                           n2979, ZN => n1759);
   U2671 : OAI22_X1 port map( A1 => n2924, A2 => n2978, B1 => n3530, B2 => 
                           n2979, ZN => n1758);
   U2672 : OAI22_X1 port map( A1 => n2925, A2 => n2978, B1 => n3529, B2 => 
                           n2979, ZN => n1757);
   U2673 : OAI22_X1 port map( A1 => n2926, A2 => n2978, B1 => n3528, B2 => 
                           n2979, ZN => n1756);
   U2674 : OAI22_X1 port map( A1 => n2927, A2 => n2978, B1 => n3527, B2 => 
                           n2979, ZN => n1755);
   U2675 : OAI22_X1 port map( A1 => n2928, A2 => n2978, B1 => n3526, B2 => 
                           n2979, ZN => n1754);
   U2676 : OAI22_X1 port map( A1 => n2929, A2 => n2978, B1 => n3525, B2 => 
                           n2979, ZN => n1753);
   U2677 : OAI22_X1 port map( A1 => n2930, A2 => n2978, B1 => n3524, B2 => 
                           n2979, ZN => n1752);
   U2678 : OAI22_X1 port map( A1 => n2931, A2 => n2978, B1 => n3523, B2 => 
                           n2979, ZN => n1751);
   U2679 : OAI22_X1 port map( A1 => n2899, A2 => n2980, B1 => n3522, B2 => 
                           n2981, ZN => n1750);
   U2680 : OAI22_X1 port map( A1 => n2901, A2 => n2980, B1 => n3521, B2 => 
                           n2981, ZN => n1749);
   U2681 : OAI22_X1 port map( A1 => n2902, A2 => n2980, B1 => n3520, B2 => 
                           n2981, ZN => n1748);
   U2682 : OAI22_X1 port map( A1 => n2903, A2 => n2980, B1 => n3519, B2 => 
                           n2981, ZN => n1747);
   U2683 : OAI22_X1 port map( A1 => n2904, A2 => n2980, B1 => n3518, B2 => 
                           n2981, ZN => n1746);
   U2684 : OAI22_X1 port map( A1 => n2905, A2 => n2980, B1 => n3517, B2 => 
                           n2981, ZN => n1745);
   U2685 : OAI22_X1 port map( A1 => n2906, A2 => n2980, B1 => n3516, B2 => 
                           n2981, ZN => n1744);
   U2686 : OAI22_X1 port map( A1 => n2907, A2 => n2980, B1 => n3515, B2 => 
                           n2981, ZN => n1743);
   U2687 : OAI22_X1 port map( A1 => n2908, A2 => n2980, B1 => n3514, B2 => 
                           n2981, ZN => n1742);
   U2688 : OAI22_X1 port map( A1 => n2909, A2 => n2980, B1 => n3513, B2 => 
                           n2981, ZN => n1741);
   U2689 : OAI22_X1 port map( A1 => n2910, A2 => n2980, B1 => n3512, B2 => 
                           n2981, ZN => n1740);
   U2690 : OAI22_X1 port map( A1 => n2911, A2 => n2980, B1 => n3511, B2 => 
                           n2981, ZN => n1739);
   U2691 : OAI22_X1 port map( A1 => n2912, A2 => n2980, B1 => n3510, B2 => 
                           n2981, ZN => n1738);
   U2692 : OAI22_X1 port map( A1 => n2913, A2 => n2980, B1 => n3509, B2 => 
                           n2981, ZN => n1737);
   U2693 : OAI22_X1 port map( A1 => n2914, A2 => n2980, B1 => n3508, B2 => 
                           n2981, ZN => n1736);
   U2694 : OAI22_X1 port map( A1 => n2915, A2 => n2980, B1 => n3507, B2 => 
                           n2981, ZN => n1735);
   U2695 : OAI22_X1 port map( A1 => n2916, A2 => n2980, B1 => n3506, B2 => 
                           n2981, ZN => n1734);
   U2696 : OAI22_X1 port map( A1 => n2917, A2 => n2980, B1 => n3505, B2 => 
                           n2981, ZN => n1733);
   U2697 : OAI22_X1 port map( A1 => n2918, A2 => n2980, B1 => n3504, B2 => 
                           n2981, ZN => n1732);
   U2698 : OAI22_X1 port map( A1 => n2919, A2 => n2980, B1 => n3503, B2 => 
                           n2981, ZN => n1731);
   U2699 : OAI22_X1 port map( A1 => n2920, A2 => n2980, B1 => n3502, B2 => 
                           n2981, ZN => n1730);
   U2700 : OAI22_X1 port map( A1 => n2921, A2 => n2980, B1 => n3501, B2 => 
                           n2981, ZN => n1729);
   U2701 : OAI22_X1 port map( A1 => n2922, A2 => n2980, B1 => n3500, B2 => 
                           n2981, ZN => n1728);
   U2702 : OAI22_X1 port map( A1 => n2923, A2 => n2980, B1 => n3499, B2 => 
                           n2981, ZN => n1727);
   U2703 : OAI22_X1 port map( A1 => n2924, A2 => n2980, B1 => n3498, B2 => 
                           n2981, ZN => n1726);
   U2704 : OAI22_X1 port map( A1 => n2925, A2 => n2980, B1 => n3497, B2 => 
                           n2981, ZN => n1725);
   U2705 : OAI22_X1 port map( A1 => n2926, A2 => n2980, B1 => n3496, B2 => 
                           n2981, ZN => n1724);
   U2706 : OAI22_X1 port map( A1 => n2927, A2 => n2980, B1 => n3495, B2 => 
                           n2981, ZN => n1723);
   U2707 : OAI22_X1 port map( A1 => n2928, A2 => n2980, B1 => n3494, B2 => 
                           n2981, ZN => n1722);
   U2708 : OAI22_X1 port map( A1 => n2929, A2 => n2980, B1 => n3493, B2 => 
                           n2981, ZN => n1721);
   U2709 : OAI22_X1 port map( A1 => n2930, A2 => n2980, B1 => n3492, B2 => 
                           n2981, ZN => n1720);
   U2710 : OAI22_X1 port map( A1 => n2931, A2 => n2980, B1 => n3491, B2 => 
                           n2981, ZN => n1719);
   U2711 : OAI22_X1 port map( A1 => n2899, A2 => n2982, B1 => n3490, B2 => 
                           n2983, ZN => n1718);
   U2712 : OAI22_X1 port map( A1 => n2901, A2 => n2982, B1 => n3489, B2 => 
                           n2983, ZN => n1717);
   U2713 : OAI22_X1 port map( A1 => n2902, A2 => n2982, B1 => n3488, B2 => 
                           n2983, ZN => n1716);
   U2714 : OAI22_X1 port map( A1 => n2903, A2 => n2982, B1 => n3487, B2 => 
                           n2983, ZN => n1715);
   U2715 : OAI22_X1 port map( A1 => n2904, A2 => n2982, B1 => n3486, B2 => 
                           n2983, ZN => n1714);
   U2716 : OAI22_X1 port map( A1 => n2905, A2 => n2982, B1 => n3485, B2 => 
                           n2983, ZN => n1713);
   U2717 : OAI22_X1 port map( A1 => n2906, A2 => n2982, B1 => n3484, B2 => 
                           n2983, ZN => n1712);
   U2718 : OAI22_X1 port map( A1 => n2907, A2 => n2982, B1 => n3483, B2 => 
                           n2983, ZN => n1711);
   U2719 : OAI22_X1 port map( A1 => n2908, A2 => n2982, B1 => n3482, B2 => 
                           n2983, ZN => n1710);
   U2720 : OAI22_X1 port map( A1 => n2909, A2 => n2982, B1 => n3481, B2 => 
                           n2983, ZN => n1709);
   U2721 : OAI22_X1 port map( A1 => n2910, A2 => n2982, B1 => n3480, B2 => 
                           n2983, ZN => n1708);
   U2722 : OAI22_X1 port map( A1 => n2911, A2 => n2982, B1 => n3479, B2 => 
                           n2983, ZN => n1707);
   U2723 : OAI22_X1 port map( A1 => n2912, A2 => n2982, B1 => n3478, B2 => 
                           n2983, ZN => n1706);
   U2724 : OAI22_X1 port map( A1 => n2913, A2 => n2982, B1 => n3477, B2 => 
                           n2983, ZN => n1705);
   U2725 : OAI22_X1 port map( A1 => n2914, A2 => n2982, B1 => n3476, B2 => 
                           n2983, ZN => n1704);
   U2726 : OAI22_X1 port map( A1 => n2915, A2 => n2982, B1 => n3475, B2 => 
                           n2983, ZN => n1703);
   U2727 : OAI22_X1 port map( A1 => n2916, A2 => n2982, B1 => n3474, B2 => 
                           n2983, ZN => n1702);
   U2728 : OAI22_X1 port map( A1 => n2917, A2 => n2982, B1 => n3473, B2 => 
                           n2983, ZN => n1701);
   U2729 : OAI22_X1 port map( A1 => n2918, A2 => n2982, B1 => n3472, B2 => 
                           n2983, ZN => n1700);
   U2730 : OAI22_X1 port map( A1 => n2919, A2 => n2982, B1 => n3471, B2 => 
                           n2983, ZN => n1699);
   U2731 : OAI22_X1 port map( A1 => n2920, A2 => n2982, B1 => n3470, B2 => 
                           n2983, ZN => n1698);
   U2732 : OAI22_X1 port map( A1 => n2921, A2 => n2982, B1 => n3469, B2 => 
                           n2983, ZN => n1697);
   U2733 : OAI22_X1 port map( A1 => n2922, A2 => n2982, B1 => n3468, B2 => 
                           n2983, ZN => n1696);
   U2734 : OAI22_X1 port map( A1 => n2923, A2 => n2982, B1 => n3467, B2 => 
                           n2983, ZN => n1695);
   U2735 : OAI22_X1 port map( A1 => n2924, A2 => n2982, B1 => n3466, B2 => 
                           n2983, ZN => n1694);
   U2736 : OAI22_X1 port map( A1 => n2925, A2 => n2982, B1 => n3465, B2 => 
                           n2983, ZN => n1693);
   U2737 : OAI22_X1 port map( A1 => n2926, A2 => n2982, B1 => n3464, B2 => 
                           n2983, ZN => n1692);
   U2738 : OAI22_X1 port map( A1 => n2927, A2 => n2982, B1 => n3463, B2 => 
                           n2983, ZN => n1691);
   U2739 : OAI22_X1 port map( A1 => n2928, A2 => n2982, B1 => n3462, B2 => 
                           n2983, ZN => n1690);
   U2740 : OAI22_X1 port map( A1 => n2929, A2 => n2982, B1 => n3461, B2 => 
                           n2983, ZN => n1689);
   U2741 : OAI22_X1 port map( A1 => n2930, A2 => n2982, B1 => n3460, B2 => 
                           n2983, ZN => n1688);
   U2742 : OAI22_X1 port map( A1 => n2931, A2 => n2982, B1 => n3459, B2 => 
                           n2983, ZN => n1687);
   U2743 : OAI22_X1 port map( A1 => n2899, A2 => n2984, B1 => n3458, B2 => 
                           n2985, ZN => n1686);
   U2744 : OAI22_X1 port map( A1 => n2901, A2 => n2984, B1 => n3457, B2 => 
                           n2985, ZN => n1685);
   U2745 : OAI22_X1 port map( A1 => n2902, A2 => n2984, B1 => n3456, B2 => 
                           n2985, ZN => n1684);
   U2746 : OAI22_X1 port map( A1 => n2903, A2 => n2984, B1 => n3455, B2 => 
                           n2985, ZN => n1683);
   U2747 : OAI22_X1 port map( A1 => n2904, A2 => n2984, B1 => n3454, B2 => 
                           n2985, ZN => n1682);
   U2748 : OAI22_X1 port map( A1 => n2905, A2 => n2984, B1 => n3453, B2 => 
                           n2985, ZN => n1681);
   U2749 : OAI22_X1 port map( A1 => n2906, A2 => n2984, B1 => n3452, B2 => 
                           n2985, ZN => n1680);
   U2750 : OAI22_X1 port map( A1 => n2907, A2 => n2984, B1 => n3451, B2 => 
                           n2985, ZN => n1679);
   U2751 : OAI22_X1 port map( A1 => n2908, A2 => n2984, B1 => n3450, B2 => 
                           n2985, ZN => n1678);
   U2752 : OAI22_X1 port map( A1 => n2909, A2 => n2984, B1 => n3449, B2 => 
                           n2985, ZN => n1677);
   U2753 : OAI22_X1 port map( A1 => n2910, A2 => n2984, B1 => n3448, B2 => 
                           n2985, ZN => n1676);
   U2754 : OAI22_X1 port map( A1 => n2911, A2 => n2984, B1 => n3447, B2 => 
                           n2985, ZN => n1675);
   U2755 : OAI22_X1 port map( A1 => n2912, A2 => n2984, B1 => n3446, B2 => 
                           n2985, ZN => n1674);
   U2756 : OAI22_X1 port map( A1 => n2913, A2 => n2984, B1 => n3445, B2 => 
                           n2985, ZN => n1673);
   U2757 : OAI22_X1 port map( A1 => n2914, A2 => n2984, B1 => n3444, B2 => 
                           n2985, ZN => n1672);
   U2758 : OAI22_X1 port map( A1 => n2915, A2 => n2984, B1 => n3443, B2 => 
                           n2985, ZN => n1671);
   U2759 : OAI22_X1 port map( A1 => n2916, A2 => n2984, B1 => n3442, B2 => 
                           n2985, ZN => n1670);
   U2760 : OAI22_X1 port map( A1 => n2917, A2 => n2984, B1 => n3441, B2 => 
                           n2985, ZN => n1669);
   U2761 : OAI22_X1 port map( A1 => n2918, A2 => n2984, B1 => n3440, B2 => 
                           n2985, ZN => n1668);
   U2762 : OAI22_X1 port map( A1 => n2919, A2 => n2984, B1 => n3439, B2 => 
                           n2985, ZN => n1667);
   U2763 : OAI22_X1 port map( A1 => n2920, A2 => n2984, B1 => n3438, B2 => 
                           n2985, ZN => n1666);
   U2764 : OAI22_X1 port map( A1 => n2921, A2 => n2984, B1 => n3437, B2 => 
                           n2985, ZN => n1665);
   U2765 : OAI22_X1 port map( A1 => n2922, A2 => n2984, B1 => n3436, B2 => 
                           n2985, ZN => n1664);
   U2766 : OAI22_X1 port map( A1 => n2923, A2 => n2984, B1 => n3435, B2 => 
                           n2985, ZN => n1663);
   U2767 : OAI22_X1 port map( A1 => n2924, A2 => n2984, B1 => n3434, B2 => 
                           n2985, ZN => n1662);
   U2768 : OAI22_X1 port map( A1 => n2925, A2 => n2984, B1 => n3433, B2 => 
                           n2985, ZN => n1661);
   U2769 : OAI22_X1 port map( A1 => n2926, A2 => n2984, B1 => n3432, B2 => 
                           n2985, ZN => n1660);
   U2770 : OAI22_X1 port map( A1 => n2927, A2 => n2984, B1 => n3431, B2 => 
                           n2985, ZN => n1659);
   U2771 : OAI22_X1 port map( A1 => n2928, A2 => n2984, B1 => n3430, B2 => 
                           n2985, ZN => n1658);
   U2772 : OAI22_X1 port map( A1 => n2929, A2 => n2984, B1 => n3429, B2 => 
                           n2985, ZN => n1657);
   U2773 : OAI22_X1 port map( A1 => n2930, A2 => n2984, B1 => n3428, B2 => 
                           n2985, ZN => n1656);
   U2774 : OAI22_X1 port map( A1 => n2931, A2 => n2984, B1 => n3427, B2 => 
                           n2985, ZN => n1655);
   U2775 : OAI22_X1 port map( A1 => n2899, A2 => n2986, B1 => n3426, B2 => 
                           n2987, ZN => n1654);
   U2776 : OAI22_X1 port map( A1 => n2901, A2 => n2986, B1 => n3425, B2 => 
                           n2987, ZN => n1653);
   U2777 : OAI22_X1 port map( A1 => n2902, A2 => n2986, B1 => n3424, B2 => 
                           n2987, ZN => n1652);
   U2778 : OAI22_X1 port map( A1 => n2903, A2 => n2986, B1 => n3423, B2 => 
                           n2987, ZN => n1651);
   U2779 : OAI22_X1 port map( A1 => n2904, A2 => n2986, B1 => n3422, B2 => 
                           n2987, ZN => n1650);
   U2780 : OAI22_X1 port map( A1 => n2905, A2 => n2986, B1 => n3421, B2 => 
                           n2987, ZN => n1649);
   U2781 : OAI22_X1 port map( A1 => n2906, A2 => n2986, B1 => n3420, B2 => 
                           n2987, ZN => n1648);
   U2782 : OAI22_X1 port map( A1 => n2907, A2 => n2986, B1 => n3419, B2 => 
                           n2987, ZN => n1647);
   U2783 : OAI22_X1 port map( A1 => n2908, A2 => n2986, B1 => n3418, B2 => 
                           n2987, ZN => n1646);
   U2784 : OAI22_X1 port map( A1 => n2909, A2 => n2986, B1 => n3417, B2 => 
                           n2987, ZN => n1645);
   U2785 : OAI22_X1 port map( A1 => n2910, A2 => n2986, B1 => n3416, B2 => 
                           n2987, ZN => n1644);
   U2786 : OAI22_X1 port map( A1 => n2911, A2 => n2986, B1 => n3415, B2 => 
                           n2987, ZN => n1643);
   U2787 : OAI22_X1 port map( A1 => n2912, A2 => n2986, B1 => n3414, B2 => 
                           n2987, ZN => n1642);
   U2788 : OAI22_X1 port map( A1 => n2913, A2 => n2986, B1 => n3413, B2 => 
                           n2987, ZN => n1641);
   U2789 : OAI22_X1 port map( A1 => n2914, A2 => n2986, B1 => n3412, B2 => 
                           n2987, ZN => n1640);
   U2790 : OAI22_X1 port map( A1 => n2915, A2 => n2986, B1 => n3411, B2 => 
                           n2987, ZN => n1639);
   U2791 : OAI22_X1 port map( A1 => n2916, A2 => n2986, B1 => n3410, B2 => 
                           n2987, ZN => n1638);
   U2792 : OAI22_X1 port map( A1 => n2917, A2 => n2986, B1 => n3409, B2 => 
                           n2987, ZN => n1637);
   U2793 : OAI22_X1 port map( A1 => n2918, A2 => n2986, B1 => n3408, B2 => 
                           n2987, ZN => n1636);
   U2794 : OAI22_X1 port map( A1 => n2919, A2 => n2986, B1 => n3407, B2 => 
                           n2987, ZN => n1635);
   U2795 : OAI22_X1 port map( A1 => n2920, A2 => n2986, B1 => n3406, B2 => 
                           n2987, ZN => n1634);
   U2796 : OAI22_X1 port map( A1 => n2921, A2 => n2986, B1 => n3405, B2 => 
                           n2987, ZN => n1633);
   U2797 : OAI22_X1 port map( A1 => n2922, A2 => n2986, B1 => n3404, B2 => 
                           n2987, ZN => n1632);
   U2798 : OAI22_X1 port map( A1 => n2923, A2 => n2986, B1 => n3403, B2 => 
                           n2987, ZN => n1631);
   U2799 : OAI22_X1 port map( A1 => n2924, A2 => n2986, B1 => n3402, B2 => 
                           n2987, ZN => n1630);
   U2800 : OAI22_X1 port map( A1 => n2925, A2 => n2986, B1 => n3401, B2 => 
                           n2987, ZN => n1629);
   U2801 : OAI22_X1 port map( A1 => n2926, A2 => n2986, B1 => n3400, B2 => 
                           n2987, ZN => n1628);
   U2802 : OAI22_X1 port map( A1 => n2927, A2 => n2986, B1 => n3399, B2 => 
                           n2987, ZN => n1627);
   U2803 : OAI22_X1 port map( A1 => n2928, A2 => n2986, B1 => n3398, B2 => 
                           n2987, ZN => n1626);
   U2804 : OAI22_X1 port map( A1 => n2929, A2 => n2986, B1 => n3397, B2 => 
                           n2987, ZN => n1625);
   U2805 : OAI22_X1 port map( A1 => n2930, A2 => n2986, B1 => n3396, B2 => 
                           n2987, ZN => n1624);
   U2806 : OAI22_X1 port map( A1 => n2931, A2 => n2986, B1 => n3395, B2 => 
                           n2987, ZN => n1623);
   U2807 : OAI22_X1 port map( A1 => n2899, A2 => n2988, B1 => n3394, B2 => 
                           n2989, ZN => n1622);
   U2808 : OAI22_X1 port map( A1 => n2901, A2 => n2988, B1 => n3393, B2 => 
                           n2989, ZN => n1621);
   U2809 : OAI22_X1 port map( A1 => n2902, A2 => n2988, B1 => n3392, B2 => 
                           n2989, ZN => n1620);
   U2810 : OAI22_X1 port map( A1 => n2903, A2 => n2988, B1 => n3391, B2 => 
                           n2989, ZN => n1619);
   U2811 : OAI22_X1 port map( A1 => n2904, A2 => n2988, B1 => n3390, B2 => 
                           n2989, ZN => n1618);
   U2812 : OAI22_X1 port map( A1 => n2905, A2 => n2988, B1 => n3389, B2 => 
                           n2989, ZN => n1617);
   U2813 : OAI22_X1 port map( A1 => n2906, A2 => n2988, B1 => n3388, B2 => 
                           n2989, ZN => n1616);
   U2814 : OAI22_X1 port map( A1 => n2907, A2 => n2988, B1 => n3387, B2 => 
                           n2989, ZN => n1615);
   U2815 : OAI22_X1 port map( A1 => n2908, A2 => n2988, B1 => n3386, B2 => 
                           n2989, ZN => n1614);
   U2816 : OAI22_X1 port map( A1 => n2909, A2 => n2988, B1 => n3385, B2 => 
                           n2989, ZN => n1613);
   U2817 : OAI22_X1 port map( A1 => n2910, A2 => n2988, B1 => n3384, B2 => 
                           n2989, ZN => n1612);
   U2818 : OAI22_X1 port map( A1 => n2911, A2 => n2988, B1 => n3383, B2 => 
                           n2989, ZN => n1611);
   U2819 : OAI22_X1 port map( A1 => n2912, A2 => n2988, B1 => n3382, B2 => 
                           n2989, ZN => n1610);
   U2820 : OAI22_X1 port map( A1 => n2913, A2 => n2988, B1 => n3381, B2 => 
                           n2989, ZN => n1609);
   U2821 : OAI22_X1 port map( A1 => n2914, A2 => n2988, B1 => n3380, B2 => 
                           n2989, ZN => n1608);
   U2822 : OAI22_X1 port map( A1 => n2915, A2 => n2988, B1 => n3379, B2 => 
                           n2989, ZN => n1607);
   U2823 : OAI22_X1 port map( A1 => n2916, A2 => n2988, B1 => n3378, B2 => 
                           n2989, ZN => n1606);
   U2824 : OAI22_X1 port map( A1 => n2917, A2 => n2988, B1 => n3377, B2 => 
                           n2989, ZN => n1605);
   U2825 : OAI22_X1 port map( A1 => n2918, A2 => n2988, B1 => n3376, B2 => 
                           n2989, ZN => n1604);
   U2826 : OAI22_X1 port map( A1 => n2919, A2 => n2988, B1 => n3375, B2 => 
                           n2989, ZN => n1603);
   U2827 : OAI22_X1 port map( A1 => n2920, A2 => n2988, B1 => n3374, B2 => 
                           n2989, ZN => n1602);
   U2828 : OAI22_X1 port map( A1 => n2921, A2 => n2988, B1 => n3373, B2 => 
                           n2989, ZN => n1601);
   U2829 : OAI22_X1 port map( A1 => n2922, A2 => n2988, B1 => n3372, B2 => 
                           n2989, ZN => n1600);
   U2830 : OAI22_X1 port map( A1 => n2923, A2 => n2988, B1 => n3371, B2 => 
                           n2989, ZN => n1599);
   U2831 : OAI22_X1 port map( A1 => n2924, A2 => n2988, B1 => n3370, B2 => 
                           n2989, ZN => n1598);
   U2832 : OAI22_X1 port map( A1 => n2925, A2 => n2988, B1 => n3369, B2 => 
                           n2989, ZN => n1597);
   U2833 : OAI22_X1 port map( A1 => n2926, A2 => n2988, B1 => n3368, B2 => 
                           n2989, ZN => n1596);
   U2834 : OAI22_X1 port map( A1 => n2927, A2 => n2988, B1 => n3367, B2 => 
                           n2989, ZN => n1595);
   U2835 : OAI22_X1 port map( A1 => n2928, A2 => n2988, B1 => n3366, B2 => 
                           n2989, ZN => n1594);
   U2836 : OAI22_X1 port map( A1 => n2929, A2 => n2988, B1 => n3365, B2 => 
                           n2989, ZN => n1593);
   U2837 : OAI22_X1 port map( A1 => n2930, A2 => n2988, B1 => n3364, B2 => 
                           n2989, ZN => n1592);
   U2838 : OAI22_X1 port map( A1 => n2931, A2 => n2988, B1 => n3363, B2 => 
                           n2989, ZN => n1591);
   U2839 : OAI22_X1 port map( A1 => n2899, A2 => n2990, B1 => n3362, B2 => 
                           n2991, ZN => n1590);
   U2840 : OAI22_X1 port map( A1 => n2901, A2 => n2990, B1 => n3361, B2 => 
                           n2991, ZN => n1589);
   U2841 : OAI22_X1 port map( A1 => n2902, A2 => n2990, B1 => n3360, B2 => 
                           n2991, ZN => n1588);
   U2842 : OAI22_X1 port map( A1 => n2903, A2 => n2990, B1 => n3359, B2 => 
                           n2991, ZN => n1587);
   U2843 : OAI22_X1 port map( A1 => n2904, A2 => n2990, B1 => n3358, B2 => 
                           n2991, ZN => n1586);
   U2844 : OAI22_X1 port map( A1 => n2905, A2 => n2990, B1 => n3357, B2 => 
                           n2991, ZN => n1585);
   U2845 : OAI22_X1 port map( A1 => n2906, A2 => n2990, B1 => n3356, B2 => 
                           n2991, ZN => n1584);
   U2846 : OAI22_X1 port map( A1 => n2907, A2 => n2990, B1 => n3355, B2 => 
                           n2991, ZN => n1583);
   U2847 : OAI22_X1 port map( A1 => n2908, A2 => n2990, B1 => n3354, B2 => 
                           n2991, ZN => n1582);
   U2848 : OAI22_X1 port map( A1 => n2909, A2 => n2990, B1 => n3353, B2 => 
                           n2991, ZN => n1581);
   U2849 : OAI22_X1 port map( A1 => n2910, A2 => n2990, B1 => n3352, B2 => 
                           n2991, ZN => n1580);
   U2850 : OAI22_X1 port map( A1 => n2911, A2 => n2990, B1 => n3351, B2 => 
                           n2991, ZN => n1579);
   U2851 : OAI22_X1 port map( A1 => n2912, A2 => n2990, B1 => n3350, B2 => 
                           n2991, ZN => n1578);
   U2852 : OAI22_X1 port map( A1 => n2913, A2 => n2990, B1 => n3349, B2 => 
                           n2991, ZN => n1577);
   U2853 : OAI22_X1 port map( A1 => n2914, A2 => n2990, B1 => n3348, B2 => 
                           n2991, ZN => n1576);
   U2854 : OAI22_X1 port map( A1 => n2915, A2 => n2990, B1 => n3347, B2 => 
                           n2991, ZN => n1575);
   U2855 : OAI22_X1 port map( A1 => n2916, A2 => n2990, B1 => n3346, B2 => 
                           n2991, ZN => n1574);
   U2856 : OAI22_X1 port map( A1 => n2917, A2 => n2990, B1 => n3345, B2 => 
                           n2991, ZN => n1573);
   U2857 : OAI22_X1 port map( A1 => n2918, A2 => n2990, B1 => n3344, B2 => 
                           n2991, ZN => n1572);
   U2858 : OAI22_X1 port map( A1 => n2919, A2 => n2990, B1 => n3343, B2 => 
                           n2991, ZN => n1571);
   U2859 : OAI22_X1 port map( A1 => n2920, A2 => n2990, B1 => n3342, B2 => 
                           n2991, ZN => n1570);
   U2860 : OAI22_X1 port map( A1 => n2921, A2 => n2990, B1 => n3341, B2 => 
                           n2991, ZN => n1569);
   U2861 : OAI22_X1 port map( A1 => n2922, A2 => n2990, B1 => n3340, B2 => 
                           n2991, ZN => n1568);
   U2862 : OAI22_X1 port map( A1 => n2923, A2 => n2990, B1 => n3339, B2 => 
                           n2991, ZN => n1567);
   U2863 : OAI22_X1 port map( A1 => n2924, A2 => n2990, B1 => n3338, B2 => 
                           n2991, ZN => n1566);
   U2864 : OAI22_X1 port map( A1 => n2925, A2 => n2990, B1 => n3337, B2 => 
                           n2991, ZN => n1565);
   U2865 : OAI22_X1 port map( A1 => n2926, A2 => n2990, B1 => n3336, B2 => 
                           n2991, ZN => n1564);
   U2866 : OAI22_X1 port map( A1 => n2927, A2 => n2990, B1 => n3335, B2 => 
                           n2991, ZN => n1563);
   U2867 : OAI22_X1 port map( A1 => n2928, A2 => n2990, B1 => n3334, B2 => 
                           n2991, ZN => n1562);
   U2868 : OAI22_X1 port map( A1 => n2929, A2 => n2990, B1 => n3333, B2 => 
                           n2991, ZN => n1561);
   U2869 : OAI22_X1 port map( A1 => n2930, A2 => n2990, B1 => n3332, B2 => 
                           n2991, ZN => n1560);
   U2870 : OAI22_X1 port map( A1 => n2931, A2 => n2990, B1 => n3331, B2 => 
                           n2991, ZN => n1559);
   U2871 : AND3_X1 port map( A1 => n2957, A2 => n2955, A3 => ADD_WR(4), ZN => 
                           n2977);
   U2872 : INV_X1 port map( A => ADD_WR(3), ZN => n2955);
   U2873 : OAI22_X1 port map( A1 => n2899, A2 => n2992, B1 => n3330, B2 => 
                           n2993, ZN => n1558);
   U2874 : OAI22_X1 port map( A1 => n2901, A2 => n2992, B1 => n3329, B2 => 
                           n2993, ZN => n1557);
   U2875 : OAI22_X1 port map( A1 => n2902, A2 => n2992, B1 => n3328, B2 => 
                           n2993, ZN => n1556);
   U2876 : OAI22_X1 port map( A1 => n2903, A2 => n2992, B1 => n3327, B2 => 
                           n2993, ZN => n1555);
   U2877 : OAI22_X1 port map( A1 => n2904, A2 => n2992, B1 => n3326, B2 => 
                           n2993, ZN => n1554);
   U2878 : OAI22_X1 port map( A1 => n2905, A2 => n2992, B1 => n3325, B2 => 
                           n2993, ZN => n1553);
   U2879 : OAI22_X1 port map( A1 => n2906, A2 => n2992, B1 => n3324, B2 => 
                           n2993, ZN => n1552);
   U2880 : OAI22_X1 port map( A1 => n2907, A2 => n2992, B1 => n3323, B2 => 
                           n2993, ZN => n1551);
   U2881 : OAI22_X1 port map( A1 => n2908, A2 => n2992, B1 => n3322, B2 => 
                           n2993, ZN => n1550);
   U2882 : OAI22_X1 port map( A1 => n2909, A2 => n2992, B1 => n3321, B2 => 
                           n2993, ZN => n1549);
   U2883 : OAI22_X1 port map( A1 => n2910, A2 => n2992, B1 => n3320, B2 => 
                           n2993, ZN => n1548);
   U2884 : OAI22_X1 port map( A1 => n2911, A2 => n2992, B1 => n3319, B2 => 
                           n2993, ZN => n1547);
   U2885 : OAI22_X1 port map( A1 => n2912, A2 => n2992, B1 => n3318, B2 => 
                           n2993, ZN => n1546);
   U2886 : OAI22_X1 port map( A1 => n2913, A2 => n2992, B1 => n3317, B2 => 
                           n2993, ZN => n1545);
   U2887 : OAI22_X1 port map( A1 => n2914, A2 => n2992, B1 => n3316, B2 => 
                           n2993, ZN => n1544);
   U2888 : OAI22_X1 port map( A1 => n2915, A2 => n2992, B1 => n3315, B2 => 
                           n2993, ZN => n1543);
   U2889 : OAI22_X1 port map( A1 => n2916, A2 => n2992, B1 => n3314, B2 => 
                           n2993, ZN => n1542);
   U2890 : OAI22_X1 port map( A1 => n2917, A2 => n2992, B1 => n3313, B2 => 
                           n2993, ZN => n1541);
   U2891 : OAI22_X1 port map( A1 => n2918, A2 => n2992, B1 => n3312, B2 => 
                           n2993, ZN => n1540);
   U2892 : OAI22_X1 port map( A1 => n2919, A2 => n2992, B1 => n3311, B2 => 
                           n2993, ZN => n1539);
   U2893 : OAI22_X1 port map( A1 => n2920, A2 => n2992, B1 => n3310, B2 => 
                           n2993, ZN => n1538);
   U2894 : OAI22_X1 port map( A1 => n2921, A2 => n2992, B1 => n3309, B2 => 
                           n2993, ZN => n1537);
   U2895 : OAI22_X1 port map( A1 => n2922, A2 => n2992, B1 => n3308, B2 => 
                           n2993, ZN => n1536);
   U2896 : OAI22_X1 port map( A1 => n2923, A2 => n2992, B1 => n3307, B2 => 
                           n2993, ZN => n1535);
   U2897 : OAI22_X1 port map( A1 => n2924, A2 => n2992, B1 => n3306, B2 => 
                           n2993, ZN => n1534);
   U2898 : OAI22_X1 port map( A1 => n2925, A2 => n2992, B1 => n3305, B2 => 
                           n2993, ZN => n1533);
   U2899 : OAI22_X1 port map( A1 => n2926, A2 => n2992, B1 => n3304, B2 => 
                           n2993, ZN => n1532);
   U2900 : OAI22_X1 port map( A1 => n2927, A2 => n2992, B1 => n3303, B2 => 
                           n2993, ZN => n1531);
   U2901 : OAI22_X1 port map( A1 => n2928, A2 => n2992, B1 => n3302, B2 => 
                           n2993, ZN => n1530);
   U2902 : OAI22_X1 port map( A1 => n2929, A2 => n2992, B1 => n3301, B2 => 
                           n2993, ZN => n1529);
   U2903 : OAI22_X1 port map( A1 => n2930, A2 => n2992, B1 => n3300, B2 => 
                           n2993, ZN => n1528);
   U2904 : OAI22_X1 port map( A1 => n2931, A2 => n2992, B1 => n3299, B2 => 
                           n2993, ZN => n1527);
   U2905 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => ADD_WR(0),
                           ZN => n2932);
   U2906 : OAI22_X1 port map( A1 => n2899, A2 => n2995, B1 => n3298, B2 => 
                           n2996, ZN => n1526);
   U2907 : OAI22_X1 port map( A1 => n2901, A2 => n2995, B1 => n3297, B2 => 
                           n2996, ZN => n1525);
   U2908 : OAI22_X1 port map( A1 => n2902, A2 => n2995, B1 => n3296, B2 => 
                           n2996, ZN => n1524);
   U2909 : OAI22_X1 port map( A1 => n2903, A2 => n2995, B1 => n3295, B2 => 
                           n2996, ZN => n1523);
   U2910 : OAI22_X1 port map( A1 => n2904, A2 => n2995, B1 => n3294, B2 => 
                           n2996, ZN => n1522);
   U2911 : OAI22_X1 port map( A1 => n2905, A2 => n2995, B1 => n3293, B2 => 
                           n2996, ZN => n1521);
   U2912 : OAI22_X1 port map( A1 => n2906, A2 => n2995, B1 => n3292, B2 => 
                           n2996, ZN => n1520);
   U2913 : OAI22_X1 port map( A1 => n2907, A2 => n2995, B1 => n3291, B2 => 
                           n2996, ZN => n1519);
   U2914 : OAI22_X1 port map( A1 => n2908, A2 => n2995, B1 => n3290, B2 => 
                           n2996, ZN => n1518);
   U2915 : OAI22_X1 port map( A1 => n2909, A2 => n2995, B1 => n3289, B2 => 
                           n2996, ZN => n1517);
   U2916 : OAI22_X1 port map( A1 => n2910, A2 => n2995, B1 => n3288, B2 => 
                           n2996, ZN => n1516);
   U2917 : OAI22_X1 port map( A1 => n2911, A2 => n2995, B1 => n3287, B2 => 
                           n2996, ZN => n1515);
   U2918 : OAI22_X1 port map( A1 => n2912, A2 => n2995, B1 => n3286, B2 => 
                           n2996, ZN => n1514);
   U2919 : OAI22_X1 port map( A1 => n2913, A2 => n2995, B1 => n3285, B2 => 
                           n2996, ZN => n1513);
   U2920 : OAI22_X1 port map( A1 => n2914, A2 => n2995, B1 => n3284, B2 => 
                           n2996, ZN => n1512);
   U2921 : OAI22_X1 port map( A1 => n2915, A2 => n2995, B1 => n3283, B2 => 
                           n2996, ZN => n1511);
   U2922 : OAI22_X1 port map( A1 => n2916, A2 => n2995, B1 => n3282, B2 => 
                           n2996, ZN => n1510);
   U2923 : OAI22_X1 port map( A1 => n2917, A2 => n2995, B1 => n3281, B2 => 
                           n2996, ZN => n1509);
   U2924 : OAI22_X1 port map( A1 => n2918, A2 => n2995, B1 => n3280, B2 => 
                           n2996, ZN => n1508);
   U2925 : OAI22_X1 port map( A1 => n2919, A2 => n2995, B1 => n3279, B2 => 
                           n2996, ZN => n1507);
   U2926 : OAI22_X1 port map( A1 => n2920, A2 => n2995, B1 => n3278, B2 => 
                           n2996, ZN => n1506);
   U2927 : OAI22_X1 port map( A1 => n2921, A2 => n2995, B1 => n3277, B2 => 
                           n2996, ZN => n1505);
   U2928 : OAI22_X1 port map( A1 => n2922, A2 => n2995, B1 => n3276, B2 => 
                           n2996, ZN => n1504);
   U2929 : OAI22_X1 port map( A1 => n2923, A2 => n2995, B1 => n3275, B2 => 
                           n2996, ZN => n1503);
   U2930 : OAI22_X1 port map( A1 => n2924, A2 => n2995, B1 => n3274, B2 => 
                           n2996, ZN => n1502);
   U2931 : OAI22_X1 port map( A1 => n2925, A2 => n2995, B1 => n3273, B2 => 
                           n2996, ZN => n1501);
   U2932 : OAI22_X1 port map( A1 => n2926, A2 => n2995, B1 => n3272, B2 => 
                           n2996, ZN => n1500);
   U2933 : OAI22_X1 port map( A1 => n2927, A2 => n2995, B1 => n3271, B2 => 
                           n2996, ZN => n1499);
   U2934 : OAI22_X1 port map( A1 => n2928, A2 => n2995, B1 => n3270, B2 => 
                           n2996, ZN => n1498);
   U2935 : OAI22_X1 port map( A1 => n2929, A2 => n2995, B1 => n3269, B2 => 
                           n2996, ZN => n1497);
   U2936 : OAI22_X1 port map( A1 => n2930, A2 => n2995, B1 => n3268, B2 => 
                           n2996, ZN => n1496);
   U2937 : OAI22_X1 port map( A1 => n2931, A2 => n2995, B1 => n3267, B2 => 
                           n2996, ZN => n1495);
   U2938 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n2997, ZN 
                           => n2936);
   U2939 : OAI22_X1 port map( A1 => n2899, A2 => n2998, B1 => n3266, B2 => 
                           n2999, ZN => n1494);
   U2940 : OAI22_X1 port map( A1 => n2901, A2 => n2998, B1 => n3265, B2 => 
                           n2999, ZN => n1493);
   U2941 : OAI22_X1 port map( A1 => n2902, A2 => n2998, B1 => n3264, B2 => 
                           n2999, ZN => n1492);
   U2942 : OAI22_X1 port map( A1 => n2903, A2 => n2998, B1 => n3263, B2 => 
                           n2999, ZN => n1491);
   U2943 : OAI22_X1 port map( A1 => n2904, A2 => n2998, B1 => n3262, B2 => 
                           n2999, ZN => n1490);
   U2944 : OAI22_X1 port map( A1 => n2905, A2 => n2998, B1 => n3261, B2 => 
                           n2999, ZN => n1489);
   U2945 : OAI22_X1 port map( A1 => n2906, A2 => n2998, B1 => n3260, B2 => 
                           n2999, ZN => n1488);
   U2946 : OAI22_X1 port map( A1 => n2907, A2 => n2998, B1 => n3259, B2 => 
                           n2999, ZN => n1487);
   U2947 : OAI22_X1 port map( A1 => n2908, A2 => n2998, B1 => n3258, B2 => 
                           n2999, ZN => n1486);
   U2948 : OAI22_X1 port map( A1 => n2909, A2 => n2998, B1 => n3257, B2 => 
                           n2999, ZN => n1485);
   U2949 : OAI22_X1 port map( A1 => n2910, A2 => n2998, B1 => n3256, B2 => 
                           n2999, ZN => n1484);
   U2950 : OAI22_X1 port map( A1 => n2911, A2 => n2998, B1 => n3255, B2 => 
                           n2999, ZN => n1483);
   U2951 : OAI22_X1 port map( A1 => n2912, A2 => n2998, B1 => n3254, B2 => 
                           n2999, ZN => n1482);
   U2952 : OAI22_X1 port map( A1 => n2913, A2 => n2998, B1 => n3253, B2 => 
                           n2999, ZN => n1481);
   U2953 : OAI22_X1 port map( A1 => n2914, A2 => n2998, B1 => n3252, B2 => 
                           n2999, ZN => n1480);
   U2954 : OAI22_X1 port map( A1 => n2915, A2 => n2998, B1 => n3251, B2 => 
                           n2999, ZN => n1479);
   U2955 : OAI22_X1 port map( A1 => n2916, A2 => n2998, B1 => n3250, B2 => 
                           n2999, ZN => n1478);
   U2956 : OAI22_X1 port map( A1 => n2917, A2 => n2998, B1 => n3249, B2 => 
                           n2999, ZN => n1477);
   U2957 : OAI22_X1 port map( A1 => n2918, A2 => n2998, B1 => n3248, B2 => 
                           n2999, ZN => n1476);
   U2958 : OAI22_X1 port map( A1 => n2919, A2 => n2998, B1 => n3247, B2 => 
                           n2999, ZN => n1475);
   U2959 : OAI22_X1 port map( A1 => n2920, A2 => n2998, B1 => n3246, B2 => 
                           n2999, ZN => n1474);
   U2960 : OAI22_X1 port map( A1 => n2921, A2 => n2998, B1 => n3245, B2 => 
                           n2999, ZN => n1473);
   U2961 : OAI22_X1 port map( A1 => n2922, A2 => n2998, B1 => n3244, B2 => 
                           n2999, ZN => n1472);
   U2962 : OAI22_X1 port map( A1 => n2923, A2 => n2998, B1 => n3243, B2 => 
                           n2999, ZN => n1471);
   U2963 : OAI22_X1 port map( A1 => n2924, A2 => n2998, B1 => n3242, B2 => 
                           n2999, ZN => n1470);
   U2964 : OAI22_X1 port map( A1 => n2925, A2 => n2998, B1 => n3241, B2 => 
                           n2999, ZN => n1469);
   U2965 : OAI22_X1 port map( A1 => n2926, A2 => n2998, B1 => n3240, B2 => 
                           n2999, ZN => n1468);
   U2966 : OAI22_X1 port map( A1 => n2927, A2 => n2998, B1 => n3239, B2 => 
                           n2999, ZN => n1467);
   U2967 : OAI22_X1 port map( A1 => n2928, A2 => n2998, B1 => n3238, B2 => 
                           n2999, ZN => n1466);
   U2968 : OAI22_X1 port map( A1 => n2929, A2 => n2998, B1 => n3237, B2 => 
                           n2999, ZN => n1465);
   U2969 : OAI22_X1 port map( A1 => n2930, A2 => n2998, B1 => n3236, B2 => 
                           n2999, ZN => n1464);
   U2970 : OAI22_X1 port map( A1 => n2931, A2 => n2998, B1 => n3235, B2 => 
                           n2999, ZN => n1463);
   U2971 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n3000, ZN 
                           => n2939);
   U2972 : OAI22_X1 port map( A1 => n2899, A2 => n3001, B1 => n3234, B2 => 
                           n3002, ZN => n1462);
   U2973 : OAI22_X1 port map( A1 => n2901, A2 => n3001, B1 => n3233, B2 => 
                           n3002, ZN => n1461);
   U2974 : OAI22_X1 port map( A1 => n2902, A2 => n3001, B1 => n3232, B2 => 
                           n3002, ZN => n1460);
   U2975 : OAI22_X1 port map( A1 => n2903, A2 => n3001, B1 => n3231, B2 => 
                           n3002, ZN => n1459);
   U2976 : OAI22_X1 port map( A1 => n2904, A2 => n3001, B1 => n3230, B2 => 
                           n3002, ZN => n1458);
   U2977 : OAI22_X1 port map( A1 => n2905, A2 => n3001, B1 => n3229, B2 => 
                           n3002, ZN => n1457);
   U2978 : OAI22_X1 port map( A1 => n2906, A2 => n3001, B1 => n3228, B2 => 
                           n3002, ZN => n1456);
   U2979 : OAI22_X1 port map( A1 => n2907, A2 => n3001, B1 => n3227, B2 => 
                           n3002, ZN => n1455);
   U2980 : OAI22_X1 port map( A1 => n2908, A2 => n3001, B1 => n3226, B2 => 
                           n3002, ZN => n1454);
   U2981 : OAI22_X1 port map( A1 => n2909, A2 => n3001, B1 => n3225, B2 => 
                           n3002, ZN => n1453);
   U2982 : OAI22_X1 port map( A1 => n2910, A2 => n3001, B1 => n3224, B2 => 
                           n3002, ZN => n1452);
   U2983 : OAI22_X1 port map( A1 => n2911, A2 => n3001, B1 => n3223, B2 => 
                           n3002, ZN => n1451);
   U2984 : OAI22_X1 port map( A1 => n2912, A2 => n3001, B1 => n3222, B2 => 
                           n3002, ZN => n1450);
   U2985 : OAI22_X1 port map( A1 => n2913, A2 => n3001, B1 => n3221, B2 => 
                           n3002, ZN => n1449);
   U2986 : OAI22_X1 port map( A1 => n2914, A2 => n3001, B1 => n3220, B2 => 
                           n3002, ZN => n1448);
   U2987 : OAI22_X1 port map( A1 => n2915, A2 => n3001, B1 => n3219, B2 => 
                           n3002, ZN => n1447);
   U2988 : OAI22_X1 port map( A1 => n2916, A2 => n3001, B1 => n3218, B2 => 
                           n3002, ZN => n1446);
   U2989 : OAI22_X1 port map( A1 => n2917, A2 => n3001, B1 => n3217, B2 => 
                           n3002, ZN => n1445);
   U2990 : OAI22_X1 port map( A1 => n2918, A2 => n3001, B1 => n3216, B2 => 
                           n3002, ZN => n1444);
   U2991 : OAI22_X1 port map( A1 => n2919, A2 => n3001, B1 => n3215, B2 => 
                           n3002, ZN => n1443);
   U2992 : OAI22_X1 port map( A1 => n2920, A2 => n3001, B1 => n3214, B2 => 
                           n3002, ZN => n1442);
   U2993 : OAI22_X1 port map( A1 => n2921, A2 => n3001, B1 => n3213, B2 => 
                           n3002, ZN => n1441);
   U2994 : OAI22_X1 port map( A1 => n2922, A2 => n3001, B1 => n3212, B2 => 
                           n3002, ZN => n1440);
   U2995 : OAI22_X1 port map( A1 => n2923, A2 => n3001, B1 => n3211, B2 => 
                           n3002, ZN => n1439);
   U2996 : OAI22_X1 port map( A1 => n2924, A2 => n3001, B1 => n3210, B2 => 
                           n3002, ZN => n1438);
   U2997 : OAI22_X1 port map( A1 => n2925, A2 => n3001, B1 => n3209, B2 => 
                           n3002, ZN => n1437);
   U2998 : OAI22_X1 port map( A1 => n2926, A2 => n3001, B1 => n3208, B2 => 
                           n3002, ZN => n1436);
   U2999 : OAI22_X1 port map( A1 => n2927, A2 => n3001, B1 => n3207, B2 => 
                           n3002, ZN => n1435);
   U3000 : OAI22_X1 port map( A1 => n2928, A2 => n3001, B1 => n3206, B2 => 
                           n3002, ZN => n1434);
   U3001 : OAI22_X1 port map( A1 => n2929, A2 => n3001, B1 => n3205, B2 => 
                           n3002, ZN => n1433);
   U3002 : OAI22_X1 port map( A1 => n2930, A2 => n3001, B1 => n3204, B2 => 
                           n3002, ZN => n1432);
   U3003 : OAI22_X1 port map( A1 => n2931, A2 => n3001, B1 => n3203, B2 => 
                           n3002, ZN => n1431);
   U3004 : NOR3_X1 port map( A1 => n2997, A2 => ADD_WR(2), A3 => n3000, ZN => 
                           n2942);
   U3005 : OAI22_X1 port map( A1 => n2899, A2 => n3003, B1 => n3202, B2 => 
                           n3004, ZN => n1430);
   U3006 : OAI22_X1 port map( A1 => n2901, A2 => n3003, B1 => n3201, B2 => 
                           n3004, ZN => n1429);
   U3007 : OAI22_X1 port map( A1 => n2902, A2 => n3003, B1 => n3200, B2 => 
                           n3004, ZN => n1428);
   U3008 : OAI22_X1 port map( A1 => n2903, A2 => n3003, B1 => n3199, B2 => 
                           n3004, ZN => n1427);
   U3009 : OAI22_X1 port map( A1 => n2904, A2 => n3003, B1 => n3198, B2 => 
                           n3004, ZN => n1426);
   U3010 : OAI22_X1 port map( A1 => n2905, A2 => n3003, B1 => n3197, B2 => 
                           n3004, ZN => n1425);
   U3011 : OAI22_X1 port map( A1 => n2906, A2 => n3003, B1 => n3196, B2 => 
                           n3004, ZN => n1424);
   U3012 : OAI22_X1 port map( A1 => n2907, A2 => n3003, B1 => n3195, B2 => 
                           n3004, ZN => n1423);
   U3013 : OAI22_X1 port map( A1 => n2908, A2 => n3003, B1 => n3194, B2 => 
                           n3004, ZN => n1422);
   U3014 : OAI22_X1 port map( A1 => n2909, A2 => n3003, B1 => n3193, B2 => 
                           n3004, ZN => n1421);
   U3015 : OAI22_X1 port map( A1 => n2910, A2 => n3003, B1 => n3192, B2 => 
                           n3004, ZN => n1420);
   U3016 : OAI22_X1 port map( A1 => n2911, A2 => n3003, B1 => n3191, B2 => 
                           n3004, ZN => n1419);
   U3017 : OAI22_X1 port map( A1 => n2912, A2 => n3003, B1 => n3190, B2 => 
                           n3004, ZN => n1418);
   U3018 : OAI22_X1 port map( A1 => n2913, A2 => n3003, B1 => n3189, B2 => 
                           n3004, ZN => n1417);
   U3019 : OAI22_X1 port map( A1 => n2914, A2 => n3003, B1 => n3188, B2 => 
                           n3004, ZN => n1416);
   U3020 : OAI22_X1 port map( A1 => n2915, A2 => n3003, B1 => n3187, B2 => 
                           n3004, ZN => n1415);
   U3021 : OAI22_X1 port map( A1 => n2916, A2 => n3003, B1 => n3186, B2 => 
                           n3004, ZN => n1414);
   U3022 : OAI22_X1 port map( A1 => n2917, A2 => n3003, B1 => n3185, B2 => 
                           n3004, ZN => n1413);
   U3023 : OAI22_X1 port map( A1 => n2918, A2 => n3003, B1 => n3184, B2 => 
                           n3004, ZN => n1412);
   U3024 : OAI22_X1 port map( A1 => n2919, A2 => n3003, B1 => n3183, B2 => 
                           n3004, ZN => n1411);
   U3025 : OAI22_X1 port map( A1 => n2920, A2 => n3003, B1 => n3182, B2 => 
                           n3004, ZN => n1410);
   U3026 : OAI22_X1 port map( A1 => n2921, A2 => n3003, B1 => n3181, B2 => 
                           n3004, ZN => n1409);
   U3027 : OAI22_X1 port map( A1 => n2922, A2 => n3003, B1 => n3180, B2 => 
                           n3004, ZN => n1408);
   U3028 : OAI22_X1 port map( A1 => n2923, A2 => n3003, B1 => n3179, B2 => 
                           n3004, ZN => n1407);
   U3029 : OAI22_X1 port map( A1 => n2924, A2 => n3003, B1 => n3178, B2 => 
                           n3004, ZN => n1406);
   U3030 : OAI22_X1 port map( A1 => n2925, A2 => n3003, B1 => n3177, B2 => 
                           n3004, ZN => n1405);
   U3031 : OAI22_X1 port map( A1 => n2926, A2 => n3003, B1 => n3176, B2 => 
                           n3004, ZN => n1404);
   U3032 : OAI22_X1 port map( A1 => n2927, A2 => n3003, B1 => n3175, B2 => 
                           n3004, ZN => n1403);
   U3033 : OAI22_X1 port map( A1 => n2928, A2 => n3003, B1 => n3174, B2 => 
                           n3004, ZN => n1402);
   U3034 : OAI22_X1 port map( A1 => n2929, A2 => n3003, B1 => n3173, B2 => 
                           n3004, ZN => n1401);
   U3035 : OAI22_X1 port map( A1 => n2930, A2 => n3003, B1 => n3172, B2 => 
                           n3004, ZN => n1400);
   U3036 : OAI22_X1 port map( A1 => n2931, A2 => n3003, B1 => n3171, B2 => 
                           n3004, ZN => n1399);
   U3037 : AND3_X1 port map( A1 => n2997, A2 => n3000, A3 => ADD_WR(2), ZN => 
                           n2945);
   U3038 : OAI22_X1 port map( A1 => n2899, A2 => n3005, B1 => n3170, B2 => 
                           n3006, ZN => n1398);
   U3039 : OAI22_X1 port map( A1 => n2901, A2 => n3005, B1 => n3169, B2 => 
                           n3006, ZN => n1397);
   U3040 : OAI22_X1 port map( A1 => n2902, A2 => n3005, B1 => n3168, B2 => 
                           n3006, ZN => n1396);
   U3041 : OAI22_X1 port map( A1 => n2903, A2 => n3005, B1 => n3167, B2 => 
                           n3006, ZN => n1395);
   U3042 : OAI22_X1 port map( A1 => n2904, A2 => n3005, B1 => n3166, B2 => 
                           n3006, ZN => n1394);
   U3043 : OAI22_X1 port map( A1 => n2905, A2 => n3005, B1 => n3165, B2 => 
                           n3006, ZN => n1393);
   U3044 : OAI22_X1 port map( A1 => n2906, A2 => n3005, B1 => n3164, B2 => 
                           n3006, ZN => n1392);
   U3045 : OAI22_X1 port map( A1 => n2907, A2 => n3005, B1 => n3163, B2 => 
                           n3006, ZN => n1391);
   U3046 : OAI22_X1 port map( A1 => n2908, A2 => n3005, B1 => n3162, B2 => 
                           n3006, ZN => n1390);
   U3047 : OAI22_X1 port map( A1 => n2909, A2 => n3005, B1 => n3161, B2 => 
                           n3006, ZN => n1389);
   U3048 : OAI22_X1 port map( A1 => n2910, A2 => n3005, B1 => n3160, B2 => 
                           n3006, ZN => n1388);
   U3049 : OAI22_X1 port map( A1 => n2911, A2 => n3005, B1 => n3159, B2 => 
                           n3006, ZN => n1387);
   U3050 : OAI22_X1 port map( A1 => n2912, A2 => n3005, B1 => n3158, B2 => 
                           n3006, ZN => n1386);
   U3051 : OAI22_X1 port map( A1 => n2913, A2 => n3005, B1 => n3157, B2 => 
                           n3006, ZN => n1385);
   U3052 : OAI22_X1 port map( A1 => n2914, A2 => n3005, B1 => n3156, B2 => 
                           n3006, ZN => n1384);
   U3053 : OAI22_X1 port map( A1 => n2915, A2 => n3005, B1 => n3155, B2 => 
                           n3006, ZN => n1383);
   U3054 : OAI22_X1 port map( A1 => n2916, A2 => n3005, B1 => n3154, B2 => 
                           n3006, ZN => n1382);
   U3055 : OAI22_X1 port map( A1 => n2917, A2 => n3005, B1 => n3153, B2 => 
                           n3006, ZN => n1381);
   U3056 : OAI22_X1 port map( A1 => n2918, A2 => n3005, B1 => n3152, B2 => 
                           n3006, ZN => n1380);
   U3057 : OAI22_X1 port map( A1 => n2919, A2 => n3005, B1 => n3151, B2 => 
                           n3006, ZN => n1379);
   U3058 : OAI22_X1 port map( A1 => n2920, A2 => n3005, B1 => n3150, B2 => 
                           n3006, ZN => n1378);
   U3059 : OAI22_X1 port map( A1 => n2921, A2 => n3005, B1 => n3149, B2 => 
                           n3006, ZN => n1377);
   U3060 : OAI22_X1 port map( A1 => n2922, A2 => n3005, B1 => n3148, B2 => 
                           n3006, ZN => n1376);
   U3061 : OAI22_X1 port map( A1 => n2923, A2 => n3005, B1 => n3147, B2 => 
                           n3006, ZN => n1375);
   U3062 : OAI22_X1 port map( A1 => n2924, A2 => n3005, B1 => n3146, B2 => 
                           n3006, ZN => n1374);
   U3063 : OAI22_X1 port map( A1 => n2925, A2 => n3005, B1 => n3145, B2 => 
                           n3006, ZN => n1373);
   U3064 : OAI22_X1 port map( A1 => n2926, A2 => n3005, B1 => n3144, B2 => 
                           n3006, ZN => n1372);
   U3065 : OAI22_X1 port map( A1 => n2927, A2 => n3005, B1 => n3143, B2 => 
                           n3006, ZN => n1371);
   U3066 : OAI22_X1 port map( A1 => n2928, A2 => n3005, B1 => n3142, B2 => 
                           n3006, ZN => n1370);
   U3067 : OAI22_X1 port map( A1 => n2929, A2 => n3005, B1 => n3141, B2 => 
                           n3006, ZN => n1369);
   U3068 : OAI22_X1 port map( A1 => n2930, A2 => n3005, B1 => n3140, B2 => 
                           n3006, ZN => n1368);
   U3069 : OAI22_X1 port map( A1 => n2931, A2 => n3005, B1 => n3139, B2 => 
                           n3006, ZN => n1367);
   U3070 : AND3_X1 port map( A1 => ADD_WR(0), A2 => n3000, A3 => ADD_WR(2), ZN 
                           => n2948);
   U3071 : INV_X1 port map( A => ADD_WR(1), ZN => n3000);
   U3072 : OAI22_X1 port map( A1 => n2899, A2 => n3007, B1 => n3138, B2 => 
                           n3008, ZN => n1366);
   U3073 : OAI22_X1 port map( A1 => n2901, A2 => n3007, B1 => n3137, B2 => 
                           n3008, ZN => n1365);
   U3074 : OAI22_X1 port map( A1 => n2902, A2 => n3007, B1 => n3136, B2 => 
                           n3008, ZN => n1364);
   U3075 : OAI22_X1 port map( A1 => n2903, A2 => n3007, B1 => n3135, B2 => 
                           n3008, ZN => n1363);
   U3076 : OAI22_X1 port map( A1 => n2904, A2 => n3007, B1 => n3134, B2 => 
                           n3008, ZN => n1362);
   U3077 : OAI22_X1 port map( A1 => n2905, A2 => n3007, B1 => n3133, B2 => 
                           n3008, ZN => n1361);
   U3078 : OAI22_X1 port map( A1 => n2906, A2 => n3007, B1 => n3132, B2 => 
                           n3008, ZN => n1360);
   U3079 : OAI22_X1 port map( A1 => n2907, A2 => n3007, B1 => n3131, B2 => 
                           n3008, ZN => n1359);
   U3080 : OAI22_X1 port map( A1 => n2908, A2 => n3007, B1 => n3130, B2 => 
                           n3008, ZN => n1358);
   U3081 : OAI22_X1 port map( A1 => n2909, A2 => n3007, B1 => n3129, B2 => 
                           n3008, ZN => n1357);
   U3082 : OAI22_X1 port map( A1 => n2910, A2 => n3007, B1 => n3128, B2 => 
                           n3008, ZN => n1356);
   U3083 : OAI22_X1 port map( A1 => n2911, A2 => n3007, B1 => n3127, B2 => 
                           n3008, ZN => n1355);
   U3084 : OAI22_X1 port map( A1 => n2912, A2 => n3007, B1 => n3126, B2 => 
                           n3008, ZN => n1354);
   U3085 : OAI22_X1 port map( A1 => n2913, A2 => n3007, B1 => n3125, B2 => 
                           n3008, ZN => n1353);
   U3086 : OAI22_X1 port map( A1 => n2914, A2 => n3007, B1 => n3124, B2 => 
                           n3008, ZN => n1352);
   U3087 : OAI22_X1 port map( A1 => n2915, A2 => n3007, B1 => n3123, B2 => 
                           n3008, ZN => n1351);
   U3088 : OAI22_X1 port map( A1 => n2916, A2 => n3007, B1 => n3122, B2 => 
                           n3008, ZN => n1350);
   U3089 : OAI22_X1 port map( A1 => n2917, A2 => n3007, B1 => n3121, B2 => 
                           n3008, ZN => n1349);
   U3090 : OAI22_X1 port map( A1 => n2918, A2 => n3007, B1 => n3120, B2 => 
                           n3008, ZN => n1348);
   U3091 : OAI22_X1 port map( A1 => n2919, A2 => n3007, B1 => n3119, B2 => 
                           n3008, ZN => n1347);
   U3092 : OAI22_X1 port map( A1 => n2920, A2 => n3007, B1 => n3118, B2 => 
                           n3008, ZN => n1346);
   U3093 : OAI22_X1 port map( A1 => n2921, A2 => n3007, B1 => n3117, B2 => 
                           n3008, ZN => n1345);
   U3094 : OAI22_X1 port map( A1 => n2922, A2 => n3007, B1 => n3116, B2 => 
                           n3008, ZN => n1344);
   U3095 : OAI22_X1 port map( A1 => n2923, A2 => n3007, B1 => n3115, B2 => 
                           n3008, ZN => n1343);
   U3096 : OAI22_X1 port map( A1 => n2924, A2 => n3007, B1 => n3114, B2 => 
                           n3008, ZN => n1342);
   U3097 : OAI22_X1 port map( A1 => n2925, A2 => n3007, B1 => n3113, B2 => 
                           n3008, ZN => n1341);
   U3098 : OAI22_X1 port map( A1 => n2926, A2 => n3007, B1 => n3112, B2 => 
                           n3008, ZN => n1340);
   U3099 : OAI22_X1 port map( A1 => n2927, A2 => n3007, B1 => n3111, B2 => 
                           n3008, ZN => n1339);
   U3100 : OAI22_X1 port map( A1 => n2928, A2 => n3007, B1 => n3110, B2 => 
                           n3008, ZN => n1338);
   U3101 : OAI22_X1 port map( A1 => n2929, A2 => n3007, B1 => n3109, B2 => 
                           n3008, ZN => n1337);
   U3102 : OAI22_X1 port map( A1 => n2930, A2 => n3007, B1 => n3108, B2 => 
                           n3008, ZN => n1336);
   U3103 : OAI22_X1 port map( A1 => n2931, A2 => n3007, B1 => n3107, B2 => 
                           n3008, ZN => n1335);
   U3104 : AND3_X1 port map( A1 => ADD_WR(1), A2 => n2997, A3 => ADD_WR(2), ZN 
                           => n2951);
   U3105 : INV_X1 port map( A => ADD_WR(0), ZN => n2997);
   U3106 : OAI22_X1 port map( A1 => n2899, A2 => n3009, B1 => n3106, B2 => 
                           n3010, ZN => n1334);
   U3107 : OAI22_X1 port map( A1 => n2901, A2 => n3009, B1 => n3105, B2 => 
                           n3010, ZN => n1333);
   U3108 : OAI22_X1 port map( A1 => n2902, A2 => n3009, B1 => n3104, B2 => 
                           n3010, ZN => n1332);
   U3109 : OAI22_X1 port map( A1 => n2903, A2 => n3009, B1 => n3103, B2 => 
                           n3010, ZN => n1331);
   U3110 : OAI22_X1 port map( A1 => n2904, A2 => n3009, B1 => n3102, B2 => 
                           n3010, ZN => n1330);
   U3111 : OAI22_X1 port map( A1 => n2905, A2 => n3009, B1 => n3101, B2 => 
                           n3010, ZN => n1329);
   U3112 : OAI22_X1 port map( A1 => n2906, A2 => n3009, B1 => n3100, B2 => 
                           n3010, ZN => n1328);
   U3113 : OAI22_X1 port map( A1 => n2907, A2 => n3009, B1 => n3099, B2 => 
                           n3010, ZN => n1327);
   U3114 : OAI22_X1 port map( A1 => n2908, A2 => n3009, B1 => n3098, B2 => 
                           n3010, ZN => n1326);
   U3115 : OAI22_X1 port map( A1 => n2909, A2 => n3009, B1 => n3097, B2 => 
                           n3010, ZN => n1325);
   U3116 : OAI22_X1 port map( A1 => n2910, A2 => n3009, B1 => n3096, B2 => 
                           n3010, ZN => n1324);
   U3117 : OAI22_X1 port map( A1 => n2911, A2 => n3009, B1 => n3095, B2 => 
                           n3010, ZN => n1323);
   U3118 : OAI22_X1 port map( A1 => n2912, A2 => n3009, B1 => n3094, B2 => 
                           n3010, ZN => n1322);
   U3119 : OAI22_X1 port map( A1 => n2913, A2 => n3009, B1 => n3093, B2 => 
                           n3010, ZN => n1321);
   U3120 : OAI22_X1 port map( A1 => n2914, A2 => n3009, B1 => n3092, B2 => 
                           n3010, ZN => n1320);
   U3121 : OAI22_X1 port map( A1 => n2915, A2 => n3009, B1 => n3091, B2 => 
                           n3010, ZN => n1319);
   U3122 : OAI22_X1 port map( A1 => n2916, A2 => n3009, B1 => n3090, B2 => 
                           n3010, ZN => n1318);
   U3123 : OAI22_X1 port map( A1 => n2917, A2 => n3009, B1 => n3089, B2 => 
                           n3010, ZN => n1317);
   U3124 : OAI22_X1 port map( A1 => n2918, A2 => n3009, B1 => n3088, B2 => 
                           n3010, ZN => n1316);
   U3125 : OAI22_X1 port map( A1 => n2919, A2 => n3009, B1 => n3087, B2 => 
                           n3010, ZN => n1315);
   U3126 : OAI22_X1 port map( A1 => n2920, A2 => n3009, B1 => n3086, B2 => 
                           n3010, ZN => n1314);
   U3127 : OAI22_X1 port map( A1 => n2921, A2 => n3009, B1 => n3085, B2 => 
                           n3010, ZN => n1313);
   U3128 : OAI22_X1 port map( A1 => n2922, A2 => n3009, B1 => n3084, B2 => 
                           n3010, ZN => n1312);
   U3129 : OAI22_X1 port map( A1 => n2923, A2 => n3009, B1 => n3083, B2 => 
                           n3010, ZN => n1311);
   U3130 : OAI22_X1 port map( A1 => n2924, A2 => n3009, B1 => n3082, B2 => 
                           n3010, ZN => n1310);
   U3131 : OAI22_X1 port map( A1 => n2925, A2 => n3009, B1 => n3081, B2 => 
                           n3010, ZN => n1309);
   U3132 : OAI22_X1 port map( A1 => n2926, A2 => n3009, B1 => n3080, B2 => 
                           n3010, ZN => n1308);
   U3133 : OAI22_X1 port map( A1 => n2927, A2 => n3009, B1 => n3079, B2 => 
                           n3010, ZN => n1307);
   U3134 : OAI22_X1 port map( A1 => n2928, A2 => n3009, B1 => n3078, B2 => 
                           n3010, ZN => n1306);
   U3135 : OAI22_X1 port map( A1 => n2929, A2 => n3009, B1 => n3077, B2 => 
                           n3010, ZN => n1305);
   U3136 : OAI22_X1 port map( A1 => n2930, A2 => n3009, B1 => n3076, B2 => 
                           n3010, ZN => n1304);
   U3137 : OAI22_X1 port map( A1 => n2931, A2 => n3009, B1 => n3075, B2 => 
                           n3010, ZN => n1303);
   U3138 : AND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2),
                           ZN => n2954);
   U3139 : AND3_X1 port map( A1 => ADD_WR(3), A2 => n2957, A3 => ADD_WR(4), ZN 
                           => n2994);
   U3140 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n2957);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity SIGN_EXT_bits16 is

   port( inputt : in std_logic_vector (15 downto 0);  outputt : out 
         std_logic_vector (31 downto 0));

end SIGN_EXT_bits16;

architecture SYN_BEHAVIORAL of SIGN_EXT_bits16 is

begin
   outputt <= ( inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), 
      inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), 
      inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), 
      inputt(14), inputt(13), inputt(12), inputt(11), inputt(10), inputt(9), 
      inputt(8), inputt(7), inputt(6), inputt(5), inputt(4), inputt(3), 
      inputt(2), inputt(1), inputt(0) );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_0 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_0;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_321
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_322
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_323
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_324
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_325
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_326
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_327
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_328
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_329
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_330
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_331
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_332
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_333
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_334
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_335
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_336
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_337
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_338
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_339
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_340
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_341
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_342
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_343
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_344
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_345
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_346
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_347
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_348
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_349
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_350
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_351
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_352
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FF_0 : FD_352 port map( D => data_in(0), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_351 port map( D => data_in(1), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_350 port map( D => data_in(2), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_349 port map( D => data_in(3), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_348 port map( D => data_in(4), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_347 port map( D => data_in(5), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_346 port map( D => data_in(6), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_345 port map( D => data_in(7), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_344 port map( D => data_in(8), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_343 port map( D => data_in(9), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_342 port map( D => data_in(10), CK => n5, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_341 port map( D => data_in(11), CK => n6, RESET => n1, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_340 port map( D => data_in(12), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(12));
   FF_13 : FD_339 port map( D => data_in(13), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(13));
   FF_14 : FD_338 port map( D => data_in(14), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(14));
   FF_15 : FD_337 port map( D => data_in(15), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(15));
   FF_16 : FD_336 port map( D => data_in(16), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(16));
   FF_17 : FD_335 port map( D => data_in(17), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(17));
   FF_18 : FD_334 port map( D => data_in(18), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(18));
   FF_19 : FD_333 port map( D => data_in(19), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(19));
   FF_20 : FD_332 port map( D => data_in(20), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(20));
   FF_21 : FD_331 port map( D => data_in(21), CK => n6, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(21));
   FF_22 : FD_330 port map( D => data_in(22), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(22));
   FF_23 : FD_329 port map( D => data_in(23), CK => n7, RESET => n2, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_328 port map( D => data_in(24), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_327 port map( D => data_in(25), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_326 port map( D => data_in(26), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_325 port map( D => data_in(27), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_324 port map( D => data_in(28), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_323 port map( D => data_in(29), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_322 port map( D => data_in(30), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_321 port map( D => data_in(31), CK => n7, RESET => n3, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n4);
   U2 : BUF_X1 port map( A => CK, Z => n8);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end RCA_NBITS32;

architecture SYN_BEHAVIORAL of RCA_NBITS32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174 : 
      std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S(9));
   U3 : XNOR2_X1 port map( A => A(9), B => n3, ZN => n2);
   U4 : XNOR2_X1 port map( A => B(9), B => Ci, ZN => n1);
   U5 : XOR2_X1 port map( A => n4, B => n5, Z => S(8));
   U6 : XNOR2_X1 port map( A => n6, B => A(8), ZN => n5);
   U7 : XNOR2_X1 port map( A => B(8), B => Ci, ZN => n4);
   U8 : XOR2_X1 port map( A => n7, B => n8, Z => S(7));
   U9 : XNOR2_X1 port map( A => n9, B => A(7), ZN => n8);
   U10 : XNOR2_X1 port map( A => B(7), B => Ci, ZN => n7);
   U11 : XOR2_X1 port map( A => n10, B => n11, Z => S(6));
   U12 : XNOR2_X1 port map( A => n12, B => A(6), ZN => n11);
   U13 : XNOR2_X1 port map( A => B(6), B => Ci, ZN => n10);
   U14 : XOR2_X1 port map( A => n13, B => n14, Z => S(5));
   U15 : XNOR2_X1 port map( A => A(5), B => n15, ZN => n14);
   U16 : XNOR2_X1 port map( A => B(5), B => Ci, ZN => n13);
   U17 : XOR2_X1 port map( A => n16, B => n17, Z => S(4));
   U18 : XNOR2_X1 port map( A => n18, B => A(4), ZN => n17);
   U19 : XNOR2_X1 port map( A => B(4), B => Ci, ZN => n16);
   U20 : XOR2_X1 port map( A => n19, B => n20, Z => S(3));
   U21 : XOR2_X1 port map( A => A(3), B => n21, Z => n20);
   U22 : XOR2_X1 port map( A => Ci, B => B(3), Z => n19);
   U23 : XOR2_X1 port map( A => n22, B => n23, Z => S(31));
   U24 : XNOR2_X1 port map( A => n24, B => A(31), ZN => n23);
   U25 : XNOR2_X1 port map( A => B(31), B => Ci, ZN => n22);
   U26 : XOR2_X1 port map( A => n25, B => n26, Z => S(30));
   U27 : XOR2_X1 port map( A => Ci, B => B(30), Z => n26);
   U28 : XNOR2_X1 port map( A => A(30), B => n27, ZN => n25);
   U29 : XOR2_X1 port map( A => n28, B => n29, Z => S(2));
   U30 : XNOR2_X1 port map( A => A(2), B => n30, ZN => n29);
   U31 : XNOR2_X1 port map( A => B(2), B => Ci, ZN => n28);
   U32 : XOR2_X1 port map( A => n31, B => n32, Z => S(29));
   U33 : XNOR2_X1 port map( A => n33, B => A(29), ZN => n32);
   U34 : XNOR2_X1 port map( A => B(29), B => Ci, ZN => n31);
   U35 : XOR2_X1 port map( A => n34, B => n35, Z => S(28));
   U36 : XNOR2_X1 port map( A => n36, B => A(28), ZN => n35);
   U37 : XNOR2_X1 port map( A => B(28), B => Ci, ZN => n34);
   U38 : XOR2_X1 port map( A => n37, B => n38, Z => S(27));
   U39 : XNOR2_X1 port map( A => n39, B => A(27), ZN => n38);
   U40 : XNOR2_X1 port map( A => B(27), B => Ci, ZN => n37);
   U41 : XOR2_X1 port map( A => n40, B => n41, Z => S(26));
   U42 : XNOR2_X1 port map( A => n42, B => A(26), ZN => n41);
   U43 : XNOR2_X1 port map( A => B(26), B => Ci, ZN => n40);
   U44 : XOR2_X1 port map( A => n43, B => n44, Z => S(25));
   U45 : XNOR2_X1 port map( A => n45, B => A(25), ZN => n44);
   U46 : XNOR2_X1 port map( A => B(25), B => Ci, ZN => n43);
   U47 : XOR2_X1 port map( A => n46, B => n47, Z => S(24));
   U48 : XNOR2_X1 port map( A => n48, B => A(24), ZN => n47);
   U49 : XNOR2_X1 port map( A => B(24), B => Ci, ZN => n46);
   U50 : XOR2_X1 port map( A => n49, B => n50, Z => S(23));
   U51 : XNOR2_X1 port map( A => n51, B => A(23), ZN => n50);
   U52 : XNOR2_X1 port map( A => B(23), B => Ci, ZN => n49);
   U53 : XOR2_X1 port map( A => n52, B => n53, Z => S(22));
   U54 : XNOR2_X1 port map( A => n54, B => A(22), ZN => n53);
   U55 : XNOR2_X1 port map( A => B(22), B => Ci, ZN => n52);
   U56 : XOR2_X1 port map( A => n55, B => n56, Z => S(21));
   U57 : XNOR2_X1 port map( A => n57, B => A(21), ZN => n56);
   U58 : XNOR2_X1 port map( A => B(21), B => Ci, ZN => n55);
   U59 : XOR2_X1 port map( A => n58, B => n59, Z => S(20));
   U60 : XNOR2_X1 port map( A => n60, B => A(20), ZN => n59);
   U61 : XNOR2_X1 port map( A => B(20), B => Ci, ZN => n58);
   U62 : XOR2_X1 port map( A => n61, B => n62, Z => S(1));
   U63 : XNOR2_X1 port map( A => n63, B => n64, ZN => n62);
   U64 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n61);
   U65 : XOR2_X1 port map( A => n65, B => n66, Z => S(19));
   U66 : XNOR2_X1 port map( A => n67, B => A(19), ZN => n66);
   U67 : XNOR2_X1 port map( A => B(19), B => Ci, ZN => n65);
   U68 : XOR2_X1 port map( A => n68, B => n69, Z => S(18));
   U69 : XNOR2_X1 port map( A => n70, B => A(18), ZN => n69);
   U70 : XNOR2_X1 port map( A => B(18), B => Ci, ZN => n68);
   U71 : XOR2_X1 port map( A => n71, B => n72, Z => S(17));
   U72 : XNOR2_X1 port map( A => n73, B => A(17), ZN => n72);
   U73 : XNOR2_X1 port map( A => B(17), B => Ci, ZN => n71);
   U74 : XOR2_X1 port map( A => n74, B => n75, Z => S(16));
   U75 : XNOR2_X1 port map( A => n76, B => A(16), ZN => n75);
   U76 : XNOR2_X1 port map( A => B(16), B => Ci, ZN => n74);
   U77 : XOR2_X1 port map( A => n77, B => n78, Z => S(15));
   U78 : XNOR2_X1 port map( A => n79, B => A(15), ZN => n78);
   U79 : XNOR2_X1 port map( A => B(15), B => Ci, ZN => n77);
   U80 : XOR2_X1 port map( A => n80, B => n81, Z => S(14));
   U81 : XNOR2_X1 port map( A => n82, B => A(14), ZN => n81);
   U82 : XNOR2_X1 port map( A => B(14), B => Ci, ZN => n80);
   U83 : XOR2_X1 port map( A => n83, B => n84, Z => S(13));
   U84 : XNOR2_X1 port map( A => n85, B => A(13), ZN => n84);
   U85 : XNOR2_X1 port map( A => B(13), B => Ci, ZN => n83);
   U86 : XOR2_X1 port map( A => n86, B => n87, Z => S(12));
   U87 : XNOR2_X1 port map( A => n88, B => A(12), ZN => n87);
   U88 : XNOR2_X1 port map( A => B(12), B => Ci, ZN => n86);
   U89 : XOR2_X1 port map( A => n89, B => n90, Z => S(11));
   U90 : XNOR2_X1 port map( A => n91, B => A(11), ZN => n90);
   U91 : XNOR2_X1 port map( A => B(11), B => Ci, ZN => n89);
   U92 : XOR2_X1 port map( A => n92, B => n93, Z => S(10));
   U93 : XNOR2_X1 port map( A => n94, B => A(10), ZN => n93);
   U94 : XNOR2_X1 port map( A => B(10), B => Ci, ZN => n92);
   U95 : MUX2_X1 port map( A => n95, B => n96, S => Ci, Z => S(0));
   U96 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n63, ZN => n96);
   U97 : XOR2_X1 port map( A => B(0), B => A(0), Z => n95);
   U98 : OAI21_X1 port map( B1 => n97, B2 => n98, A => n99, ZN => Co);
   U99 : OAI21_X1 port map( B1 => n24, B2 => A(31), A => B(31), ZN => n99);
   U100 : INV_X1 port map( A => n98, ZN => n24);
   U101 : OAI22_X1 port map( A1 => A(30), A2 => n100, B1 => B(30), B2 => n101, 
                           ZN => n98);
   U102 : AND2_X1 port map( A1 => n100, A2 => A(30), ZN => n101);
   U103 : INV_X1 port map( A => n27, ZN => n100);
   U104 : AOI21_X1 port map( B1 => n33, B2 => A(29), A => n102, ZN => n27);
   U105 : INV_X1 port map( A => n103, ZN => n102);
   U106 : OAI21_X1 port map( B1 => n33, B2 => A(29), A => B(29), ZN => n103);
   U107 : AOI21_X1 port map( B1 => n104, B2 => n105, A => n106, ZN => n33);
   U108 : AOI21_X1 port map( B1 => n36, B2 => A(28), A => B(28), ZN => n106);
   U109 : INV_X1 port map( A => n36, ZN => n105);
   U110 : AOI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => n36);
   U111 : AOI21_X1 port map( B1 => n39, B2 => A(27), A => B(27), ZN => n109);
   U112 : INV_X1 port map( A => n39, ZN => n108);
   U113 : AOI21_X1 port map( B1 => n110, B2 => n111, A => n112, ZN => n39);
   U114 : AOI21_X1 port map( B1 => n42, B2 => A(26), A => B(26), ZN => n112);
   U115 : INV_X1 port map( A => n42, ZN => n111);
   U116 : AOI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n42);
   U117 : AOI21_X1 port map( B1 => n45, B2 => A(25), A => B(25), ZN => n115);
   U118 : INV_X1 port map( A => n45, ZN => n114);
   U119 : AOI21_X1 port map( B1 => n116, B2 => n117, A => n118, ZN => n45);
   U120 : AOI21_X1 port map( B1 => n48, B2 => A(24), A => B(24), ZN => n118);
   U121 : INV_X1 port map( A => n48, ZN => n117);
   U122 : AOI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n48);
   U123 : AOI21_X1 port map( B1 => n51, B2 => A(23), A => B(23), ZN => n121);
   U124 : INV_X1 port map( A => n51, ZN => n120);
   U125 : AOI21_X1 port map( B1 => n122, B2 => n123, A => n124, ZN => n51);
   U126 : AOI21_X1 port map( B1 => n54, B2 => A(22), A => B(22), ZN => n124);
   U127 : INV_X1 port map( A => n54, ZN => n123);
   U128 : AOI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n54);
   U129 : AOI21_X1 port map( B1 => n57, B2 => A(21), A => B(21), ZN => n127);
   U130 : INV_X1 port map( A => n57, ZN => n126);
   U131 : AOI21_X1 port map( B1 => n128, B2 => n129, A => n130, ZN => n57);
   U132 : AOI21_X1 port map( B1 => n60, B2 => A(20), A => B(20), ZN => n130);
   U133 : INV_X1 port map( A => n60, ZN => n129);
   U134 : AOI21_X1 port map( B1 => n131, B2 => n132, A => n133, ZN => n60);
   U135 : AOI21_X1 port map( B1 => n67, B2 => A(19), A => B(19), ZN => n133);
   U136 : INV_X1 port map( A => n67, ZN => n132);
   U137 : AOI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n67);
   U138 : AOI21_X1 port map( B1 => n70, B2 => A(18), A => B(18), ZN => n136);
   U139 : INV_X1 port map( A => n70, ZN => n135);
   U140 : AOI21_X1 port map( B1 => n137, B2 => n138, A => n139, ZN => n70);
   U141 : AOI21_X1 port map( B1 => n73, B2 => A(17), A => B(17), ZN => n139);
   U142 : INV_X1 port map( A => n73, ZN => n138);
   U143 : AOI21_X1 port map( B1 => n140, B2 => n141, A => n142, ZN => n73);
   U144 : AOI21_X1 port map( B1 => n76, B2 => A(16), A => B(16), ZN => n142);
   U145 : INV_X1 port map( A => n141, ZN => n76);
   U146 : OAI22_X1 port map( A1 => A(15), A2 => n79, B1 => B(15), B2 => n143, 
                           ZN => n141);
   U147 : AND2_X1 port map( A1 => n79, A2 => A(15), ZN => n143);
   U148 : INV_X1 port map( A => n144, ZN => n79);
   U149 : OAI22_X1 port map( A1 => A(14), A2 => n82, B1 => B(14), B2 => n145, 
                           ZN => n144);
   U150 : AND2_X1 port map( A1 => n82, A2 => A(14), ZN => n145);
   U151 : INV_X1 port map( A => n146, ZN => n82);
   U152 : OAI22_X1 port map( A1 => A(13), A2 => n85, B1 => B(13), B2 => n147, 
                           ZN => n146);
   U153 : AND2_X1 port map( A1 => n85, A2 => A(13), ZN => n147);
   U154 : INV_X1 port map( A => n148, ZN => n85);
   U155 : OAI22_X1 port map( A1 => A(12), A2 => n88, B1 => B(12), B2 => n149, 
                           ZN => n148);
   U156 : AND2_X1 port map( A1 => n88, A2 => A(12), ZN => n149);
   U157 : INV_X1 port map( A => n150, ZN => n88);
   U158 : OAI22_X1 port map( A1 => A(11), A2 => n91, B1 => B(11), B2 => n151, 
                           ZN => n150);
   U159 : AND2_X1 port map( A1 => n91, A2 => A(11), ZN => n151);
   U160 : AOI21_X1 port map( B1 => n152, B2 => n153, A => n154, ZN => n91);
   U161 : AOI21_X1 port map( B1 => n94, B2 => A(10), A => B(10), ZN => n154);
   U162 : INV_X1 port map( A => n153, ZN => n94);
   U163 : OAI21_X1 port map( B1 => A(9), B2 => n3, A => n155, ZN => n153);
   U164 : INV_X1 port map( A => n156, ZN => n155);
   U165 : AOI21_X1 port map( B1 => n3, B2 => A(9), A => B(9), ZN => n156);
   U166 : OAI21_X1 port map( B1 => n157, B2 => n158, A => n159, ZN => n3);
   U167 : OAI21_X1 port map( B1 => n6, B2 => A(8), A => B(8), ZN => n159);
   U168 : INV_X1 port map( A => n157, ZN => n6);
   U169 : INV_X1 port map( A => A(8), ZN => n158);
   U170 : OAI22_X1 port map( A1 => A(7), A2 => n9, B1 => B(7), B2 => n160, ZN 
                           => n157);
   U171 : AND2_X1 port map( A1 => n9, A2 => A(7), ZN => n160);
   U172 : AOI21_X1 port map( B1 => n161, B2 => n162, A => n163, ZN => n9);
   U173 : AOI21_X1 port map( B1 => n12, B2 => A(6), A => B(6), ZN => n163);
   U174 : INV_X1 port map( A => n162, ZN => n12);
   U175 : OAI21_X1 port map( B1 => A(5), B2 => n15, A => n164, ZN => n162);
   U176 : INV_X1 port map( A => n165, ZN => n164);
   U177 : AOI21_X1 port map( B1 => n15, B2 => A(5), A => B(5), ZN => n165);
   U178 : OAI21_X1 port map( B1 => n166, B2 => n167, A => n168, ZN => n15);
   U179 : OAI21_X1 port map( B1 => n18, B2 => A(4), A => B(4), ZN => n168);
   U180 : INV_X1 port map( A => n166, ZN => n18);
   U181 : INV_X1 port map( A => A(4), ZN => n167);
   U182 : OAI22_X1 port map( A1 => A(3), A2 => n21, B1 => B(3), B2 => n169, ZN 
                           => n166);
   U183 : AND2_X1 port map( A1 => n21, A2 => A(3), ZN => n169);
   U184 : AOI21_X1 port map( B1 => n170, B2 => n171, A => n172, ZN => n21);
   U185 : AOI21_X1 port map( B1 => n30, B2 => A(2), A => B(2), ZN => n172);
   U186 : INV_X1 port map( A => n30, ZN => n171);
   U187 : OAI22_X1 port map( A1 => n64, A2 => n173, B1 => n174, B2 => n63, ZN 
                           => n30);
   U188 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n63);
   U189 : NOR2_X1 port map( A1 => B(1), A2 => A(1), ZN => n174);
   U190 : INV_X1 port map( A => B(1), ZN => n173);
   U191 : INV_X1 port map( A => A(1), ZN => n64);
   U192 : INV_X1 port map( A => A(2), ZN => n170);
   U193 : INV_X1 port map( A => A(6), ZN => n161);
   U194 : INV_X1 port map( A => A(10), ZN => n152);
   U195 : INV_X1 port map( A => A(16), ZN => n140);
   U196 : INV_X1 port map( A => A(17), ZN => n137);
   U197 : INV_X1 port map( A => A(18), ZN => n134);
   U198 : INV_X1 port map( A => A(19), ZN => n131);
   U199 : INV_X1 port map( A => A(20), ZN => n128);
   U200 : INV_X1 port map( A => A(21), ZN => n125);
   U201 : INV_X1 port map( A => A(22), ZN => n122);
   U202 : INV_X1 port map( A => A(23), ZN => n119);
   U203 : INV_X1 port map( A => A(24), ZN => n116);
   U204 : INV_X1 port map( A => A(25), ZN => n113);
   U205 : INV_X1 port map( A => A(26), ZN => n110);
   U206 : INV_X1 port map( A => A(27), ZN => n107);
   U207 : INV_X1 port map( A => A(28), ZN => n104);
   U208 : INV_X1 port map( A => A(31), ZN => n97);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity writeBack_nbits32 is

   port( LMD_OUT, ALUREG_OUTPUT : in std_logic_vector (31 downto 0);  
         WB_MUX_SEL : in std_logic;  DATAIN_RF : out std_logic_vector (31 
         downto 0));

end writeBack_nbits32;

architecture SYN_STRUCTURAL of writeBack_nbits32 is

   component MUX21_GENERIC_bits32_1
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;

begin
   
   MUXWB : MUX21_GENERIC_bits32_1 port map( A(31) => ALUREG_OUTPUT(31), A(30) 
                           => ALUREG_OUTPUT(30), A(29) => ALUREG_OUTPUT(29), 
                           A(28) => ALUREG_OUTPUT(28), A(27) => 
                           ALUREG_OUTPUT(27), A(26) => ALUREG_OUTPUT(26), A(25)
                           => ALUREG_OUTPUT(25), A(24) => ALUREG_OUTPUT(24), 
                           A(23) => ALUREG_OUTPUT(23), A(22) => 
                           ALUREG_OUTPUT(22), A(21) => ALUREG_OUTPUT(21), A(20)
                           => ALUREG_OUTPUT(20), A(19) => ALUREG_OUTPUT(19), 
                           A(18) => ALUREG_OUTPUT(18), A(17) => 
                           ALUREG_OUTPUT(17), A(16) => ALUREG_OUTPUT(16), A(15)
                           => ALUREG_OUTPUT(15), A(14) => ALUREG_OUTPUT(14), 
                           A(13) => ALUREG_OUTPUT(13), A(12) => 
                           ALUREG_OUTPUT(12), A(11) => ALUREG_OUTPUT(11), A(10)
                           => ALUREG_OUTPUT(10), A(9) => ALUREG_OUTPUT(9), A(8)
                           => ALUREG_OUTPUT(8), A(7) => ALUREG_OUTPUT(7), A(6) 
                           => ALUREG_OUTPUT(6), A(5) => ALUREG_OUTPUT(5), A(4) 
                           => ALUREG_OUTPUT(4), A(3) => ALUREG_OUTPUT(3), A(2) 
                           => ALUREG_OUTPUT(2), A(1) => ALUREG_OUTPUT(1), A(0) 
                           => ALUREG_OUTPUT(0), B(31) => LMD_OUT(31), B(30) => 
                           LMD_OUT(30), B(29) => LMD_OUT(29), B(28) => 
                           LMD_OUT(28), B(27) => LMD_OUT(27), B(26) => 
                           LMD_OUT(26), B(25) => LMD_OUT(25), B(24) => 
                           LMD_OUT(24), B(23) => LMD_OUT(23), B(22) => 
                           LMD_OUT(22), B(21) => LMD_OUT(21), B(20) => 
                           LMD_OUT(20), B(19) => LMD_OUT(19), B(18) => 
                           LMD_OUT(18), B(17) => LMD_OUT(17), B(16) => 
                           LMD_OUT(16), B(15) => LMD_OUT(15), B(14) => 
                           LMD_OUT(14), B(13) => LMD_OUT(13), B(12) => 
                           LMD_OUT(12), B(11) => LMD_OUT(11), B(10) => 
                           LMD_OUT(10), B(9) => LMD_OUT(9), B(8) => LMD_OUT(8),
                           B(7) => LMD_OUT(7), B(6) => LMD_OUT(6), B(5) => 
                           LMD_OUT(5), B(4) => LMD_OUT(4), B(3) => LMD_OUT(3), 
                           B(2) => LMD_OUT(2), B(1) => LMD_OUT(1), B(0) => 
                           LMD_OUT(0), S => WB_MUX_SEL, Y(31) => DATAIN_RF(31),
                           Y(30) => DATAIN_RF(30), Y(29) => DATAIN_RF(29), 
                           Y(28) => DATAIN_RF(28), Y(27) => DATAIN_RF(27), 
                           Y(26) => DATAIN_RF(26), Y(25) => DATAIN_RF(25), 
                           Y(24) => DATAIN_RF(24), Y(23) => DATAIN_RF(23), 
                           Y(22) => DATAIN_RF(22), Y(21) => DATAIN_RF(21), 
                           Y(20) => DATAIN_RF(20), Y(19) => DATAIN_RF(19), 
                           Y(18) => DATAIN_RF(18), Y(17) => DATAIN_RF(17), 
                           Y(16) => DATAIN_RF(16), Y(15) => DATAIN_RF(15), 
                           Y(14) => DATAIN_RF(14), Y(13) => DATAIN_RF(13), 
                           Y(12) => DATAIN_RF(12), Y(11) => DATAIN_RF(11), 
                           Y(10) => DATAIN_RF(10), Y(9) => DATAIN_RF(9), Y(8) 
                           => DATAIN_RF(8), Y(7) => DATAIN_RF(7), Y(6) => 
                           DATAIN_RF(6), Y(5) => DATAIN_RF(5), Y(4) => 
                           DATAIN_RF(4), Y(3) => DATAIN_RF(3), Y(2) => 
                           DATAIN_RF(2), Y(1) => DATAIN_RF(1), Y(0) => 
                           DATAIN_RF(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity memoryUnit_nbits32 is

   port( clk, rst, LMD_LATCH_EN, JUMP_EN : in std_logic;  DRAM_DATA, 
         ALUREG_OUTPUT, NPC_OUT : in std_logic_vector (31 downto 0);  COND_OUT 
         : in std_logic;  DRAM_DATAout, TO_PC_OUT, ALU_OUT2 : out 
         std_logic_vector (31 downto 0);  IR_IN4 : in std_logic_vector (31 
         downto 0);  IR_OUT4 : out std_logic_vector (31 downto 0));

end memoryUnit_nbits32;

architecture SYN_STRUCTURAL of memoryUnit_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component register_generic_nbits32_1
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_2
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_bits32_2
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, muxjmp_to_mux, n1, n2 : std_logic;

begin
   DRAM_DATAout <= ( DRAM_DATA(31), DRAM_DATA(30), DRAM_DATA(29), DRAM_DATA(28)
      , DRAM_DATA(27), DRAM_DATA(26), DRAM_DATA(25), DRAM_DATA(24), 
      DRAM_DATA(23), DRAM_DATA(22), DRAM_DATA(21), DRAM_DATA(20), DRAM_DATA(19)
      , DRAM_DATA(18), DRAM_DATA(17), DRAM_DATA(16), DRAM_DATA(15), 
      DRAM_DATA(14), DRAM_DATA(13), DRAM_DATA(12), DRAM_DATA(11), DRAM_DATA(10)
      , DRAM_DATA(9), DRAM_DATA(8), DRAM_DATA(7), DRAM_DATA(6), DRAM_DATA(5), 
      DRAM_DATA(4), DRAM_DATA(3), DRAM_DATA(2), DRAM_DATA(1), DRAM_DATA(0) );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   JUMPMUX : MUX21 port map( A => COND_OUT, B => X_Logic0_port, S => JUMP_EN, Y
                           => muxjmp_to_mux);
   MUX_PC : MUX21_GENERIC_bits32_2 port map( A(31) => ALUREG_OUTPUT(31), A(30) 
                           => ALUREG_OUTPUT(30), A(29) => ALUREG_OUTPUT(29), 
                           A(28) => ALUREG_OUTPUT(28), A(27) => 
                           ALUREG_OUTPUT(27), A(26) => ALUREG_OUTPUT(26), A(25)
                           => ALUREG_OUTPUT(25), A(24) => ALUREG_OUTPUT(24), 
                           A(23) => ALUREG_OUTPUT(23), A(22) => 
                           ALUREG_OUTPUT(22), A(21) => ALUREG_OUTPUT(21), A(20)
                           => ALUREG_OUTPUT(20), A(19) => ALUREG_OUTPUT(19), 
                           A(18) => ALUREG_OUTPUT(18), A(17) => 
                           ALUREG_OUTPUT(17), A(16) => ALUREG_OUTPUT(16), A(15)
                           => ALUREG_OUTPUT(15), A(14) => ALUREG_OUTPUT(14), 
                           A(13) => ALUREG_OUTPUT(13), A(12) => 
                           ALUREG_OUTPUT(12), A(11) => ALUREG_OUTPUT(11), A(10)
                           => ALUREG_OUTPUT(10), A(9) => ALUREG_OUTPUT(9), A(8)
                           => ALUREG_OUTPUT(8), A(7) => ALUREG_OUTPUT(7), A(6) 
                           => ALUREG_OUTPUT(6), A(5) => ALUREG_OUTPUT(5), A(4) 
                           => ALUREG_OUTPUT(4), A(3) => ALUREG_OUTPUT(3), A(2) 
                           => ALUREG_OUTPUT(2), A(1) => ALUREG_OUTPUT(1), A(0) 
                           => ALUREG_OUTPUT(0), B(31) => NPC_OUT(31), B(30) => 
                           NPC_OUT(30), B(29) => NPC_OUT(29), B(28) => 
                           NPC_OUT(28), B(27) => NPC_OUT(27), B(26) => 
                           NPC_OUT(26), B(25) => NPC_OUT(25), B(24) => 
                           NPC_OUT(24), B(23) => NPC_OUT(23), B(22) => 
                           NPC_OUT(22), B(21) => NPC_OUT(21), B(20) => 
                           NPC_OUT(20), B(19) => NPC_OUT(19), B(18) => 
                           NPC_OUT(18), B(17) => NPC_OUT(17), B(16) => 
                           NPC_OUT(16), B(15) => NPC_OUT(15), B(14) => 
                           NPC_OUT(14), B(13) => NPC_OUT(13), B(12) => 
                           NPC_OUT(12), B(11) => NPC_OUT(11), B(10) => 
                           NPC_OUT(10), B(9) => NPC_OUT(9), B(8) => NPC_OUT(8),
                           B(7) => NPC_OUT(7), B(6) => NPC_OUT(6), B(5) => 
                           NPC_OUT(5), B(4) => NPC_OUT(4), B(3) => NPC_OUT(3), 
                           B(2) => NPC_OUT(2), B(1) => NPC_OUT(1), B(0) => 
                           NPC_OUT(0), S => muxjmp_to_mux, Y(31) => 
                           TO_PC_OUT(31), Y(30) => TO_PC_OUT(30), Y(29) => 
                           TO_PC_OUT(29), Y(28) => TO_PC_OUT(28), Y(27) => 
                           TO_PC_OUT(27), Y(26) => TO_PC_OUT(26), Y(25) => 
                           TO_PC_OUT(25), Y(24) => TO_PC_OUT(24), Y(23) => 
                           TO_PC_OUT(23), Y(22) => TO_PC_OUT(22), Y(21) => 
                           TO_PC_OUT(21), Y(20) => TO_PC_OUT(20), Y(19) => 
                           TO_PC_OUT(19), Y(18) => TO_PC_OUT(18), Y(17) => 
                           TO_PC_OUT(17), Y(16) => TO_PC_OUT(16), Y(15) => 
                           TO_PC_OUT(15), Y(14) => TO_PC_OUT(14), Y(13) => 
                           TO_PC_OUT(13), Y(12) => TO_PC_OUT(12), Y(11) => 
                           TO_PC_OUT(11), Y(10) => TO_PC_OUT(10), Y(9) => 
                           TO_PC_OUT(9), Y(8) => TO_PC_OUT(8), Y(7) => 
                           TO_PC_OUT(7), Y(6) => TO_PC_OUT(6), Y(5) => 
                           TO_PC_OUT(5), Y(4) => TO_PC_OUT(4), Y(3) => 
                           TO_PC_OUT(3), Y(2) => TO_PC_OUT(2), Y(1) => 
                           TO_PC_OUT(1), Y(0) => TO_PC_OUT(0));
   ALU_OUT2r : register_generic_nbits32_2 port map( data_in(31) => 
                           ALUREG_OUTPUT(31), data_in(30) => ALUREG_OUTPUT(30),
                           data_in(29) => ALUREG_OUTPUT(29), data_in(28) => 
                           ALUREG_OUTPUT(28), data_in(27) => ALUREG_OUTPUT(27),
                           data_in(26) => ALUREG_OUTPUT(26), data_in(25) => 
                           ALUREG_OUTPUT(25), data_in(24) => ALUREG_OUTPUT(24),
                           data_in(23) => ALUREG_OUTPUT(23), data_in(22) => 
                           ALUREG_OUTPUT(22), data_in(21) => ALUREG_OUTPUT(21),
                           data_in(20) => ALUREG_OUTPUT(20), data_in(19) => 
                           ALUREG_OUTPUT(19), data_in(18) => ALUREG_OUTPUT(18),
                           data_in(17) => ALUREG_OUTPUT(17), data_in(16) => 
                           ALUREG_OUTPUT(16), data_in(15) => ALUREG_OUTPUT(15),
                           data_in(14) => ALUREG_OUTPUT(14), data_in(13) => 
                           ALUREG_OUTPUT(13), data_in(12) => ALUREG_OUTPUT(12),
                           data_in(11) => ALUREG_OUTPUT(11), data_in(10) => 
                           ALUREG_OUTPUT(10), data_in(9) => ALUREG_OUTPUT(9), 
                           data_in(8) => ALUREG_OUTPUT(8), data_in(7) => 
                           ALUREG_OUTPUT(7), data_in(6) => ALUREG_OUTPUT(6), 
                           data_in(5) => ALUREG_OUTPUT(5), data_in(4) => 
                           ALUREG_OUTPUT(4), data_in(3) => ALUREG_OUTPUT(3), 
                           data_in(2) => ALUREG_OUTPUT(2), data_in(1) => 
                           ALUREG_OUTPUT(1), data_in(0) => ALUREG_OUTPUT(0), CK
                           => n2, RESET => n1, ENABLE => X_Logic1_port, 
                           data_out(31) => ALU_OUT2(31), data_out(30) => 
                           ALU_OUT2(30), data_out(29) => ALU_OUT2(29), 
                           data_out(28) => ALU_OUT2(28), data_out(27) => 
                           ALU_OUT2(27), data_out(26) => ALU_OUT2(26), 
                           data_out(25) => ALU_OUT2(25), data_out(24) => 
                           ALU_OUT2(24), data_out(23) => ALU_OUT2(23), 
                           data_out(22) => ALU_OUT2(22), data_out(21) => 
                           ALU_OUT2(21), data_out(20) => ALU_OUT2(20), 
                           data_out(19) => ALU_OUT2(19), data_out(18) => 
                           ALU_OUT2(18), data_out(17) => ALU_OUT2(17), 
                           data_out(16) => ALU_OUT2(16), data_out(15) => 
                           ALU_OUT2(15), data_out(14) => ALU_OUT2(14), 
                           data_out(13) => ALU_OUT2(13), data_out(12) => 
                           ALU_OUT2(12), data_out(11) => ALU_OUT2(11), 
                           data_out(10) => ALU_OUT2(10), data_out(9) => 
                           ALU_OUT2(9), data_out(8) => ALU_OUT2(8), data_out(7)
                           => ALU_OUT2(7), data_out(6) => ALU_OUT2(6), 
                           data_out(5) => ALU_OUT2(5), data_out(4) => 
                           ALU_OUT2(4), data_out(3) => ALU_OUT2(3), data_out(2)
                           => ALU_OUT2(2), data_out(1) => ALU_OUT2(1), 
                           data_out(0) => ALU_OUT2(0));
   IR4 : register_generic_nbits32_1 port map( data_in(31) => IR_IN4(31), 
                           data_in(30) => IR_IN4(30), data_in(29) => IR_IN4(29)
                           , data_in(28) => IR_IN4(28), data_in(27) => 
                           IR_IN4(27), data_in(26) => IR_IN4(26), data_in(25) 
                           => IR_IN4(25), data_in(24) => IR_IN4(24), 
                           data_in(23) => IR_IN4(23), data_in(22) => IR_IN4(22)
                           , data_in(21) => IR_IN4(21), data_in(20) => 
                           IR_IN4(20), data_in(19) => IR_IN4(19), data_in(18) 
                           => IR_IN4(18), data_in(17) => IR_IN4(17), 
                           data_in(16) => IR_IN4(16), data_in(15) => IR_IN4(15)
                           , data_in(14) => IR_IN4(14), data_in(13) => 
                           IR_IN4(13), data_in(12) => IR_IN4(12), data_in(11) 
                           => IR_IN4(11), data_in(10) => IR_IN4(10), data_in(9)
                           => IR_IN4(9), data_in(8) => IR_IN4(8), data_in(7) =>
                           IR_IN4(7), data_in(6) => IR_IN4(6), data_in(5) => 
                           IR_IN4(5), data_in(4) => IR_IN4(4), data_in(3) => 
                           IR_IN4(3), data_in(2) => IR_IN4(2), data_in(1) => 
                           IR_IN4(1), data_in(0) => IR_IN4(0), CK => n2, RESET 
                           => n1, ENABLE => X_Logic1_port, data_out(31) => 
                           IR_OUT4(31), data_out(30) => IR_OUT4(30), 
                           data_out(29) => IR_OUT4(29), data_out(28) => 
                           IR_OUT4(28), data_out(27) => IR_OUT4(27), 
                           data_out(26) => IR_OUT4(26), data_out(25) => 
                           IR_OUT4(25), data_out(24) => IR_OUT4(24), 
                           data_out(23) => IR_OUT4(23), data_out(22) => 
                           IR_OUT4(22), data_out(21) => IR_OUT4(21), 
                           data_out(20) => IR_OUT4(20), data_out(19) => 
                           IR_OUT4(19), data_out(18) => IR_OUT4(18), 
                           data_out(17) => IR_OUT4(17), data_out(16) => 
                           IR_OUT4(16), data_out(15) => IR_OUT4(15), 
                           data_out(14) => IR_OUT4(14), data_out(13) => 
                           IR_OUT4(13), data_out(12) => IR_OUT4(12), 
                           data_out(11) => IR_OUT4(11), data_out(10) => 
                           IR_OUT4(10), data_out(9) => IR_OUT4(9), data_out(8) 
                           => IR_OUT4(8), data_out(7) => IR_OUT4(7), 
                           data_out(6) => IR_OUT4(6), data_out(5) => IR_OUT4(5)
                           , data_out(4) => IR_OUT4(4), data_out(3) => 
                           IR_OUT4(3), data_out(2) => IR_OUT4(2), data_out(1) 
                           => IR_OUT4(1), data_out(0) => IR_OUT4(0));
   U3 : BUF_X1 port map( A => rst, Z => n1);
   U4 : BUF_X1 port map( A => clk, Z => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity executionUnit_nbits32 is

   port( clk, rst, ALU_OUTREG_ENABLE, MUXA_SEL, MUXB_SEL, COND_ENABLE : in 
         std_logic;  ALU_BITS : in std_logic_vector (0 to 3);  NPC_OUT, A_out, 
         B_out, Imm_out : in std_logic_vector (31 downto 0);  ALUREG_OUTPUT : 
         out std_logic_vector (31 downto 0);  COND_OUT : out std_logic;  IR_IN3
         : in std_logic_vector (31 downto 0);  IR_OUT3, B_outreg : out 
         std_logic_vector (31 downto 0));

end executionUnit_nbits32;

architecture SYN_STRUCTURAL of executionUnit_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_0
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component XNOR_logic
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component alu_nbits32
      port( FUNC : in std_logic_vector (0 to 3);  A, B : in std_logic_vector 
            (31 downto 0);  OUTALU : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_3
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_4
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_5
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_bits32_3
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_bits32_0
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component ZERO_DEC_bits32
      port( data : in std_logic_vector (31 downto 0);  zero_detect : out 
            std_logic);
   end component;
   
   signal X_Logic1_port, ZERO_DEC_OUT, MUX1_OUT_31_port, MUX1_OUT_30_port, 
      MUX1_OUT_29_port, MUX1_OUT_28_port, MUX1_OUT_27_port, MUX1_OUT_26_port, 
      MUX1_OUT_25_port, MUX1_OUT_24_port, MUX1_OUT_23_port, MUX1_OUT_22_port, 
      MUX1_OUT_21_port, MUX1_OUT_20_port, MUX1_OUT_19_port, MUX1_OUT_18_port, 
      MUX1_OUT_17_port, MUX1_OUT_16_port, MUX1_OUT_15_port, MUX1_OUT_14_port, 
      MUX1_OUT_13_port, MUX1_OUT_12_port, MUX1_OUT_11_port, MUX1_OUT_10_port, 
      MUX1_OUT_9_port, MUX1_OUT_8_port, MUX1_OUT_7_port, MUX1_OUT_6_port, 
      MUX1_OUT_5_port, MUX1_OUT_4_port, MUX1_OUT_3_port, MUX1_OUT_2_port, 
      MUX1_OUT_1_port, MUX1_OUT_0_port, MUX2_OUT_31_port, MUX2_OUT_30_port, 
      MUX2_OUT_29_port, MUX2_OUT_28_port, MUX2_OUT_27_port, MUX2_OUT_26_port, 
      MUX2_OUT_25_port, MUX2_OUT_24_port, MUX2_OUT_23_port, MUX2_OUT_22_port, 
      MUX2_OUT_21_port, MUX2_OUT_20_port, MUX2_OUT_19_port, MUX2_OUT_18_port, 
      MUX2_OUT_17_port, MUX2_OUT_16_port, MUX2_OUT_15_port, MUX2_OUT_14_port, 
      MUX2_OUT_13_port, MUX2_OUT_12_port, MUX2_OUT_11_port, MUX2_OUT_10_port, 
      MUX2_OUT_9_port, MUX2_OUT_8_port, MUX2_OUT_7_port, MUX2_OUT_6_port, 
      MUX2_OUT_5_port, MUX2_OUT_4_port, MUX2_OUT_3_port, MUX2_OUT_2_port, 
      MUX2_OUT_1_port, MUX2_OUT_0_port, ALU_output_31_port, ALU_output_30_port,
      ALU_output_29_port, ALU_output_28_port, ALU_output_27_port, 
      ALU_output_26_port, ALU_output_25_port, ALU_output_24_port, 
      ALU_output_23_port, ALU_output_22_port, ALU_output_21_port, 
      ALU_output_20_port, ALU_output_19_port, ALU_output_18_port, 
      ALU_output_17_port, ALU_output_16_port, ALU_output_15_port, 
      ALU_output_14_port, ALU_output_13_port, ALU_output_12_port, 
      ALU_output_11_port, ALU_output_10_port, ALU_output_9_port, 
      ALU_output_8_port, ALU_output_7_port, ALU_output_6_port, 
      ALU_output_5_port, ALU_output_4_port, ALU_output_3_port, 
      ALU_output_2_port, ALU_output_1_port, ALU_output_0_port, XNOR_OUT, n1, n2
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   zerodec : ZERO_DEC_bits32 port map( data(31) => A_out(31), data(30) => 
                           A_out(30), data(29) => A_out(29), data(28) => 
                           A_out(28), data(27) => A_out(27), data(26) => 
                           A_out(26), data(25) => A_out(25), data(24) => 
                           A_out(24), data(23) => A_out(23), data(22) => 
                           A_out(22), data(21) => A_out(21), data(20) => 
                           A_out(20), data(19) => A_out(19), data(18) => 
                           A_out(18), data(17) => A_out(17), data(16) => 
                           A_out(16), data(15) => A_out(15), data(14) => 
                           A_out(14), data(13) => A_out(13), data(12) => 
                           A_out(12), data(11) => A_out(11), data(10) => 
                           A_out(10), data(9) => A_out(9), data(8) => A_out(8),
                           data(7) => A_out(7), data(6) => A_out(6), data(5) =>
                           A_out(5), data(4) => A_out(4), data(3) => A_out(3), 
                           data(2) => A_out(2), data(1) => A_out(1), data(0) =>
                           A_out(0), zero_detect => ZERO_DEC_OUT);
   mux1 : MUX21_GENERIC_bits32_0 port map( A(31) => A_out(31), A(30) => 
                           A_out(30), A(29) => A_out(29), A(28) => A_out(28), 
                           A(27) => A_out(27), A(26) => A_out(26), A(25) => 
                           A_out(25), A(24) => A_out(24), A(23) => A_out(23), 
                           A(22) => A_out(22), A(21) => A_out(21), A(20) => 
                           A_out(20), A(19) => A_out(19), A(18) => A_out(18), 
                           A(17) => A_out(17), A(16) => A_out(16), A(15) => 
                           A_out(15), A(14) => A_out(14), A(13) => A_out(13), 
                           A(12) => A_out(12), A(11) => A_out(11), A(10) => 
                           A_out(10), A(9) => A_out(9), A(8) => A_out(8), A(7) 
                           => A_out(7), A(6) => A_out(6), A(5) => A_out(5), 
                           A(4) => A_out(4), A(3) => A_out(3), A(2) => A_out(2)
                           , A(1) => A_out(1), A(0) => A_out(0), B(31) => 
                           NPC_OUT(31), B(30) => NPC_OUT(30), B(29) => 
                           NPC_OUT(29), B(28) => NPC_OUT(28), B(27) => 
                           NPC_OUT(27), B(26) => NPC_OUT(26), B(25) => 
                           NPC_OUT(25), B(24) => NPC_OUT(24), B(23) => 
                           NPC_OUT(23), B(22) => NPC_OUT(22), B(21) => 
                           NPC_OUT(21), B(20) => NPC_OUT(20), B(19) => 
                           NPC_OUT(19), B(18) => NPC_OUT(18), B(17) => 
                           NPC_OUT(17), B(16) => NPC_OUT(16), B(15) => 
                           NPC_OUT(15), B(14) => NPC_OUT(14), B(13) => 
                           NPC_OUT(13), B(12) => NPC_OUT(12), B(11) => 
                           NPC_OUT(11), B(10) => NPC_OUT(10), B(9) => 
                           NPC_OUT(9), B(8) => NPC_OUT(8), B(7) => NPC_OUT(7), 
                           B(6) => NPC_OUT(6), B(5) => NPC_OUT(5), B(4) => 
                           NPC_OUT(4), B(3) => NPC_OUT(3), B(2) => NPC_OUT(2), 
                           B(1) => NPC_OUT(1), B(0) => NPC_OUT(0), S => 
                           MUXA_SEL, Y(31) => MUX1_OUT_31_port, Y(30) => 
                           MUX1_OUT_30_port, Y(29) => MUX1_OUT_29_port, Y(28) 
                           => MUX1_OUT_28_port, Y(27) => MUX1_OUT_27_port, 
                           Y(26) => MUX1_OUT_26_port, Y(25) => MUX1_OUT_25_port
                           , Y(24) => MUX1_OUT_24_port, Y(23) => 
                           MUX1_OUT_23_port, Y(22) => MUX1_OUT_22_port, Y(21) 
                           => MUX1_OUT_21_port, Y(20) => MUX1_OUT_20_port, 
                           Y(19) => MUX1_OUT_19_port, Y(18) => MUX1_OUT_18_port
                           , Y(17) => MUX1_OUT_17_port, Y(16) => 
                           MUX1_OUT_16_port, Y(15) => MUX1_OUT_15_port, Y(14) 
                           => MUX1_OUT_14_port, Y(13) => MUX1_OUT_13_port, 
                           Y(12) => MUX1_OUT_12_port, Y(11) => MUX1_OUT_11_port
                           , Y(10) => MUX1_OUT_10_port, Y(9) => MUX1_OUT_9_port
                           , Y(8) => MUX1_OUT_8_port, Y(7) => MUX1_OUT_7_port, 
                           Y(6) => MUX1_OUT_6_port, Y(5) => MUX1_OUT_5_port, 
                           Y(4) => MUX1_OUT_4_port, Y(3) => MUX1_OUT_3_port, 
                           Y(2) => MUX1_OUT_2_port, Y(1) => MUX1_OUT_1_port, 
                           Y(0) => MUX1_OUT_0_port);
   mux2 : MUX21_GENERIC_bits32_3 port map( A(31) => Imm_out(31), A(30) => 
                           Imm_out(30), A(29) => Imm_out(29), A(28) => 
                           Imm_out(28), A(27) => Imm_out(27), A(26) => 
                           Imm_out(26), A(25) => Imm_out(25), A(24) => 
                           Imm_out(24), A(23) => Imm_out(23), A(22) => 
                           Imm_out(22), A(21) => Imm_out(21), A(20) => 
                           Imm_out(20), A(19) => Imm_out(19), A(18) => 
                           Imm_out(18), A(17) => Imm_out(17), A(16) => 
                           Imm_out(16), A(15) => Imm_out(15), A(14) => 
                           Imm_out(14), A(13) => Imm_out(13), A(12) => 
                           Imm_out(12), A(11) => Imm_out(11), A(10) => 
                           Imm_out(10), A(9) => Imm_out(9), A(8) => Imm_out(8),
                           A(7) => Imm_out(7), A(6) => Imm_out(6), A(5) => 
                           Imm_out(5), A(4) => Imm_out(4), A(3) => Imm_out(3), 
                           A(2) => Imm_out(2), A(1) => Imm_out(1), A(0) => 
                           Imm_out(0), B(31) => B_out(31), B(30) => B_out(30), 
                           B(29) => B_out(29), B(28) => B_out(28), B(27) => 
                           B_out(27), B(26) => B_out(26), B(25) => B_out(25), 
                           B(24) => B_out(24), B(23) => B_out(23), B(22) => 
                           B_out(22), B(21) => B_out(21), B(20) => B_out(20), 
                           B(19) => B_out(19), B(18) => B_out(18), B(17) => 
                           B_out(17), B(16) => B_out(16), B(15) => B_out(15), 
                           B(14) => B_out(14), B(13) => B_out(13), B(12) => 
                           B_out(12), B(11) => B_out(11), B(10) => B_out(10), 
                           B(9) => B_out(9), B(8) => B_out(8), B(7) => B_out(7)
                           , B(6) => B_out(6), B(5) => B_out(5), B(4) => 
                           B_out(4), B(3) => B_out(3), B(2) => B_out(2), B(1) 
                           => B_out(1), B(0) => B_out(0), S => MUXB_SEL, Y(31) 
                           => MUX2_OUT_31_port, Y(30) => MUX2_OUT_30_port, 
                           Y(29) => MUX2_OUT_29_port, Y(28) => MUX2_OUT_28_port
                           , Y(27) => MUX2_OUT_27_port, Y(26) => 
                           MUX2_OUT_26_port, Y(25) => MUX2_OUT_25_port, Y(24) 
                           => MUX2_OUT_24_port, Y(23) => MUX2_OUT_23_port, 
                           Y(22) => MUX2_OUT_22_port, Y(21) => MUX2_OUT_21_port
                           , Y(20) => MUX2_OUT_20_port, Y(19) => 
                           MUX2_OUT_19_port, Y(18) => MUX2_OUT_18_port, Y(17) 
                           => MUX2_OUT_17_port, Y(16) => MUX2_OUT_16_port, 
                           Y(15) => MUX2_OUT_15_port, Y(14) => MUX2_OUT_14_port
                           , Y(13) => MUX2_OUT_13_port, Y(12) => 
                           MUX2_OUT_12_port, Y(11) => MUX2_OUT_11_port, Y(10) 
                           => MUX2_OUT_10_port, Y(9) => MUX2_OUT_9_port, Y(8) 
                           => MUX2_OUT_8_port, Y(7) => MUX2_OUT_7_port, Y(6) =>
                           MUX2_OUT_6_port, Y(5) => MUX2_OUT_5_port, Y(4) => 
                           MUX2_OUT_4_port, Y(3) => MUX2_OUT_3_port, Y(2) => 
                           MUX2_OUT_2_port, Y(1) => MUX2_OUT_1_port, Y(0) => 
                           MUX2_OUT_0_port);
   ALUoutput : register_generic_nbits32_5 port map( data_in(31) => 
                           ALU_output_31_port, data_in(30) => 
                           ALU_output_30_port, data_in(29) => 
                           ALU_output_29_port, data_in(28) => 
                           ALU_output_28_port, data_in(27) => 
                           ALU_output_27_port, data_in(26) => 
                           ALU_output_26_port, data_in(25) => 
                           ALU_output_25_port, data_in(24) => 
                           ALU_output_24_port, data_in(23) => 
                           ALU_output_23_port, data_in(22) => 
                           ALU_output_22_port, data_in(21) => 
                           ALU_output_21_port, data_in(20) => 
                           ALU_output_20_port, data_in(19) => 
                           ALU_output_19_port, data_in(18) => 
                           ALU_output_18_port, data_in(17) => 
                           ALU_output_17_port, data_in(16) => 
                           ALU_output_16_port, data_in(15) => 
                           ALU_output_15_port, data_in(14) => 
                           ALU_output_14_port, data_in(13) => 
                           ALU_output_13_port, data_in(12) => 
                           ALU_output_12_port, data_in(11) => 
                           ALU_output_11_port, data_in(10) => 
                           ALU_output_10_port, data_in(9) => ALU_output_9_port,
                           data_in(8) => ALU_output_8_port, data_in(7) => 
                           ALU_output_7_port, data_in(6) => ALU_output_6_port, 
                           data_in(5) => ALU_output_5_port, data_in(4) => 
                           ALU_output_4_port, data_in(3) => ALU_output_3_port, 
                           data_in(2) => ALU_output_2_port, data_in(1) => 
                           ALU_output_1_port, data_in(0) => ALU_output_0_port, 
                           CK => n2, RESET => n1, ENABLE => ALU_OUTREG_ENABLE, 
                           data_out(31) => ALUREG_OUTPUT(31), data_out(30) => 
                           ALUREG_OUTPUT(30), data_out(29) => ALUREG_OUTPUT(29)
                           , data_out(28) => ALUREG_OUTPUT(28), data_out(27) =>
                           ALUREG_OUTPUT(27), data_out(26) => ALUREG_OUTPUT(26)
                           , data_out(25) => ALUREG_OUTPUT(25), data_out(24) =>
                           ALUREG_OUTPUT(24), data_out(23) => ALUREG_OUTPUT(23)
                           , data_out(22) => ALUREG_OUTPUT(22), data_out(21) =>
                           ALUREG_OUTPUT(21), data_out(20) => ALUREG_OUTPUT(20)
                           , data_out(19) => ALUREG_OUTPUT(19), data_out(18) =>
                           ALUREG_OUTPUT(18), data_out(17) => ALUREG_OUTPUT(17)
                           , data_out(16) => ALUREG_OUTPUT(16), data_out(15) =>
                           ALUREG_OUTPUT(15), data_out(14) => ALUREG_OUTPUT(14)
                           , data_out(13) => ALUREG_OUTPUT(13), data_out(12) =>
                           ALUREG_OUTPUT(12), data_out(11) => ALUREG_OUTPUT(11)
                           , data_out(10) => ALUREG_OUTPUT(10), data_out(9) => 
                           ALUREG_OUTPUT(9), data_out(8) => ALUREG_OUTPUT(8), 
                           data_out(7) => ALUREG_OUTPUT(7), data_out(6) => 
                           ALUREG_OUTPUT(6), data_out(5) => ALUREG_OUTPUT(5), 
                           data_out(4) => ALUREG_OUTPUT(4), data_out(3) => 
                           ALUREG_OUTPUT(3), data_out(2) => ALUREG_OUTPUT(2), 
                           data_out(1) => ALUREG_OUTPUT(1), data_out(0) => 
                           ALUREG_OUTPUT(0));
   IR3 : register_generic_nbits32_4 port map( data_in(31) => IR_IN3(31), 
                           data_in(30) => IR_IN3(30), data_in(29) => IR_IN3(29)
                           , data_in(28) => IR_IN3(28), data_in(27) => 
                           IR_IN3(27), data_in(26) => IR_IN3(26), data_in(25) 
                           => IR_IN3(25), data_in(24) => IR_IN3(24), 
                           data_in(23) => IR_IN3(23), data_in(22) => IR_IN3(22)
                           , data_in(21) => IR_IN3(21), data_in(20) => 
                           IR_IN3(20), data_in(19) => IR_IN3(19), data_in(18) 
                           => IR_IN3(18), data_in(17) => IR_IN3(17), 
                           data_in(16) => IR_IN3(16), data_in(15) => IR_IN3(15)
                           , data_in(14) => IR_IN3(14), data_in(13) => 
                           IR_IN3(13), data_in(12) => IR_IN3(12), data_in(11) 
                           => IR_IN3(11), data_in(10) => IR_IN3(10), data_in(9)
                           => IR_IN3(9), data_in(8) => IR_IN3(8), data_in(7) =>
                           IR_IN3(7), data_in(6) => IR_IN3(6), data_in(5) => 
                           IR_IN3(5), data_in(4) => IR_IN3(4), data_in(3) => 
                           IR_IN3(3), data_in(2) => IR_IN3(2), data_in(1) => 
                           IR_IN3(1), data_in(0) => IR_IN3(0), CK => n2, RESET 
                           => n1, ENABLE => X_Logic1_port, data_out(31) => 
                           IR_OUT3(31), data_out(30) => IR_OUT3(30), 
                           data_out(29) => IR_OUT3(29), data_out(28) => 
                           IR_OUT3(28), data_out(27) => IR_OUT3(27), 
                           data_out(26) => IR_OUT3(26), data_out(25) => 
                           IR_OUT3(25), data_out(24) => IR_OUT3(24), 
                           data_out(23) => IR_OUT3(23), data_out(22) => 
                           IR_OUT3(22), data_out(21) => IR_OUT3(21), 
                           data_out(20) => IR_OUT3(20), data_out(19) => 
                           IR_OUT3(19), data_out(18) => IR_OUT3(18), 
                           data_out(17) => IR_OUT3(17), data_out(16) => 
                           IR_OUT3(16), data_out(15) => IR_OUT3(15), 
                           data_out(14) => IR_OUT3(14), data_out(13) => 
                           IR_OUT3(13), data_out(12) => IR_OUT3(12), 
                           data_out(11) => IR_OUT3(11), data_out(10) => 
                           IR_OUT3(10), data_out(9) => IR_OUT3(9), data_out(8) 
                           => IR_OUT3(8), data_out(7) => IR_OUT3(7), 
                           data_out(6) => IR_OUT3(6), data_out(5) => IR_OUT3(5)
                           , data_out(4) => IR_OUT3(4), data_out(3) => 
                           IR_OUT3(3), data_out(2) => IR_OUT3(2), data_out(1) 
                           => IR_OUT3(1), data_out(0) => IR_OUT3(0));
   B_outregister : register_generic_nbits32_3 port map( data_in(31) => 
                           B_out(31), data_in(30) => B_out(30), data_in(29) => 
                           B_out(29), data_in(28) => B_out(28), data_in(27) => 
                           B_out(27), data_in(26) => B_out(26), data_in(25) => 
                           B_out(25), data_in(24) => B_out(24), data_in(23) => 
                           B_out(23), data_in(22) => B_out(22), data_in(21) => 
                           B_out(21), data_in(20) => B_out(20), data_in(19) => 
                           B_out(19), data_in(18) => B_out(18), data_in(17) => 
                           B_out(17), data_in(16) => B_out(16), data_in(15) => 
                           B_out(15), data_in(14) => B_out(14), data_in(13) => 
                           B_out(13), data_in(12) => B_out(12), data_in(11) => 
                           B_out(11), data_in(10) => B_out(10), data_in(9) => 
                           B_out(9), data_in(8) => B_out(8), data_in(7) => 
                           B_out(7), data_in(6) => B_out(6), data_in(5) => 
                           B_out(5), data_in(4) => B_out(4), data_in(3) => 
                           B_out(3), data_in(2) => B_out(2), data_in(1) => 
                           B_out(1), data_in(0) => B_out(0), CK => n2, RESET =>
                           n1, ENABLE => X_Logic1_port, data_out(31) => 
                           B_outreg(31), data_out(30) => B_outreg(30), 
                           data_out(29) => B_outreg(29), data_out(28) => 
                           B_outreg(28), data_out(27) => B_outreg(27), 
                           data_out(26) => B_outreg(26), data_out(25) => 
                           B_outreg(25), data_out(24) => B_outreg(24), 
                           data_out(23) => B_outreg(23), data_out(22) => 
                           B_outreg(22), data_out(21) => B_outreg(21), 
                           data_out(20) => B_outreg(20), data_out(19) => 
                           B_outreg(19), data_out(18) => B_outreg(18), 
                           data_out(17) => B_outreg(17), data_out(16) => 
                           B_outreg(16), data_out(15) => B_outreg(15), 
                           data_out(14) => B_outreg(14), data_out(13) => 
                           B_outreg(13), data_out(12) => B_outreg(12), 
                           data_out(11) => B_outreg(11), data_out(10) => 
                           B_outreg(10), data_out(9) => B_outreg(9), 
                           data_out(8) => B_outreg(8), data_out(7) => 
                           B_outreg(7), data_out(6) => B_outreg(6), data_out(5)
                           => B_outreg(5), data_out(4) => B_outreg(4), 
                           data_out(3) => B_outreg(3), data_out(2) => 
                           B_outreg(2), data_out(1) => B_outreg(1), data_out(0)
                           => B_outreg(0));
   alu1 : alu_nbits32 port map( FUNC(0) => ALU_BITS(0), FUNC(1) => ALU_BITS(1),
                           FUNC(2) => ALU_BITS(2), FUNC(3) => ALU_BITS(3), 
                           A(31) => MUX1_OUT_31_port, A(30) => MUX1_OUT_30_port
                           , A(29) => MUX1_OUT_29_port, A(28) => 
                           MUX1_OUT_28_port, A(27) => MUX1_OUT_27_port, A(26) 
                           => MUX1_OUT_26_port, A(25) => MUX1_OUT_25_port, 
                           A(24) => MUX1_OUT_24_port, A(23) => MUX1_OUT_23_port
                           , A(22) => MUX1_OUT_22_port, A(21) => 
                           MUX1_OUT_21_port, A(20) => MUX1_OUT_20_port, A(19) 
                           => MUX1_OUT_19_port, A(18) => MUX1_OUT_18_port, 
                           A(17) => MUX1_OUT_17_port, A(16) => MUX1_OUT_16_port
                           , A(15) => MUX1_OUT_15_port, A(14) => 
                           MUX1_OUT_14_port, A(13) => MUX1_OUT_13_port, A(12) 
                           => MUX1_OUT_12_port, A(11) => MUX1_OUT_11_port, 
                           A(10) => MUX1_OUT_10_port, A(9) => MUX1_OUT_9_port, 
                           A(8) => MUX1_OUT_8_port, A(7) => MUX1_OUT_7_port, 
                           A(6) => MUX1_OUT_6_port, A(5) => MUX1_OUT_5_port, 
                           A(4) => MUX1_OUT_4_port, A(3) => MUX1_OUT_3_port, 
                           A(2) => MUX1_OUT_2_port, A(1) => MUX1_OUT_1_port, 
                           A(0) => MUX1_OUT_0_port, B(31) => MUX2_OUT_31_port, 
                           B(30) => MUX2_OUT_30_port, B(29) => MUX2_OUT_29_port
                           , B(28) => MUX2_OUT_28_port, B(27) => 
                           MUX2_OUT_27_port, B(26) => MUX2_OUT_26_port, B(25) 
                           => MUX2_OUT_25_port, B(24) => MUX2_OUT_24_port, 
                           B(23) => MUX2_OUT_23_port, B(22) => MUX2_OUT_22_port
                           , B(21) => MUX2_OUT_21_port, B(20) => 
                           MUX2_OUT_20_port, B(19) => MUX2_OUT_19_port, B(18) 
                           => MUX2_OUT_18_port, B(17) => MUX2_OUT_17_port, 
                           B(16) => MUX2_OUT_16_port, B(15) => MUX2_OUT_15_port
                           , B(14) => MUX2_OUT_14_port, B(13) => 
                           MUX2_OUT_13_port, B(12) => MUX2_OUT_12_port, B(11) 
                           => MUX2_OUT_11_port, B(10) => MUX2_OUT_10_port, B(9)
                           => MUX2_OUT_9_port, B(8) => MUX2_OUT_8_port, B(7) =>
                           MUX2_OUT_7_port, B(6) => MUX2_OUT_6_port, B(5) => 
                           MUX2_OUT_5_port, B(4) => MUX2_OUT_4_port, B(3) => 
                           MUX2_OUT_3_port, B(2) => MUX2_OUT_2_port, B(1) => 
                           MUX2_OUT_1_port, B(0) => MUX2_OUT_0_port, OUTALU(31)
                           => ALU_output_31_port, OUTALU(30) => 
                           ALU_output_30_port, OUTALU(29) => ALU_output_29_port
                           , OUTALU(28) => ALU_output_28_port, OUTALU(27) => 
                           ALU_output_27_port, OUTALU(26) => ALU_output_26_port
                           , OUTALU(25) => ALU_output_25_port, OUTALU(24) => 
                           ALU_output_24_port, OUTALU(23) => ALU_output_23_port
                           , OUTALU(22) => ALU_output_22_port, OUTALU(21) => 
                           ALU_output_21_port, OUTALU(20) => ALU_output_20_port
                           , OUTALU(19) => ALU_output_19_port, OUTALU(18) => 
                           ALU_output_18_port, OUTALU(17) => ALU_output_17_port
                           , OUTALU(16) => ALU_output_16_port, OUTALU(15) => 
                           ALU_output_15_port, OUTALU(14) => ALU_output_14_port
                           , OUTALU(13) => ALU_output_13_port, OUTALU(12) => 
                           ALU_output_12_port, OUTALU(11) => ALU_output_11_port
                           , OUTALU(10) => ALU_output_10_port, OUTALU(9) => 
                           ALU_output_9_port, OUTALU(8) => ALU_output_8_port, 
                           OUTALU(7) => ALU_output_7_port, OUTALU(6) => 
                           ALU_output_6_port, OUTALU(5) => ALU_output_5_port, 
                           OUTALU(4) => ALU_output_4_port, OUTALU(3) => 
                           ALU_output_3_port, OUTALU(2) => ALU_output_2_port, 
                           OUTALU(1) => ALU_output_1_port, OUTALU(0) => 
                           ALU_output_0_port);
   XNOR_2 : XNOR_logic port map( A => ZERO_DEC_OUT, B => COND_ENABLE, Y => 
                           XNOR_OUT);
   COND : FD_0 port map( D => XNOR_OUT, CK => n2, RESET => n1, ENABLE => 
                           X_Logic1_port, Q => COND_OUT);
   U2 : BUF_X1 port map( A => rst, Z => n1);
   U3 : BUF_X1 port map( A => clk, Z => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity decodeUnit_nbits32 is

   port( clk, rst, RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE : in 
         std_logic;  DATAIN, IR_OUT : in std_logic_vector (31 downto 0);  A_out
         , B_out, Imm_out : out std_logic_vector (31 downto 0);  IR_IN2 : in 
         std_logic_vector (31 downto 0);  IR_OUT2 : out std_logic_vector (31 
         downto 0);  NPC_IN : in std_logic_vector (31 downto 0);  NPC2_OUT : 
         out std_logic_vector (31 downto 0));

end decodeUnit_nbits32;

architecture SYN_STRUCTURAL of decodeUnit_nbits32 is

   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component REGISTER_FILE_NBITS32_NREGISTERS32
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component SIGN_EXT_bits16
      port( inputt : in std_logic_vector (15 downto 0);  outputt : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_6
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_7
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_8
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, signExtOut_31_port, signExtOut_30_port, 
      signExtOut_29_port, signExtOut_28_port, signExtOut_27_port, 
      signExtOut_26_port, signExtOut_25_port, signExtOut_24_port, 
      signExtOut_23_port, signExtOut_22_port, signExtOut_21_port, 
      signExtOut_20_port, signExtOut_19_port, signExtOut_18_port, 
      signExtOut_17_port, signExtOut_16_port, signExtOut_15_port, 
      signExtOut_14_port, signExtOut_13_port, signExtOut_12_port, 
      signExtOut_11_port, signExtOut_10_port, signExtOut_9_port, 
      signExtOut_8_port, signExtOut_7_port, signExtOut_6_port, 
      signExtOut_5_port, signExtOut_4_port, signExtOut_3_port, 
      signExtOut_2_port, signExtOut_1_port, signExtOut_0_port, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9 : std_logic;

begin
   
   X_Logic1_port <= '1';
   NPC2 : register_generic_nbits32_8 port map( data_in(31) => NPC_IN(31), 
                           data_in(30) => NPC_IN(30), data_in(29) => NPC_IN(29)
                           , data_in(28) => NPC_IN(28), data_in(27) => 
                           NPC_IN(27), data_in(26) => NPC_IN(26), data_in(25) 
                           => NPC_IN(25), data_in(24) => NPC_IN(24), 
                           data_in(23) => NPC_IN(23), data_in(22) => NPC_IN(22)
                           , data_in(21) => NPC_IN(21), data_in(20) => 
                           NPC_IN(20), data_in(19) => NPC_IN(19), data_in(18) 
                           => NPC_IN(18), data_in(17) => NPC_IN(17), 
                           data_in(16) => NPC_IN(16), data_in(15) => NPC_IN(15)
                           , data_in(14) => NPC_IN(14), data_in(13) => 
                           NPC_IN(13), data_in(12) => NPC_IN(12), data_in(11) 
                           => NPC_IN(11), data_in(10) => NPC_IN(10), data_in(9)
                           => NPC_IN(9), data_in(8) => NPC_IN(8), data_in(7) =>
                           NPC_IN(7), data_in(6) => NPC_IN(6), data_in(5) => 
                           NPC_IN(5), data_in(4) => NPC_IN(4), data_in(3) => 
                           NPC_IN(3), data_in(2) => NPC_IN(2), data_in(1) => 
                           NPC_IN(1), data_in(0) => NPC_IN(0), CK => n2, RESET 
                           => n1, ENABLE => X_Logic1_port, data_out(31) => 
                           NPC2_OUT(31), data_out(30) => NPC2_OUT(30), 
                           data_out(29) => NPC2_OUT(29), data_out(28) => 
                           NPC2_OUT(28), data_out(27) => NPC2_OUT(27), 
                           data_out(26) => NPC2_OUT(26), data_out(25) => 
                           NPC2_OUT(25), data_out(24) => NPC2_OUT(24), 
                           data_out(23) => NPC2_OUT(23), data_out(22) => 
                           NPC2_OUT(22), data_out(21) => NPC2_OUT(21), 
                           data_out(20) => NPC2_OUT(20), data_out(19) => 
                           NPC2_OUT(19), data_out(18) => NPC2_OUT(18), 
                           data_out(17) => NPC2_OUT(17), data_out(16) => 
                           NPC2_OUT(16), data_out(15) => NPC2_OUT(15), 
                           data_out(14) => NPC2_OUT(14), data_out(13) => 
                           NPC2_OUT(13), data_out(12) => NPC2_OUT(12), 
                           data_out(11) => NPC2_OUT(11), data_out(10) => 
                           NPC2_OUT(10), data_out(9) => NPC2_OUT(9), 
                           data_out(8) => NPC2_OUT(8), data_out(7) => 
                           NPC2_OUT(7), data_out(6) => NPC2_OUT(6), data_out(5)
                           => NPC2_OUT(5), data_out(4) => NPC2_OUT(4), 
                           data_out(3) => NPC2_OUT(3), data_out(2) => 
                           NPC2_OUT(2), data_out(1) => NPC2_OUT(1), data_out(0)
                           => NPC2_OUT(0));
   Imm : register_generic_nbits32_7 port map( data_in(31) => signExtOut_31_port
                           , data_in(30) => signExtOut_30_port, data_in(29) => 
                           signExtOut_29_port, data_in(28) => 
                           signExtOut_28_port, data_in(27) => 
                           signExtOut_27_port, data_in(26) => 
                           signExtOut_26_port, data_in(25) => 
                           signExtOut_25_port, data_in(24) => 
                           signExtOut_24_port, data_in(23) => 
                           signExtOut_23_port, data_in(22) => 
                           signExtOut_22_port, data_in(21) => 
                           signExtOut_21_port, data_in(20) => 
                           signExtOut_20_port, data_in(19) => 
                           signExtOut_19_port, data_in(18) => 
                           signExtOut_18_port, data_in(17) => 
                           signExtOut_17_port, data_in(16) => 
                           signExtOut_16_port, data_in(15) => 
                           signExtOut_15_port, data_in(14) => 
                           signExtOut_14_port, data_in(13) => 
                           signExtOut_13_port, data_in(12) => 
                           signExtOut_12_port, data_in(11) => 
                           signExtOut_11_port, data_in(10) => 
                           signExtOut_10_port, data_in(9) => signExtOut_9_port,
                           data_in(8) => signExtOut_8_port, data_in(7) => 
                           signExtOut_7_port, data_in(6) => signExtOut_6_port, 
                           data_in(5) => signExtOut_5_port, data_in(4) => 
                           signExtOut_4_port, data_in(3) => signExtOut_3_port, 
                           data_in(2) => signExtOut_2_port, data_in(1) => 
                           signExtOut_1_port, data_in(0) => signExtOut_0_port, 
                           CK => n2, RESET => n1, ENABLE => RegIMM_LATCH_EN, 
                           data_out(31) => Imm_out(31), data_out(30) => 
                           Imm_out(30), data_out(29) => Imm_out(29), 
                           data_out(28) => Imm_out(28), data_out(27) => 
                           Imm_out(27), data_out(26) => Imm_out(26), 
                           data_out(25) => Imm_out(25), data_out(24) => 
                           Imm_out(24), data_out(23) => Imm_out(23), 
                           data_out(22) => Imm_out(22), data_out(21) => 
                           Imm_out(21), data_out(20) => Imm_out(20), 
                           data_out(19) => Imm_out(19), data_out(18) => 
                           Imm_out(18), data_out(17) => Imm_out(17), 
                           data_out(16) => Imm_out(16), data_out(15) => 
                           Imm_out(15), data_out(14) => Imm_out(14), 
                           data_out(13) => Imm_out(13), data_out(12) => 
                           Imm_out(12), data_out(11) => Imm_out(11), 
                           data_out(10) => Imm_out(10), data_out(9) => 
                           Imm_out(9), data_out(8) => Imm_out(8), data_out(7) 
                           => Imm_out(7), data_out(6) => Imm_out(6), 
                           data_out(5) => Imm_out(5), data_out(4) => Imm_out(4)
                           , data_out(3) => Imm_out(3), data_out(2) => 
                           Imm_out(2), data_out(1) => Imm_out(1), data_out(0) 
                           => Imm_out(0));
   IR2 : register_generic_nbits32_6 port map( data_in(31) => IR_OUT(31), 
                           data_in(30) => IR_OUT(30), data_in(29) => IR_OUT(29)
                           , data_in(28) => IR_OUT(28), data_in(27) => 
                           IR_OUT(27), data_in(26) => IR_OUT(26), data_in(25) 
                           => IR_OUT(25), data_in(24) => IR_OUT(24), 
                           data_in(23) => IR_OUT(23), data_in(22) => IR_OUT(22)
                           , data_in(21) => IR_OUT(21), data_in(20) => 
                           IR_OUT(20), data_in(19) => IR_OUT(19), data_in(18) 
                           => IR_OUT(18), data_in(17) => IR_OUT(17), 
                           data_in(16) => IR_OUT(16), data_in(15) => IR_OUT(15)
                           , data_in(14) => IR_OUT(14), data_in(13) => 
                           IR_OUT(13), data_in(12) => IR_OUT(12), data_in(11) 
                           => IR_OUT(11), data_in(10) => IR_OUT(10), data_in(9)
                           => IR_OUT(9), data_in(8) => IR_OUT(8), data_in(7) =>
                           IR_OUT(7), data_in(6) => IR_OUT(6), data_in(5) => 
                           IR_OUT(5), data_in(4) => IR_OUT(4), data_in(3) => 
                           IR_OUT(3), data_in(2) => IR_OUT(2), data_in(1) => 
                           IR_OUT(1), data_in(0) => IR_OUT(0), CK => n2, RESET 
                           => n1, ENABLE => X_Logic1_port, data_out(31) => 
                           IR_OUT2(31), data_out(30) => IR_OUT2(30), 
                           data_out(29) => IR_OUT2(29), data_out(28) => 
                           IR_OUT2(28), data_out(27) => IR_OUT2(27), 
                           data_out(26) => IR_OUT2(26), data_out(25) => 
                           IR_OUT2(25), data_out(24) => IR_OUT2(24), 
                           data_out(23) => IR_OUT2(23), data_out(22) => 
                           IR_OUT2(22), data_out(21) => IR_OUT2(21), 
                           data_out(20) => IR_OUT2(20), data_out(19) => 
                           IR_OUT2(19), data_out(18) => IR_OUT2(18), 
                           data_out(17) => IR_OUT2(17), data_out(16) => 
                           IR_OUT2(16), data_out(15) => IR_OUT2(15), 
                           data_out(14) => IR_OUT2(14), data_out(13) => 
                           IR_OUT2(13), data_out(12) => IR_OUT2(12), 
                           data_out(11) => IR_OUT2(11), data_out(10) => 
                           IR_OUT2(10), data_out(9) => IR_OUT2(9), data_out(8) 
                           => IR_OUT2(8), data_out(7) => IR_OUT2(7), 
                           data_out(6) => IR_OUT2(6), data_out(5) => IR_OUT2(5)
                           , data_out(4) => IR_OUT2(4), data_out(3) => 
                           IR_OUT2(3), data_out(2) => IR_OUT2(2), data_out(1) 
                           => IR_OUT2(1), data_out(0) => IR_OUT2(0));
   Signext : SIGN_EXT_bits16 port map( inputt(15) => IR_OUT(15), inputt(14) => 
                           IR_OUT(14), inputt(13) => IR_OUT(13), inputt(12) => 
                           IR_OUT(12), inputt(11) => IR_OUT(11), inputt(10) => 
                           IR_OUT(10), inputt(9) => IR_OUT(9), inputt(8) => 
                           IR_OUT(8), inputt(7) => IR_OUT(7), inputt(6) => 
                           IR_OUT(6), inputt(5) => IR_OUT(5), inputt(4) => 
                           IR_OUT(4), inputt(3) => IR_OUT(3), inputt(2) => 
                           IR_OUT(2), inputt(1) => IR_OUT(1), inputt(0) => 
                           IR_OUT(0), outputt(31) => signExtOut_31_port, 
                           outputt(30) => signExtOut_30_port, outputt(29) => 
                           signExtOut_29_port, outputt(28) => 
                           signExtOut_28_port, outputt(27) => 
                           signExtOut_27_port, outputt(26) => 
                           signExtOut_26_port, outputt(25) => 
                           signExtOut_25_port, outputt(24) => 
                           signExtOut_24_port, outputt(23) => 
                           signExtOut_23_port, outputt(22) => 
                           signExtOut_22_port, outputt(21) => 
                           signExtOut_21_port, outputt(20) => 
                           signExtOut_20_port, outputt(19) => 
                           signExtOut_19_port, outputt(18) => 
                           signExtOut_18_port, outputt(17) => 
                           signExtOut_17_port, outputt(16) => 
                           signExtOut_16_port, outputt(15) => 
                           signExtOut_15_port, outputt(14) => 
                           signExtOut_14_port, outputt(13) => 
                           signExtOut_13_port, outputt(12) => 
                           signExtOut_12_port, outputt(11) => 
                           signExtOut_11_port, outputt(10) => 
                           signExtOut_10_port, outputt(9) => signExtOut_9_port,
                           outputt(8) => signExtOut_8_port, outputt(7) => 
                           signExtOut_7_port, outputt(6) => signExtOut_6_port, 
                           outputt(5) => signExtOut_5_port, outputt(4) => 
                           signExtOut_4_port, outputt(3) => signExtOut_3_port, 
                           outputt(2) => signExtOut_2_port, outputt(1) => 
                           signExtOut_1_port, outputt(0) => signExtOut_0_port);
   RF : REGISTER_FILE_NBITS32_NREGISTERS32 port map( CLK => n2, RESET => n1, 
                           ENABLE => X_Logic1_port, RD1 => X_Logic1_port, RD2 
                           => X_Logic1_port, WR => RF_WE, ADD_WR(4) => n9, 
                           ADD_WR(3) => n8, ADD_WR(2) => n7, ADD_WR(1) => n6, 
                           ADD_WR(0) => n5, ADD_RD1(4) => IR_OUT(25), 
                           ADD_RD1(3) => IR_OUT(24), ADD_RD1(2) => IR_OUT(23), 
                           ADD_RD1(1) => IR_OUT(22), ADD_RD1(0) => IR_OUT(21), 
                           ADD_RD2(4) => IR_OUT(20), ADD_RD2(3) => IR_OUT(19), 
                           ADD_RD2(2) => IR_OUT(18), ADD_RD2(1) => IR_OUT(17), 
                           ADD_RD2(0) => IR_OUT(16), DATAIN(31) => DATAIN(31), 
                           DATAIN(30) => DATAIN(30), DATAIN(29) => DATAIN(29), 
                           DATAIN(28) => DATAIN(28), DATAIN(27) => DATAIN(27), 
                           DATAIN(26) => DATAIN(26), DATAIN(25) => DATAIN(25), 
                           DATAIN(24) => DATAIN(24), DATAIN(23) => DATAIN(23), 
                           DATAIN(22) => DATAIN(22), DATAIN(21) => DATAIN(21), 
                           DATAIN(20) => DATAIN(20), DATAIN(19) => DATAIN(19), 
                           DATAIN(18) => DATAIN(18), DATAIN(17) => DATAIN(17), 
                           DATAIN(16) => DATAIN(16), DATAIN(15) => DATAIN(15), 
                           DATAIN(14) => DATAIN(14), DATAIN(13) => DATAIN(13), 
                           DATAIN(12) => DATAIN(12), DATAIN(11) => DATAIN(11), 
                           DATAIN(10) => DATAIN(10), DATAIN(9) => DATAIN(9), 
                           DATAIN(8) => DATAIN(8), DATAIN(7) => DATAIN(7), 
                           DATAIN(6) => DATAIN(6), DATAIN(5) => DATAIN(5), 
                           DATAIN(4) => DATAIN(4), DATAIN(3) => DATAIN(3), 
                           DATAIN(2) => DATAIN(2), DATAIN(1) => DATAIN(1), 
                           DATAIN(0) => DATAIN(0), OUT1(31) => A_out(31), 
                           OUT1(30) => A_out(30), OUT1(29) => A_out(29), 
                           OUT1(28) => A_out(28), OUT1(27) => A_out(27), 
                           OUT1(26) => A_out(26), OUT1(25) => A_out(25), 
                           OUT1(24) => A_out(24), OUT1(23) => A_out(23), 
                           OUT1(22) => A_out(22), OUT1(21) => A_out(21), 
                           OUT1(20) => A_out(20), OUT1(19) => A_out(19), 
                           OUT1(18) => A_out(18), OUT1(17) => A_out(17), 
                           OUT1(16) => A_out(16), OUT1(15) => A_out(15), 
                           OUT1(14) => A_out(14), OUT1(13) => A_out(13), 
                           OUT1(12) => A_out(12), OUT1(11) => A_out(11), 
                           OUT1(10) => A_out(10), OUT1(9) => A_out(9), OUT1(8) 
                           => A_out(8), OUT1(7) => A_out(7), OUT1(6) => 
                           A_out(6), OUT1(5) => A_out(5), OUT1(4) => A_out(4), 
                           OUT1(3) => A_out(3), OUT1(2) => A_out(2), OUT1(1) =>
                           A_out(1), OUT1(0) => A_out(0), OUT2(31) => B_out(31)
                           , OUT2(30) => B_out(30), OUT2(29) => B_out(29), 
                           OUT2(28) => B_out(28), OUT2(27) => B_out(27), 
                           OUT2(26) => B_out(26), OUT2(25) => B_out(25), 
                           OUT2(24) => B_out(24), OUT2(23) => B_out(23), 
                           OUT2(22) => B_out(22), OUT2(21) => B_out(21), 
                           OUT2(20) => B_out(20), OUT2(19) => B_out(19), 
                           OUT2(18) => B_out(18), OUT2(17) => B_out(17), 
                           OUT2(16) => B_out(16), OUT2(15) => B_out(15), 
                           OUT2(14) => B_out(14), OUT2(13) => B_out(13), 
                           OUT2(12) => B_out(12), OUT2(11) => B_out(11), 
                           OUT2(10) => B_out(10), OUT2(9) => B_out(9), OUT2(8) 
                           => B_out(8), OUT2(7) => B_out(7), OUT2(6) => 
                           B_out(6), OUT2(5) => B_out(5), OUT2(4) => B_out(4), 
                           OUT2(3) => B_out(3), OUT2(2) => B_out(2), OUT2(1) =>
                           B_out(1), OUT2(0) => B_out(0));
   U2 : NOR4_X2 port map( A1 => IR_IN2(28), A2 => IR_IN2(27), A3 => IR_IN2(26),
                           A4 => n4, ZN => n3);
   U3 : BUF_X1 port map( A => clk, Z => n2);
   U4 : BUF_X1 port map( A => rst, Z => n1);
   U5 : MUX2_X1 port map( A => IR_IN2(16), B => IR_IN2(11), S => n3, Z => n5);
   U6 : MUX2_X1 port map( A => IR_IN2(17), B => IR_IN2(12), S => n3, Z => n6);
   U7 : MUX2_X1 port map( A => IR_IN2(18), B => IR_IN2(13), S => n3, Z => n7);
   U8 : MUX2_X1 port map( A => IR_IN2(19), B => IR_IN2(14), S => n3, Z => n8);
   U9 : MUX2_X1 port map( A => IR_IN2(20), B => IR_IN2(15), S => n3, Z => n9);
   U10 : OR3_X1 port map( A1 => IR_IN2(31), A2 => IR_IN2(30), A3 => IR_IN2(29),
                           ZN => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity fetchUnit_nbits32 is

   port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 downto 
         0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN : in std_logic;  PC_IN : 
         in std_logic_vector (31 downto 0);  ADDRESS_IRAM, NPC_OUT, IR_OUT, 
         ADDERPC_OUT : out std_logic_vector (31 downto 0));

end fetchUnit_nbits32;

architecture SYN_STRUCTURAL of fetchUnit_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component register_generic_nbits32_9
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_10
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_0
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component RCA_NBITS32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ADDRESS_IRAM_31_port, 
      ADDRESS_IRAM_30_port, ADDRESS_IRAM_29_port, ADDRESS_IRAM_28_port, 
      ADDRESS_IRAM_27_port, ADDRESS_IRAM_26_port, ADDRESS_IRAM_25_port, 
      ADDRESS_IRAM_24_port, ADDRESS_IRAM_23_port, ADDRESS_IRAM_22_port, 
      ADDRESS_IRAM_21_port, ADDRESS_IRAM_20_port, ADDRESS_IRAM_19_port, 
      ADDRESS_IRAM_18_port, ADDRESS_IRAM_17_port, ADDRESS_IRAM_16_port, 
      ADDRESS_IRAM_15_port, ADDRESS_IRAM_14_port, ADDRESS_IRAM_13_port, 
      ADDRESS_IRAM_12_port, ADDRESS_IRAM_11_port, ADDRESS_IRAM_10_port, 
      ADDRESS_IRAM_9_port, ADDRESS_IRAM_8_port, ADDRESS_IRAM_7_port, 
      ADDRESS_IRAM_6_port, ADDRESS_IRAM_5_port, ADDRESS_IRAM_4_port, 
      ADDRESS_IRAM_3_port, ADDRESS_IRAM_2_port, ADDRESS_IRAM_1_port, 
      ADDRESS_IRAM_0_port, ADDERPC_OUT_31_port, ADDERPC_OUT_30_port, 
      ADDERPC_OUT_29_port, ADDERPC_OUT_28_port, ADDERPC_OUT_27_port, 
      ADDERPC_OUT_26_port, ADDERPC_OUT_25_port, ADDERPC_OUT_24_port, 
      ADDERPC_OUT_23_port, ADDERPC_OUT_22_port, ADDERPC_OUT_21_port, 
      ADDERPC_OUT_20_port, ADDERPC_OUT_19_port, ADDERPC_OUT_18_port, 
      ADDERPC_OUT_17_port, ADDERPC_OUT_16_port, ADDERPC_OUT_15_port, 
      ADDERPC_OUT_14_port, ADDERPC_OUT_13_port, ADDERPC_OUT_12_port, 
      ADDERPC_OUT_11_port, ADDERPC_OUT_10_port, ADDERPC_OUT_9_port, 
      ADDERPC_OUT_8_port, ADDERPC_OUT_7_port, ADDERPC_OUT_6_port, 
      ADDERPC_OUT_5_port, ADDERPC_OUT_4_port, ADDERPC_OUT_3_port, 
      ADDERPC_OUT_2_port, ADDERPC_OUT_1_port, ADDERPC_OUT_0_port, n1, n2, 
      n_1404 : std_logic;

begin
   ADDRESS_IRAM <= ( ADDRESS_IRAM_31_port, ADDRESS_IRAM_30_port, 
      ADDRESS_IRAM_29_port, ADDRESS_IRAM_28_port, ADDRESS_IRAM_27_port, 
      ADDRESS_IRAM_26_port, ADDRESS_IRAM_25_port, ADDRESS_IRAM_24_port, 
      ADDRESS_IRAM_23_port, ADDRESS_IRAM_22_port, ADDRESS_IRAM_21_port, 
      ADDRESS_IRAM_20_port, ADDRESS_IRAM_19_port, ADDRESS_IRAM_18_port, 
      ADDRESS_IRAM_17_port, ADDRESS_IRAM_16_port, ADDRESS_IRAM_15_port, 
      ADDRESS_IRAM_14_port, ADDRESS_IRAM_13_port, ADDRESS_IRAM_12_port, 
      ADDRESS_IRAM_11_port, ADDRESS_IRAM_10_port, ADDRESS_IRAM_9_port, 
      ADDRESS_IRAM_8_port, ADDRESS_IRAM_7_port, ADDRESS_IRAM_6_port, 
      ADDRESS_IRAM_5_port, ADDRESS_IRAM_4_port, ADDRESS_IRAM_3_port, 
      ADDRESS_IRAM_2_port, ADDRESS_IRAM_1_port, ADDRESS_IRAM_0_port );
   ADDERPC_OUT <= ( ADDERPC_OUT_31_port, ADDERPC_OUT_30_port, 
      ADDERPC_OUT_29_port, ADDERPC_OUT_28_port, ADDERPC_OUT_27_port, 
      ADDERPC_OUT_26_port, ADDERPC_OUT_25_port, ADDERPC_OUT_24_port, 
      ADDERPC_OUT_23_port, ADDERPC_OUT_22_port, ADDERPC_OUT_21_port, 
      ADDERPC_OUT_20_port, ADDERPC_OUT_19_port, ADDERPC_OUT_18_port, 
      ADDERPC_OUT_17_port, ADDERPC_OUT_16_port, ADDERPC_OUT_15_port, 
      ADDERPC_OUT_14_port, ADDERPC_OUT_13_port, ADDERPC_OUT_12_port, 
      ADDERPC_OUT_11_port, ADDERPC_OUT_10_port, ADDERPC_OUT_9_port, 
      ADDERPC_OUT_8_port, ADDERPC_OUT_7_port, ADDERPC_OUT_6_port, 
      ADDERPC_OUT_5_port, ADDERPC_OUT_4_port, ADDERPC_OUT_3_port, 
      ADDERPC_OUT_2_port, ADDERPC_OUT_1_port, ADDERPC_OUT_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADD : RCA_NBITS32 port map( A(31) => ADDRESS_IRAM_31_port, A(30) => 
                           ADDRESS_IRAM_30_port, A(29) => ADDRESS_IRAM_29_port,
                           A(28) => ADDRESS_IRAM_28_port, A(27) => 
                           ADDRESS_IRAM_27_port, A(26) => ADDRESS_IRAM_26_port,
                           A(25) => ADDRESS_IRAM_25_port, A(24) => 
                           ADDRESS_IRAM_24_port, A(23) => ADDRESS_IRAM_23_port,
                           A(22) => ADDRESS_IRAM_22_port, A(21) => 
                           ADDRESS_IRAM_21_port, A(20) => ADDRESS_IRAM_20_port,
                           A(19) => ADDRESS_IRAM_19_port, A(18) => 
                           ADDRESS_IRAM_18_port, A(17) => ADDRESS_IRAM_17_port,
                           A(16) => ADDRESS_IRAM_16_port, A(15) => 
                           ADDRESS_IRAM_15_port, A(14) => ADDRESS_IRAM_14_port,
                           A(13) => ADDRESS_IRAM_13_port, A(12) => 
                           ADDRESS_IRAM_12_port, A(11) => ADDRESS_IRAM_11_port,
                           A(10) => ADDRESS_IRAM_10_port, A(9) => 
                           ADDRESS_IRAM_9_port, A(8) => ADDRESS_IRAM_8_port, 
                           A(7) => ADDRESS_IRAM_7_port, A(6) => 
                           ADDRESS_IRAM_6_port, A(5) => ADDRESS_IRAM_5_port, 
                           A(4) => ADDRESS_IRAM_4_port, A(3) => 
                           ADDRESS_IRAM_3_port, A(2) => ADDRESS_IRAM_2_port, 
                           A(1) => ADDRESS_IRAM_1_port, A(0) => 
                           ADDRESS_IRAM_0_port, B(31) => X_Logic0_port, B(30) 
                           => X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic1_port, Ci => X_Logic0_port, S(31) => 
                           ADDERPC_OUT_31_port, S(30) => ADDERPC_OUT_30_port, 
                           S(29) => ADDERPC_OUT_29_port, S(28) => 
                           ADDERPC_OUT_28_port, S(27) => ADDERPC_OUT_27_port, 
                           S(26) => ADDERPC_OUT_26_port, S(25) => 
                           ADDERPC_OUT_25_port, S(24) => ADDERPC_OUT_24_port, 
                           S(23) => ADDERPC_OUT_23_port, S(22) => 
                           ADDERPC_OUT_22_port, S(21) => ADDERPC_OUT_21_port, 
                           S(20) => ADDERPC_OUT_20_port, S(19) => 
                           ADDERPC_OUT_19_port, S(18) => ADDERPC_OUT_18_port, 
                           S(17) => ADDERPC_OUT_17_port, S(16) => 
                           ADDERPC_OUT_16_port, S(15) => ADDERPC_OUT_15_port, 
                           S(14) => ADDERPC_OUT_14_port, S(13) => 
                           ADDERPC_OUT_13_port, S(12) => ADDERPC_OUT_12_port, 
                           S(11) => ADDERPC_OUT_11_port, S(10) => 
                           ADDERPC_OUT_10_port, S(9) => ADDERPC_OUT_9_port, 
                           S(8) => ADDERPC_OUT_8_port, S(7) => 
                           ADDERPC_OUT_7_port, S(6) => ADDERPC_OUT_6_port, S(5)
                           => ADDERPC_OUT_5_port, S(4) => ADDERPC_OUT_4_port, 
                           S(3) => ADDERPC_OUT_3_port, S(2) => 
                           ADDERPC_OUT_2_port, S(1) => ADDERPC_OUT_1_port, S(0)
                           => ADDERPC_OUT_0_port, Co => n_1404);
   PC : register_generic_nbits32_0 port map( data_in(31) => PC_IN(31), 
                           data_in(30) => PC_IN(30), data_in(29) => PC_IN(29), 
                           data_in(28) => PC_IN(28), data_in(27) => PC_IN(27), 
                           data_in(26) => PC_IN(26), data_in(25) => PC_IN(25), 
                           data_in(24) => PC_IN(24), data_in(23) => PC_IN(23), 
                           data_in(22) => PC_IN(22), data_in(21) => PC_IN(21), 
                           data_in(20) => PC_IN(20), data_in(19) => PC_IN(19), 
                           data_in(18) => PC_IN(18), data_in(17) => PC_IN(17), 
                           data_in(16) => PC_IN(16), data_in(15) => PC_IN(15), 
                           data_in(14) => PC_IN(14), data_in(13) => PC_IN(13), 
                           data_in(12) => PC_IN(12), data_in(11) => PC_IN(11), 
                           data_in(10) => PC_IN(10), data_in(9) => PC_IN(9), 
                           data_in(8) => PC_IN(8), data_in(7) => PC_IN(7), 
                           data_in(6) => PC_IN(6), data_in(5) => PC_IN(5), 
                           data_in(4) => PC_IN(4), data_in(3) => PC_IN(3), 
                           data_in(2) => PC_IN(2), data_in(1) => PC_IN(1), 
                           data_in(0) => PC_IN(0), CK => n2, RESET => n1, 
                           ENABLE => PC_LATCH_EN, data_out(31) => 
                           ADDRESS_IRAM_31_port, data_out(30) => 
                           ADDRESS_IRAM_30_port, data_out(29) => 
                           ADDRESS_IRAM_29_port, data_out(28) => 
                           ADDRESS_IRAM_28_port, data_out(27) => 
                           ADDRESS_IRAM_27_port, data_out(26) => 
                           ADDRESS_IRAM_26_port, data_out(25) => 
                           ADDRESS_IRAM_25_port, data_out(24) => 
                           ADDRESS_IRAM_24_port, data_out(23) => 
                           ADDRESS_IRAM_23_port, data_out(22) => 
                           ADDRESS_IRAM_22_port, data_out(21) => 
                           ADDRESS_IRAM_21_port, data_out(20) => 
                           ADDRESS_IRAM_20_port, data_out(19) => 
                           ADDRESS_IRAM_19_port, data_out(18) => 
                           ADDRESS_IRAM_18_port, data_out(17) => 
                           ADDRESS_IRAM_17_port, data_out(16) => 
                           ADDRESS_IRAM_16_port, data_out(15) => 
                           ADDRESS_IRAM_15_port, data_out(14) => 
                           ADDRESS_IRAM_14_port, data_out(13) => 
                           ADDRESS_IRAM_13_port, data_out(12) => 
                           ADDRESS_IRAM_12_port, data_out(11) => 
                           ADDRESS_IRAM_11_port, data_out(10) => 
                           ADDRESS_IRAM_10_port, data_out(9) => 
                           ADDRESS_IRAM_9_port, data_out(8) => 
                           ADDRESS_IRAM_8_port, data_out(7) => 
                           ADDRESS_IRAM_7_port, data_out(6) => 
                           ADDRESS_IRAM_6_port, data_out(5) => 
                           ADDRESS_IRAM_5_port, data_out(4) => 
                           ADDRESS_IRAM_4_port, data_out(3) => 
                           ADDRESS_IRAM_3_port, data_out(2) => 
                           ADDRESS_IRAM_2_port, data_out(1) => 
                           ADDRESS_IRAM_1_port, data_out(0) => 
                           ADDRESS_IRAM_0_port);
   IR : register_generic_nbits32_10 port map( data_in(31) => DATA_IRAM(31), 
                           data_in(30) => DATA_IRAM(30), data_in(29) => 
                           DATA_IRAM(29), data_in(28) => DATA_IRAM(28), 
                           data_in(27) => DATA_IRAM(27), data_in(26) => 
                           DATA_IRAM(26), data_in(25) => DATA_IRAM(25), 
                           data_in(24) => DATA_IRAM(24), data_in(23) => 
                           DATA_IRAM(23), data_in(22) => DATA_IRAM(22), 
                           data_in(21) => DATA_IRAM(21), data_in(20) => 
                           DATA_IRAM(20), data_in(19) => DATA_IRAM(19), 
                           data_in(18) => DATA_IRAM(18), data_in(17) => 
                           DATA_IRAM(17), data_in(16) => DATA_IRAM(16), 
                           data_in(15) => DATA_IRAM(15), data_in(14) => 
                           DATA_IRAM(14), data_in(13) => DATA_IRAM(13), 
                           data_in(12) => DATA_IRAM(12), data_in(11) => 
                           DATA_IRAM(11), data_in(10) => DATA_IRAM(10), 
                           data_in(9) => DATA_IRAM(9), data_in(8) => 
                           DATA_IRAM(8), data_in(7) => DATA_IRAM(7), data_in(6)
                           => DATA_IRAM(6), data_in(5) => DATA_IRAM(5), 
                           data_in(4) => DATA_IRAM(4), data_in(3) => 
                           DATA_IRAM(3), data_in(2) => DATA_IRAM(2), data_in(1)
                           => DATA_IRAM(1), data_in(0) => DATA_IRAM(0), CK => 
                           n2, RESET => n1, ENABLE => IR_LATCH_EN, data_out(31)
                           => IR_OUT(31), data_out(30) => IR_OUT(30), 
                           data_out(29) => IR_OUT(29), data_out(28) => 
                           IR_OUT(28), data_out(27) => IR_OUT(27), data_out(26)
                           => IR_OUT(26), data_out(25) => IR_OUT(25), 
                           data_out(24) => IR_OUT(24), data_out(23) => 
                           IR_OUT(23), data_out(22) => IR_OUT(22), data_out(21)
                           => IR_OUT(21), data_out(20) => IR_OUT(20), 
                           data_out(19) => IR_OUT(19), data_out(18) => 
                           IR_OUT(18), data_out(17) => IR_OUT(17), data_out(16)
                           => IR_OUT(16), data_out(15) => IR_OUT(15), 
                           data_out(14) => IR_OUT(14), data_out(13) => 
                           IR_OUT(13), data_out(12) => IR_OUT(12), data_out(11)
                           => IR_OUT(11), data_out(10) => IR_OUT(10), 
                           data_out(9) => IR_OUT(9), data_out(8) => IR_OUT(8), 
                           data_out(7) => IR_OUT(7), data_out(6) => IR_OUT(6), 
                           data_out(5) => IR_OUT(5), data_out(4) => IR_OUT(4), 
                           data_out(3) => IR_OUT(3), data_out(2) => IR_OUT(2), 
                           data_out(1) => IR_OUT(1), data_out(0) => IR_OUT(0));
   NPC : register_generic_nbits32_9 port map( data_in(31) => 
                           ADDERPC_OUT_31_port, data_in(30) => 
                           ADDERPC_OUT_30_port, data_in(29) => 
                           ADDERPC_OUT_29_port, data_in(28) => 
                           ADDERPC_OUT_28_port, data_in(27) => 
                           ADDERPC_OUT_27_port, data_in(26) => 
                           ADDERPC_OUT_26_port, data_in(25) => 
                           ADDERPC_OUT_25_port, data_in(24) => 
                           ADDERPC_OUT_24_port, data_in(23) => 
                           ADDERPC_OUT_23_port, data_in(22) => 
                           ADDERPC_OUT_22_port, data_in(21) => 
                           ADDERPC_OUT_21_port, data_in(20) => 
                           ADDERPC_OUT_20_port, data_in(19) => 
                           ADDERPC_OUT_19_port, data_in(18) => 
                           ADDERPC_OUT_18_port, data_in(17) => 
                           ADDERPC_OUT_17_port, data_in(16) => 
                           ADDERPC_OUT_16_port, data_in(15) => 
                           ADDERPC_OUT_15_port, data_in(14) => 
                           ADDERPC_OUT_14_port, data_in(13) => 
                           ADDERPC_OUT_13_port, data_in(12) => 
                           ADDERPC_OUT_12_port, data_in(11) => 
                           ADDERPC_OUT_11_port, data_in(10) => 
                           ADDERPC_OUT_10_port, data_in(9) => 
                           ADDERPC_OUT_9_port, data_in(8) => ADDERPC_OUT_8_port
                           , data_in(7) => ADDERPC_OUT_7_port, data_in(6) => 
                           ADDERPC_OUT_6_port, data_in(5) => ADDERPC_OUT_5_port
                           , data_in(4) => ADDERPC_OUT_4_port, data_in(3) => 
                           ADDERPC_OUT_3_port, data_in(2) => ADDERPC_OUT_2_port
                           , data_in(1) => ADDERPC_OUT_1_port, data_in(0) => 
                           ADDERPC_OUT_0_port, CK => n2, RESET => n1, ENABLE =>
                           NPC_LATCH_EN, data_out(31) => NPC_OUT(31), 
                           data_out(30) => NPC_OUT(30), data_out(29) => 
                           NPC_OUT(29), data_out(28) => NPC_OUT(28), 
                           data_out(27) => NPC_OUT(27), data_out(26) => 
                           NPC_OUT(26), data_out(25) => NPC_OUT(25), 
                           data_out(24) => NPC_OUT(24), data_out(23) => 
                           NPC_OUT(23), data_out(22) => NPC_OUT(22), 
                           data_out(21) => NPC_OUT(21), data_out(20) => 
                           NPC_OUT(20), data_out(19) => NPC_OUT(19), 
                           data_out(18) => NPC_OUT(18), data_out(17) => 
                           NPC_OUT(17), data_out(16) => NPC_OUT(16), 
                           data_out(15) => NPC_OUT(15), data_out(14) => 
                           NPC_OUT(14), data_out(13) => NPC_OUT(13), 
                           data_out(12) => NPC_OUT(12), data_out(11) => 
                           NPC_OUT(11), data_out(10) => NPC_OUT(10), 
                           data_out(9) => NPC_OUT(9), data_out(8) => NPC_OUT(8)
                           , data_out(7) => NPC_OUT(7), data_out(6) => 
                           NPC_OUT(6), data_out(5) => NPC_OUT(5), data_out(4) 
                           => NPC_OUT(4), data_out(3) => NPC_OUT(3), 
                           data_out(2) => NPC_OUT(2), data_out(1) => NPC_OUT(1)
                           , data_out(0) => NPC_OUT(0));
   U3 : BUF_X1 port map( A => rst, Z => n1);
   U4 : BUF_X1 port map( A => clk, Z => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity datapath_nbits32 is

   port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 downto 
         0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN, RegA_LATCH_EN, 
         RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE, MUXA_SEL, MUXB_SEL, 
         ALU_OUTREG_EN, EQ_COND : in std_logic;  ALU_OPCODE : in 
         std_logic_vector (0 to 3);  DRAM_DATA : in std_logic_vector (31 downto
         0);  LMD_LATCH_EN, JUMP_EN, WB_MUX_SEL : in std_logic;  B, ALU_OUT, 
         ADDRESS_IRAM, IR_OUT : out std_logic_vector (31 downto 0));

end datapath_nbits32;

architecture SYN_STRUCTURAL of datapath_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component writeBack_nbits32
      port( LMD_OUT, ALUREG_OUTPUT : in std_logic_vector (31 downto 0);  
            WB_MUX_SEL : in std_logic;  DATAIN_RF : out std_logic_vector (31 
            downto 0));
   end component;
   
   component memoryUnit_nbits32
      port( clk, rst, LMD_LATCH_EN, JUMP_EN : in std_logic;  DRAM_DATA, 
            ALUREG_OUTPUT, NPC_OUT : in std_logic_vector (31 downto 0);  
            COND_OUT : in std_logic;  DRAM_DATAout, TO_PC_OUT, ALU_OUT2 : out 
            std_logic_vector (31 downto 0);  IR_IN4 : in std_logic_vector (31 
            downto 0);  IR_OUT4 : out std_logic_vector (31 downto 0));
   end component;
   
   component executionUnit_nbits32
      port( clk, rst, ALU_OUTREG_ENABLE, MUXA_SEL, MUXB_SEL, COND_ENABLE : in 
            std_logic;  ALU_BITS : in std_logic_vector (0 to 3);  NPC_OUT, 
            A_out, B_out, Imm_out : in std_logic_vector (31 downto 0);  
            ALUREG_OUTPUT : out std_logic_vector (31 downto 0);  COND_OUT : out
            std_logic;  IR_IN3 : in std_logic_vector (31 downto 0);  IR_OUT3, 
            B_outreg : out std_logic_vector (31 downto 0));
   end component;
   
   component decodeUnit_nbits32
      port( clk, rst, RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE : in
            std_logic;  DATAIN, IR_OUT : in std_logic_vector (31 downto 0);  
            A_out, B_out, Imm_out : out std_logic_vector (31 downto 0);  IR_IN2
            : in std_logic_vector (31 downto 0);  IR_OUT2 : out 
            std_logic_vector (31 downto 0);  NPC_IN : in std_logic_vector (31 
            downto 0);  NPC2_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component fetchUnit_nbits32
      port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 
            downto 0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN : in std_logic; 
            PC_IN : in std_logic_vector (31 downto 0);  ADDRESS_IRAM, NPC_OUT, 
            IR_OUT, ADDERPC_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal ALU_OUT_31_port, ALU_OUT_30_port, ALU_OUT_29_port, ALU_OUT_28_port, 
      ALU_OUT_27_port, ALU_OUT_26_port, ALU_OUT_25_port, ALU_OUT_24_port, 
      ALU_OUT_23_port, ALU_OUT_22_port, ALU_OUT_21_port, ALU_OUT_20_port, 
      ALU_OUT_19_port, ALU_OUT_18_port, ALU_OUT_17_port, ALU_OUT_16_port, 
      ALU_OUT_15_port, ALU_OUT_14_port, ALU_OUT_13_port, ALU_OUT_12_port, 
      ALU_OUT_11_port, ALU_OUT_10_port, ALU_OUT_9_port, ALU_OUT_8_port, 
      ALU_OUT_7_port, ALU_OUT_6_port, ALU_OUT_5_port, ALU_OUT_4_port, 
      ALU_OUT_3_port, ALU_OUT_2_port, ALU_OUT_1_port, ALU_OUT_0_port, 
      IR_OUT_31_port, IR_OUT_30_port, IR_OUT_29_port, IR_OUT_28_port, 
      IR_OUT_27_port, IR_OUT_26_port, IR_OUT_25_port, IR_OUT_24_port, 
      IR_OUT_23_port, IR_OUT_22_port, IR_OUT_21_port, IR_OUT_20_port, 
      IR_OUT_19_port, IR_OUT_18_port, IR_OUT_17_port, IR_OUT_16_port, 
      IR_OUT_15_port, IR_OUT_14_port, IR_OUT_13_port, IR_OUT_12_port, 
      IR_OUT_11_port, IR_OUT_10_port, IR_OUT_9_port, IR_OUT_8_port, 
      IR_OUT_7_port, IR_OUT_6_port, IR_OUT_5_port, IR_OUT_4_port, IR_OUT_3_port
      , IR_OUT_2_port, IR_OUT_1_port, IR_OUT_0_port, TO_PC_OUTs_31_port, 
      TO_PC_OUTs_30_port, TO_PC_OUTs_29_port, TO_PC_OUTs_28_port, 
      TO_PC_OUTs_27_port, TO_PC_OUTs_26_port, TO_PC_OUTs_25_port, 
      TO_PC_OUTs_24_port, TO_PC_OUTs_23_port, TO_PC_OUTs_22_port, 
      TO_PC_OUTs_21_port, TO_PC_OUTs_20_port, TO_PC_OUTs_19_port, 
      TO_PC_OUTs_18_port, TO_PC_OUTs_17_port, TO_PC_OUTs_16_port, 
      TO_PC_OUTs_15_port, TO_PC_OUTs_14_port, TO_PC_OUTs_13_port, 
      TO_PC_OUTs_12_port, TO_PC_OUTs_11_port, TO_PC_OUTs_10_port, 
      TO_PC_OUTs_9_port, TO_PC_OUTs_8_port, TO_PC_OUTs_7_port, 
      TO_PC_OUTs_6_port, TO_PC_OUTs_5_port, TO_PC_OUTs_4_port, 
      TO_PC_OUTs_3_port, TO_PC_OUTs_2_port, TO_PC_OUTs_1_port, 
      TO_PC_OUTs_0_port, NPC_OUTs_31_port, NPC_OUTs_30_port, NPC_OUTs_29_port, 
      NPC_OUTs_28_port, NPC_OUTs_27_port, NPC_OUTs_26_port, NPC_OUTs_25_port, 
      NPC_OUTs_24_port, NPC_OUTs_23_port, NPC_OUTs_22_port, NPC_OUTs_21_port, 
      NPC_OUTs_20_port, NPC_OUTs_19_port, NPC_OUTs_18_port, NPC_OUTs_17_port, 
      NPC_OUTs_16_port, NPC_OUTs_15_port, NPC_OUTs_14_port, NPC_OUTs_13_port, 
      NPC_OUTs_12_port, NPC_OUTs_11_port, NPC_OUTs_10_port, NPC_OUTs_9_port, 
      NPC_OUTs_8_port, NPC_OUTs_7_port, NPC_OUTs_6_port, NPC_OUTs_5_port, 
      NPC_OUTs_4_port, NPC_OUTs_3_port, NPC_OUTs_2_port, NPC_OUTs_1_port, 
      NPC_OUTs_0_port, ADDERPC_OUTs_31_port, ADDERPC_OUTs_30_port, 
      ADDERPC_OUTs_29_port, ADDERPC_OUTs_28_port, ADDERPC_OUTs_27_port, 
      ADDERPC_OUTs_26_port, ADDERPC_OUTs_25_port, ADDERPC_OUTs_24_port, 
      ADDERPC_OUTs_23_port, ADDERPC_OUTs_22_port, ADDERPC_OUTs_21_port, 
      ADDERPC_OUTs_20_port, ADDERPC_OUTs_19_port, ADDERPC_OUTs_18_port, 
      ADDERPC_OUTs_17_port, ADDERPC_OUTs_16_port, ADDERPC_OUTs_15_port, 
      ADDERPC_OUTs_14_port, ADDERPC_OUTs_13_port, ADDERPC_OUTs_12_port, 
      ADDERPC_OUTs_11_port, ADDERPC_OUTs_10_port, ADDERPC_OUTs_9_port, 
      ADDERPC_OUTs_8_port, ADDERPC_OUTs_7_port, ADDERPC_OUTs_6_port, 
      ADDERPC_OUTs_5_port, ADDERPC_OUTs_4_port, ADDERPC_OUTs_3_port, 
      ADDERPC_OUTs_2_port, ADDERPC_OUTs_1_port, ADDERPC_OUTs_0_port, 
      DATAIN_RFs_31_port, DATAIN_RFs_30_port, DATAIN_RFs_29_port, 
      DATAIN_RFs_28_port, DATAIN_RFs_27_port, DATAIN_RFs_26_port, 
      DATAIN_RFs_25_port, DATAIN_RFs_24_port, DATAIN_RFs_23_port, 
      DATAIN_RFs_22_port, DATAIN_RFs_21_port, DATAIN_RFs_20_port, 
      DATAIN_RFs_19_port, DATAIN_RFs_18_port, DATAIN_RFs_17_port, 
      DATAIN_RFs_16_port, DATAIN_RFs_15_port, DATAIN_RFs_14_port, 
      DATAIN_RFs_13_port, DATAIN_RFs_12_port, DATAIN_RFs_11_port, 
      DATAIN_RFs_10_port, DATAIN_RFs_9_port, DATAIN_RFs_8_port, 
      DATAIN_RFs_7_port, DATAIN_RFs_6_port, DATAIN_RFs_5_port, 
      DATAIN_RFs_4_port, DATAIN_RFs_3_port, DATAIN_RFs_2_port, 
      DATAIN_RFs_1_port, DATAIN_RFs_0_port, A_outs_31_port, A_outs_30_port, 
      A_outs_29_port, A_outs_28_port, A_outs_27_port, A_outs_26_port, 
      A_outs_25_port, A_outs_24_port, A_outs_23_port, A_outs_22_port, 
      A_outs_21_port, A_outs_20_port, A_outs_19_port, A_outs_18_port, 
      A_outs_17_port, A_outs_16_port, A_outs_15_port, A_outs_14_port, 
      A_outs_13_port, A_outs_12_port, A_outs_11_port, A_outs_10_port, 
      A_outs_9_port, A_outs_8_port, A_outs_7_port, A_outs_6_port, A_outs_5_port
      , A_outs_4_port, A_outs_3_port, A_outs_2_port, A_outs_1_port, 
      A_outs_0_port, B_outs_31_port, B_outs_30_port, B_outs_29_port, 
      B_outs_28_port, B_outs_27_port, B_outs_26_port, B_outs_25_port, 
      B_outs_24_port, B_outs_23_port, B_outs_22_port, B_outs_21_port, 
      B_outs_20_port, B_outs_19_port, B_outs_18_port, B_outs_17_port, 
      B_outs_16_port, B_outs_15_port, B_outs_14_port, B_outs_13_port, 
      B_outs_12_port, B_outs_11_port, B_outs_10_port, B_outs_9_port, 
      B_outs_8_port, B_outs_7_port, B_outs_6_port, B_outs_5_port, B_outs_4_port
      , B_outs_3_port, B_outs_2_port, B_outs_1_port, B_outs_0_port, 
      Imm_outs_31_port, Imm_outs_30_port, Imm_outs_29_port, Imm_outs_28_port, 
      Imm_outs_27_port, Imm_outs_26_port, Imm_outs_25_port, Imm_outs_24_port, 
      Imm_outs_23_port, Imm_outs_22_port, Imm_outs_21_port, Imm_outs_20_port, 
      Imm_outs_19_port, Imm_outs_18_port, Imm_outs_17_port, Imm_outs_16_port, 
      Imm_outs_15_port, Imm_outs_14_port, Imm_outs_13_port, Imm_outs_12_port, 
      Imm_outs_11_port, Imm_outs_10_port, Imm_outs_9_port, Imm_outs_8_port, 
      Imm_outs_7_port, Imm_outs_6_port, Imm_outs_5_port, Imm_outs_4_port, 
      Imm_outs_3_port, Imm_outs_2_port, Imm_outs_1_port, Imm_outs_0_port, 
      IR_OUT4s_31_port, IR_OUT4s_30_port, IR_OUT4s_29_port, IR_OUT4s_28_port, 
      IR_OUT4s_27_port, IR_OUT4s_26_port, IR_OUT4s_25_port, IR_OUT4s_24_port, 
      IR_OUT4s_23_port, IR_OUT4s_22_port, IR_OUT4s_21_port, IR_OUT4s_20_port, 
      IR_OUT4s_19_port, IR_OUT4s_18_port, IR_OUT4s_17_port, IR_OUT4s_16_port, 
      IR_OUT4s_15_port, IR_OUT4s_14_port, IR_OUT4s_13_port, IR_OUT4s_12_port, 
      IR_OUT4s_11_port, IR_OUT4s_10_port, IR_OUT4s_9_port, IR_OUT4s_8_port, 
      IR_OUT4s_7_port, IR_OUT4s_6_port, IR_OUT4s_5_port, IR_OUT4s_4_port, 
      IR_OUT4s_3_port, IR_OUT4s_2_port, IR_OUT4s_1_port, IR_OUT4s_0_port, 
      IR_OUT2s_31_port, IR_OUT2s_30_port, IR_OUT2s_29_port, IR_OUT2s_28_port, 
      IR_OUT2s_27_port, IR_OUT2s_26_port, IR_OUT2s_25_port, IR_OUT2s_24_port, 
      IR_OUT2s_23_port, IR_OUT2s_22_port, IR_OUT2s_21_port, IR_OUT2s_20_port, 
      IR_OUT2s_19_port, IR_OUT2s_18_port, IR_OUT2s_17_port, IR_OUT2s_16_port, 
      IR_OUT2s_15_port, IR_OUT2s_14_port, IR_OUT2s_13_port, IR_OUT2s_12_port, 
      IR_OUT2s_11_port, IR_OUT2s_10_port, IR_OUT2s_9_port, IR_OUT2s_8_port, 
      IR_OUT2s_7_port, IR_OUT2s_6_port, IR_OUT2s_5_port, IR_OUT2s_4_port, 
      IR_OUT2s_3_port, IR_OUT2s_2_port, IR_OUT2s_1_port, IR_OUT2s_0_port, 
      NPC2_OUTs_31_port, NPC2_OUTs_30_port, NPC2_OUTs_29_port, 
      NPC2_OUTs_28_port, NPC2_OUTs_27_port, NPC2_OUTs_26_port, 
      NPC2_OUTs_25_port, NPC2_OUTs_24_port, NPC2_OUTs_23_port, 
      NPC2_OUTs_22_port, NPC2_OUTs_21_port, NPC2_OUTs_20_port, 
      NPC2_OUTs_19_port, NPC2_OUTs_18_port, NPC2_OUTs_17_port, 
      NPC2_OUTs_16_port, NPC2_OUTs_15_port, NPC2_OUTs_14_port, 
      NPC2_OUTs_13_port, NPC2_OUTs_12_port, NPC2_OUTs_11_port, 
      NPC2_OUTs_10_port, NPC2_OUTs_9_port, NPC2_OUTs_8_port, NPC2_OUTs_7_port, 
      NPC2_OUTs_6_port, NPC2_OUTs_5_port, NPC2_OUTs_4_port, NPC2_OUTs_3_port, 
      NPC2_OUTs_2_port, NPC2_OUTs_1_port, NPC2_OUTs_0_port, COND_OUTs, 
      IR_OUT3s_31_port, IR_OUT3s_30_port, IR_OUT3s_29_port, IR_OUT3s_28_port, 
      IR_OUT3s_27_port, IR_OUT3s_26_port, IR_OUT3s_25_port, IR_OUT3s_24_port, 
      IR_OUT3s_23_port, IR_OUT3s_22_port, IR_OUT3s_21_port, IR_OUT3s_20_port, 
      IR_OUT3s_19_port, IR_OUT3s_18_port, IR_OUT3s_17_port, IR_OUT3s_16_port, 
      IR_OUT3s_15_port, IR_OUT3s_14_port, IR_OUT3s_13_port, IR_OUT3s_12_port, 
      IR_OUT3s_11_port, IR_OUT3s_10_port, IR_OUT3s_9_port, IR_OUT3s_8_port, 
      IR_OUT3s_7_port, IR_OUT3s_6_port, IR_OUT3s_5_port, IR_OUT3s_4_port, 
      IR_OUT3s_3_port, IR_OUT3s_2_port, IR_OUT3s_1_port, IR_OUT3s_0_port, 
      LMD_OUTs_31_port, LMD_OUTs_30_port, LMD_OUTs_29_port, LMD_OUTs_28_port, 
      LMD_OUTs_27_port, LMD_OUTs_26_port, LMD_OUTs_25_port, LMD_OUTs_24_port, 
      LMD_OUTs_23_port, LMD_OUTs_22_port, LMD_OUTs_21_port, LMD_OUTs_20_port, 
      LMD_OUTs_19_port, LMD_OUTs_18_port, LMD_OUTs_17_port, LMD_OUTs_16_port, 
      LMD_OUTs_15_port, LMD_OUTs_14_port, LMD_OUTs_13_port, LMD_OUTs_12_port, 
      LMD_OUTs_11_port, LMD_OUTs_10_port, LMD_OUTs_9_port, LMD_OUTs_8_port, 
      LMD_OUTs_7_port, LMD_OUTs_6_port, LMD_OUTs_5_port, LMD_OUTs_4_port, 
      LMD_OUTs_3_port, LMD_OUTs_2_port, LMD_OUTs_1_port, LMD_OUTs_0_port, 
      ALU_OUT2s_31_port, ALU_OUT2s_30_port, ALU_OUT2s_29_port, 
      ALU_OUT2s_28_port, ALU_OUT2s_27_port, ALU_OUT2s_26_port, 
      ALU_OUT2s_25_port, ALU_OUT2s_24_port, ALU_OUT2s_23_port, 
      ALU_OUT2s_22_port, ALU_OUT2s_21_port, ALU_OUT2s_20_port, 
      ALU_OUT2s_19_port, ALU_OUT2s_18_port, ALU_OUT2s_17_port, 
      ALU_OUT2s_16_port, ALU_OUT2s_15_port, ALU_OUT2s_14_port, 
      ALU_OUT2s_13_port, ALU_OUT2s_12_port, ALU_OUT2s_11_port, 
      ALU_OUT2s_10_port, ALU_OUT2s_9_port, ALU_OUT2s_8_port, ALU_OUT2s_7_port, 
      ALU_OUT2s_6_port, ALU_OUT2s_5_port, ALU_OUT2s_4_port, ALU_OUT2s_3_port, 
      ALU_OUT2s_2_port, ALU_OUT2s_1_port, ALU_OUT2s_0_port, n1, n2 : std_logic;

begin
   ALU_OUT <= ( ALU_OUT_31_port, ALU_OUT_30_port, ALU_OUT_29_port, 
      ALU_OUT_28_port, ALU_OUT_27_port, ALU_OUT_26_port, ALU_OUT_25_port, 
      ALU_OUT_24_port, ALU_OUT_23_port, ALU_OUT_22_port, ALU_OUT_21_port, 
      ALU_OUT_20_port, ALU_OUT_19_port, ALU_OUT_18_port, ALU_OUT_17_port, 
      ALU_OUT_16_port, ALU_OUT_15_port, ALU_OUT_14_port, ALU_OUT_13_port, 
      ALU_OUT_12_port, ALU_OUT_11_port, ALU_OUT_10_port, ALU_OUT_9_port, 
      ALU_OUT_8_port, ALU_OUT_7_port, ALU_OUT_6_port, ALU_OUT_5_port, 
      ALU_OUT_4_port, ALU_OUT_3_port, ALU_OUT_2_port, ALU_OUT_1_port, 
      ALU_OUT_0_port );
   IR_OUT <= ( IR_OUT_31_port, IR_OUT_30_port, IR_OUT_29_port, IR_OUT_28_port, 
      IR_OUT_27_port, IR_OUT_26_port, IR_OUT_25_port, IR_OUT_24_port, 
      IR_OUT_23_port, IR_OUT_22_port, IR_OUT_21_port, IR_OUT_20_port, 
      IR_OUT_19_port, IR_OUT_18_port, IR_OUT_17_port, IR_OUT_16_port, 
      IR_OUT_15_port, IR_OUT_14_port, IR_OUT_13_port, IR_OUT_12_port, 
      IR_OUT_11_port, IR_OUT_10_port, IR_OUT_9_port, IR_OUT_8_port, 
      IR_OUT_7_port, IR_OUT_6_port, IR_OUT_5_port, IR_OUT_4_port, IR_OUT_3_port
      , IR_OUT_2_port, IR_OUT_1_port, IR_OUT_0_port );
   
   FETCH : fetchUnit_nbits32 port map( clk => n2, rst => n1, DATA_IRAM(31) => 
                           DATA_IRAM(31), DATA_IRAM(30) => DATA_IRAM(30), 
                           DATA_IRAM(29) => DATA_IRAM(29), DATA_IRAM(28) => 
                           DATA_IRAM(28), DATA_IRAM(27) => DATA_IRAM(27), 
                           DATA_IRAM(26) => DATA_IRAM(26), DATA_IRAM(25) => 
                           DATA_IRAM(25), DATA_IRAM(24) => DATA_IRAM(24), 
                           DATA_IRAM(23) => DATA_IRAM(23), DATA_IRAM(22) => 
                           DATA_IRAM(22), DATA_IRAM(21) => DATA_IRAM(21), 
                           DATA_IRAM(20) => DATA_IRAM(20), DATA_IRAM(19) => 
                           DATA_IRAM(19), DATA_IRAM(18) => DATA_IRAM(18), 
                           DATA_IRAM(17) => DATA_IRAM(17), DATA_IRAM(16) => 
                           DATA_IRAM(16), DATA_IRAM(15) => DATA_IRAM(15), 
                           DATA_IRAM(14) => DATA_IRAM(14), DATA_IRAM(13) => 
                           DATA_IRAM(13), DATA_IRAM(12) => DATA_IRAM(12), 
                           DATA_IRAM(11) => DATA_IRAM(11), DATA_IRAM(10) => 
                           DATA_IRAM(10), DATA_IRAM(9) => DATA_IRAM(9), 
                           DATA_IRAM(8) => DATA_IRAM(8), DATA_IRAM(7) => 
                           DATA_IRAM(7), DATA_IRAM(6) => DATA_IRAM(6), 
                           DATA_IRAM(5) => DATA_IRAM(5), DATA_IRAM(4) => 
                           DATA_IRAM(4), DATA_IRAM(3) => DATA_IRAM(3), 
                           DATA_IRAM(2) => DATA_IRAM(2), DATA_IRAM(1) => 
                           DATA_IRAM(1), DATA_IRAM(0) => DATA_IRAM(0), 
                           IR_LATCH_EN => IR_LATCH_EN, NPC_LATCH_EN => 
                           NPC_LATCH_EN, PC_LATCH_EN => PC_LATCH_EN, PC_IN(31) 
                           => TO_PC_OUTs_31_port, PC_IN(30) => 
                           TO_PC_OUTs_30_port, PC_IN(29) => TO_PC_OUTs_29_port,
                           PC_IN(28) => TO_PC_OUTs_28_port, PC_IN(27) => 
                           TO_PC_OUTs_27_port, PC_IN(26) => TO_PC_OUTs_26_port,
                           PC_IN(25) => TO_PC_OUTs_25_port, PC_IN(24) => 
                           TO_PC_OUTs_24_port, PC_IN(23) => TO_PC_OUTs_23_port,
                           PC_IN(22) => TO_PC_OUTs_22_port, PC_IN(21) => 
                           TO_PC_OUTs_21_port, PC_IN(20) => TO_PC_OUTs_20_port,
                           PC_IN(19) => TO_PC_OUTs_19_port, PC_IN(18) => 
                           TO_PC_OUTs_18_port, PC_IN(17) => TO_PC_OUTs_17_port,
                           PC_IN(16) => TO_PC_OUTs_16_port, PC_IN(15) => 
                           TO_PC_OUTs_15_port, PC_IN(14) => TO_PC_OUTs_14_port,
                           PC_IN(13) => TO_PC_OUTs_13_port, PC_IN(12) => 
                           TO_PC_OUTs_12_port, PC_IN(11) => TO_PC_OUTs_11_port,
                           PC_IN(10) => TO_PC_OUTs_10_port, PC_IN(9) => 
                           TO_PC_OUTs_9_port, PC_IN(8) => TO_PC_OUTs_8_port, 
                           PC_IN(7) => TO_PC_OUTs_7_port, PC_IN(6) => 
                           TO_PC_OUTs_6_port, PC_IN(5) => TO_PC_OUTs_5_port, 
                           PC_IN(4) => TO_PC_OUTs_4_port, PC_IN(3) => 
                           TO_PC_OUTs_3_port, PC_IN(2) => TO_PC_OUTs_2_port, 
                           PC_IN(1) => TO_PC_OUTs_1_port, PC_IN(0) => 
                           TO_PC_OUTs_0_port, ADDRESS_IRAM(31) => 
                           ADDRESS_IRAM(31), ADDRESS_IRAM(30) => 
                           ADDRESS_IRAM(30), ADDRESS_IRAM(29) => 
                           ADDRESS_IRAM(29), ADDRESS_IRAM(28) => 
                           ADDRESS_IRAM(28), ADDRESS_IRAM(27) => 
                           ADDRESS_IRAM(27), ADDRESS_IRAM(26) => 
                           ADDRESS_IRAM(26), ADDRESS_IRAM(25) => 
                           ADDRESS_IRAM(25), ADDRESS_IRAM(24) => 
                           ADDRESS_IRAM(24), ADDRESS_IRAM(23) => 
                           ADDRESS_IRAM(23), ADDRESS_IRAM(22) => 
                           ADDRESS_IRAM(22), ADDRESS_IRAM(21) => 
                           ADDRESS_IRAM(21), ADDRESS_IRAM(20) => 
                           ADDRESS_IRAM(20), ADDRESS_IRAM(19) => 
                           ADDRESS_IRAM(19), ADDRESS_IRAM(18) => 
                           ADDRESS_IRAM(18), ADDRESS_IRAM(17) => 
                           ADDRESS_IRAM(17), ADDRESS_IRAM(16) => 
                           ADDRESS_IRAM(16), ADDRESS_IRAM(15) => 
                           ADDRESS_IRAM(15), ADDRESS_IRAM(14) => 
                           ADDRESS_IRAM(14), ADDRESS_IRAM(13) => 
                           ADDRESS_IRAM(13), ADDRESS_IRAM(12) => 
                           ADDRESS_IRAM(12), ADDRESS_IRAM(11) => 
                           ADDRESS_IRAM(11), ADDRESS_IRAM(10) => 
                           ADDRESS_IRAM(10), ADDRESS_IRAM(9) => ADDRESS_IRAM(9)
                           , ADDRESS_IRAM(8) => ADDRESS_IRAM(8), 
                           ADDRESS_IRAM(7) => ADDRESS_IRAM(7), ADDRESS_IRAM(6) 
                           => ADDRESS_IRAM(6), ADDRESS_IRAM(5) => 
                           ADDRESS_IRAM(5), ADDRESS_IRAM(4) => ADDRESS_IRAM(4),
                           ADDRESS_IRAM(3) => ADDRESS_IRAM(3), ADDRESS_IRAM(2) 
                           => ADDRESS_IRAM(2), ADDRESS_IRAM(1) => 
                           ADDRESS_IRAM(1), ADDRESS_IRAM(0) => ADDRESS_IRAM(0),
                           NPC_OUT(31) => NPC_OUTs_31_port, NPC_OUT(30) => 
                           NPC_OUTs_30_port, NPC_OUT(29) => NPC_OUTs_29_port, 
                           NPC_OUT(28) => NPC_OUTs_28_port, NPC_OUT(27) => 
                           NPC_OUTs_27_port, NPC_OUT(26) => NPC_OUTs_26_port, 
                           NPC_OUT(25) => NPC_OUTs_25_port, NPC_OUT(24) => 
                           NPC_OUTs_24_port, NPC_OUT(23) => NPC_OUTs_23_port, 
                           NPC_OUT(22) => NPC_OUTs_22_port, NPC_OUT(21) => 
                           NPC_OUTs_21_port, NPC_OUT(20) => NPC_OUTs_20_port, 
                           NPC_OUT(19) => NPC_OUTs_19_port, NPC_OUT(18) => 
                           NPC_OUTs_18_port, NPC_OUT(17) => NPC_OUTs_17_port, 
                           NPC_OUT(16) => NPC_OUTs_16_port, NPC_OUT(15) => 
                           NPC_OUTs_15_port, NPC_OUT(14) => NPC_OUTs_14_port, 
                           NPC_OUT(13) => NPC_OUTs_13_port, NPC_OUT(12) => 
                           NPC_OUTs_12_port, NPC_OUT(11) => NPC_OUTs_11_port, 
                           NPC_OUT(10) => NPC_OUTs_10_port, NPC_OUT(9) => 
                           NPC_OUTs_9_port, NPC_OUT(8) => NPC_OUTs_8_port, 
                           NPC_OUT(7) => NPC_OUTs_7_port, NPC_OUT(6) => 
                           NPC_OUTs_6_port, NPC_OUT(5) => NPC_OUTs_5_port, 
                           NPC_OUT(4) => NPC_OUTs_4_port, NPC_OUT(3) => 
                           NPC_OUTs_3_port, NPC_OUT(2) => NPC_OUTs_2_port, 
                           NPC_OUT(1) => NPC_OUTs_1_port, NPC_OUT(0) => 
                           NPC_OUTs_0_port, IR_OUT(31) => IR_OUT_31_port, 
                           IR_OUT(30) => IR_OUT_30_port, IR_OUT(29) => 
                           IR_OUT_29_port, IR_OUT(28) => IR_OUT_28_port, 
                           IR_OUT(27) => IR_OUT_27_port, IR_OUT(26) => 
                           IR_OUT_26_port, IR_OUT(25) => IR_OUT_25_port, 
                           IR_OUT(24) => IR_OUT_24_port, IR_OUT(23) => 
                           IR_OUT_23_port, IR_OUT(22) => IR_OUT_22_port, 
                           IR_OUT(21) => IR_OUT_21_port, IR_OUT(20) => 
                           IR_OUT_20_port, IR_OUT(19) => IR_OUT_19_port, 
                           IR_OUT(18) => IR_OUT_18_port, IR_OUT(17) => 
                           IR_OUT_17_port, IR_OUT(16) => IR_OUT_16_port, 
                           IR_OUT(15) => IR_OUT_15_port, IR_OUT(14) => 
                           IR_OUT_14_port, IR_OUT(13) => IR_OUT_13_port, 
                           IR_OUT(12) => IR_OUT_12_port, IR_OUT(11) => 
                           IR_OUT_11_port, IR_OUT(10) => IR_OUT_10_port, 
                           IR_OUT(9) => IR_OUT_9_port, IR_OUT(8) => 
                           IR_OUT_8_port, IR_OUT(7) => IR_OUT_7_port, IR_OUT(6)
                           => IR_OUT_6_port, IR_OUT(5) => IR_OUT_5_port, 
                           IR_OUT(4) => IR_OUT_4_port, IR_OUT(3) => 
                           IR_OUT_3_port, IR_OUT(2) => IR_OUT_2_port, IR_OUT(1)
                           => IR_OUT_1_port, IR_OUT(0) => IR_OUT_0_port, 
                           ADDERPC_OUT(31) => ADDERPC_OUTs_31_port, 
                           ADDERPC_OUT(30) => ADDERPC_OUTs_30_port, 
                           ADDERPC_OUT(29) => ADDERPC_OUTs_29_port, 
                           ADDERPC_OUT(28) => ADDERPC_OUTs_28_port, 
                           ADDERPC_OUT(27) => ADDERPC_OUTs_27_port, 
                           ADDERPC_OUT(26) => ADDERPC_OUTs_26_port, 
                           ADDERPC_OUT(25) => ADDERPC_OUTs_25_port, 
                           ADDERPC_OUT(24) => ADDERPC_OUTs_24_port, 
                           ADDERPC_OUT(23) => ADDERPC_OUTs_23_port, 
                           ADDERPC_OUT(22) => ADDERPC_OUTs_22_port, 
                           ADDERPC_OUT(21) => ADDERPC_OUTs_21_port, 
                           ADDERPC_OUT(20) => ADDERPC_OUTs_20_port, 
                           ADDERPC_OUT(19) => ADDERPC_OUTs_19_port, 
                           ADDERPC_OUT(18) => ADDERPC_OUTs_18_port, 
                           ADDERPC_OUT(17) => ADDERPC_OUTs_17_port, 
                           ADDERPC_OUT(16) => ADDERPC_OUTs_16_port, 
                           ADDERPC_OUT(15) => ADDERPC_OUTs_15_port, 
                           ADDERPC_OUT(14) => ADDERPC_OUTs_14_port, 
                           ADDERPC_OUT(13) => ADDERPC_OUTs_13_port, 
                           ADDERPC_OUT(12) => ADDERPC_OUTs_12_port, 
                           ADDERPC_OUT(11) => ADDERPC_OUTs_11_port, 
                           ADDERPC_OUT(10) => ADDERPC_OUTs_10_port, 
                           ADDERPC_OUT(9) => ADDERPC_OUTs_9_port, 
                           ADDERPC_OUT(8) => ADDERPC_OUTs_8_port, 
                           ADDERPC_OUT(7) => ADDERPC_OUTs_7_port, 
                           ADDERPC_OUT(6) => ADDERPC_OUTs_6_port, 
                           ADDERPC_OUT(5) => ADDERPC_OUTs_5_port, 
                           ADDERPC_OUT(4) => ADDERPC_OUTs_4_port, 
                           ADDERPC_OUT(3) => ADDERPC_OUTs_3_port, 
                           ADDERPC_OUT(2) => ADDERPC_OUTs_2_port, 
                           ADDERPC_OUT(1) => ADDERPC_OUTs_1_port, 
                           ADDERPC_OUT(0) => ADDERPC_OUTs_0_port);
   DECODE : decodeUnit_nbits32 port map( clk => n2, rst => n1, RegA_LATCH_EN =>
                           RegA_LATCH_EN, RegB_LATCH_EN => RegB_LATCH_EN, 
                           RegIMM_LATCH_EN => RegIMM_LATCH_EN, RF_WE => RF_WE, 
                           DATAIN(31) => DATAIN_RFs_31_port, DATAIN(30) => 
                           DATAIN_RFs_30_port, DATAIN(29) => DATAIN_RFs_29_port
                           , DATAIN(28) => DATAIN_RFs_28_port, DATAIN(27) => 
                           DATAIN_RFs_27_port, DATAIN(26) => DATAIN_RFs_26_port
                           , DATAIN(25) => DATAIN_RFs_25_port, DATAIN(24) => 
                           DATAIN_RFs_24_port, DATAIN(23) => DATAIN_RFs_23_port
                           , DATAIN(22) => DATAIN_RFs_22_port, DATAIN(21) => 
                           DATAIN_RFs_21_port, DATAIN(20) => DATAIN_RFs_20_port
                           , DATAIN(19) => DATAIN_RFs_19_port, DATAIN(18) => 
                           DATAIN_RFs_18_port, DATAIN(17) => DATAIN_RFs_17_port
                           , DATAIN(16) => DATAIN_RFs_16_port, DATAIN(15) => 
                           DATAIN_RFs_15_port, DATAIN(14) => DATAIN_RFs_14_port
                           , DATAIN(13) => DATAIN_RFs_13_port, DATAIN(12) => 
                           DATAIN_RFs_12_port, DATAIN(11) => DATAIN_RFs_11_port
                           , DATAIN(10) => DATAIN_RFs_10_port, DATAIN(9) => 
                           DATAIN_RFs_9_port, DATAIN(8) => DATAIN_RFs_8_port, 
                           DATAIN(7) => DATAIN_RFs_7_port, DATAIN(6) => 
                           DATAIN_RFs_6_port, DATAIN(5) => DATAIN_RFs_5_port, 
                           DATAIN(4) => DATAIN_RFs_4_port, DATAIN(3) => 
                           DATAIN_RFs_3_port, DATAIN(2) => DATAIN_RFs_2_port, 
                           DATAIN(1) => DATAIN_RFs_1_port, DATAIN(0) => 
                           DATAIN_RFs_0_port, IR_OUT(31) => IR_OUT_31_port, 
                           IR_OUT(30) => IR_OUT_30_port, IR_OUT(29) => 
                           IR_OUT_29_port, IR_OUT(28) => IR_OUT_28_port, 
                           IR_OUT(27) => IR_OUT_27_port, IR_OUT(26) => 
                           IR_OUT_26_port, IR_OUT(25) => IR_OUT_25_port, 
                           IR_OUT(24) => IR_OUT_24_port, IR_OUT(23) => 
                           IR_OUT_23_port, IR_OUT(22) => IR_OUT_22_port, 
                           IR_OUT(21) => IR_OUT_21_port, IR_OUT(20) => 
                           IR_OUT_20_port, IR_OUT(19) => IR_OUT_19_port, 
                           IR_OUT(18) => IR_OUT_18_port, IR_OUT(17) => 
                           IR_OUT_17_port, IR_OUT(16) => IR_OUT_16_port, 
                           IR_OUT(15) => IR_OUT_15_port, IR_OUT(14) => 
                           IR_OUT_14_port, IR_OUT(13) => IR_OUT_13_port, 
                           IR_OUT(12) => IR_OUT_12_port, IR_OUT(11) => 
                           IR_OUT_11_port, IR_OUT(10) => IR_OUT_10_port, 
                           IR_OUT(9) => IR_OUT_9_port, IR_OUT(8) => 
                           IR_OUT_8_port, IR_OUT(7) => IR_OUT_7_port, IR_OUT(6)
                           => IR_OUT_6_port, IR_OUT(5) => IR_OUT_5_port, 
                           IR_OUT(4) => IR_OUT_4_port, IR_OUT(3) => 
                           IR_OUT_3_port, IR_OUT(2) => IR_OUT_2_port, IR_OUT(1)
                           => IR_OUT_1_port, IR_OUT(0) => IR_OUT_0_port, 
                           A_out(31) => A_outs_31_port, A_out(30) => 
                           A_outs_30_port, A_out(29) => A_outs_29_port, 
                           A_out(28) => A_outs_28_port, A_out(27) => 
                           A_outs_27_port, A_out(26) => A_outs_26_port, 
                           A_out(25) => A_outs_25_port, A_out(24) => 
                           A_outs_24_port, A_out(23) => A_outs_23_port, 
                           A_out(22) => A_outs_22_port, A_out(21) => 
                           A_outs_21_port, A_out(20) => A_outs_20_port, 
                           A_out(19) => A_outs_19_port, A_out(18) => 
                           A_outs_18_port, A_out(17) => A_outs_17_port, 
                           A_out(16) => A_outs_16_port, A_out(15) => 
                           A_outs_15_port, A_out(14) => A_outs_14_port, 
                           A_out(13) => A_outs_13_port, A_out(12) => 
                           A_outs_12_port, A_out(11) => A_outs_11_port, 
                           A_out(10) => A_outs_10_port, A_out(9) => 
                           A_outs_9_port, A_out(8) => A_outs_8_port, A_out(7) 
                           => A_outs_7_port, A_out(6) => A_outs_6_port, 
                           A_out(5) => A_outs_5_port, A_out(4) => A_outs_4_port
                           , A_out(3) => A_outs_3_port, A_out(2) => 
                           A_outs_2_port, A_out(1) => A_outs_1_port, A_out(0) 
                           => A_outs_0_port, B_out(31) => B_outs_31_port, 
                           B_out(30) => B_outs_30_port, B_out(29) => 
                           B_outs_29_port, B_out(28) => B_outs_28_port, 
                           B_out(27) => B_outs_27_port, B_out(26) => 
                           B_outs_26_port, B_out(25) => B_outs_25_port, 
                           B_out(24) => B_outs_24_port, B_out(23) => 
                           B_outs_23_port, B_out(22) => B_outs_22_port, 
                           B_out(21) => B_outs_21_port, B_out(20) => 
                           B_outs_20_port, B_out(19) => B_outs_19_port, 
                           B_out(18) => B_outs_18_port, B_out(17) => 
                           B_outs_17_port, B_out(16) => B_outs_16_port, 
                           B_out(15) => B_outs_15_port, B_out(14) => 
                           B_outs_14_port, B_out(13) => B_outs_13_port, 
                           B_out(12) => B_outs_12_port, B_out(11) => 
                           B_outs_11_port, B_out(10) => B_outs_10_port, 
                           B_out(9) => B_outs_9_port, B_out(8) => B_outs_8_port
                           , B_out(7) => B_outs_7_port, B_out(6) => 
                           B_outs_6_port, B_out(5) => B_outs_5_port, B_out(4) 
                           => B_outs_4_port, B_out(3) => B_outs_3_port, 
                           B_out(2) => B_outs_2_port, B_out(1) => B_outs_1_port
                           , B_out(0) => B_outs_0_port, Imm_out(31) => 
                           Imm_outs_31_port, Imm_out(30) => Imm_outs_30_port, 
                           Imm_out(29) => Imm_outs_29_port, Imm_out(28) => 
                           Imm_outs_28_port, Imm_out(27) => Imm_outs_27_port, 
                           Imm_out(26) => Imm_outs_26_port, Imm_out(25) => 
                           Imm_outs_25_port, Imm_out(24) => Imm_outs_24_port, 
                           Imm_out(23) => Imm_outs_23_port, Imm_out(22) => 
                           Imm_outs_22_port, Imm_out(21) => Imm_outs_21_port, 
                           Imm_out(20) => Imm_outs_20_port, Imm_out(19) => 
                           Imm_outs_19_port, Imm_out(18) => Imm_outs_18_port, 
                           Imm_out(17) => Imm_outs_17_port, Imm_out(16) => 
                           Imm_outs_16_port, Imm_out(15) => Imm_outs_15_port, 
                           Imm_out(14) => Imm_outs_14_port, Imm_out(13) => 
                           Imm_outs_13_port, Imm_out(12) => Imm_outs_12_port, 
                           Imm_out(11) => Imm_outs_11_port, Imm_out(10) => 
                           Imm_outs_10_port, Imm_out(9) => Imm_outs_9_port, 
                           Imm_out(8) => Imm_outs_8_port, Imm_out(7) => 
                           Imm_outs_7_port, Imm_out(6) => Imm_outs_6_port, 
                           Imm_out(5) => Imm_outs_5_port, Imm_out(4) => 
                           Imm_outs_4_port, Imm_out(3) => Imm_outs_3_port, 
                           Imm_out(2) => Imm_outs_2_port, Imm_out(1) => 
                           Imm_outs_1_port, Imm_out(0) => Imm_outs_0_port, 
                           IR_IN2(31) => IR_OUT4s_31_port, IR_IN2(30) => 
                           IR_OUT4s_30_port, IR_IN2(29) => IR_OUT4s_29_port, 
                           IR_IN2(28) => IR_OUT4s_28_port, IR_IN2(27) => 
                           IR_OUT4s_27_port, IR_IN2(26) => IR_OUT4s_26_port, 
                           IR_IN2(25) => IR_OUT4s_25_port, IR_IN2(24) => 
                           IR_OUT4s_24_port, IR_IN2(23) => IR_OUT4s_23_port, 
                           IR_IN2(22) => IR_OUT4s_22_port, IR_IN2(21) => 
                           IR_OUT4s_21_port, IR_IN2(20) => IR_OUT4s_20_port, 
                           IR_IN2(19) => IR_OUT4s_19_port, IR_IN2(18) => 
                           IR_OUT4s_18_port, IR_IN2(17) => IR_OUT4s_17_port, 
                           IR_IN2(16) => IR_OUT4s_16_port, IR_IN2(15) => 
                           IR_OUT4s_15_port, IR_IN2(14) => IR_OUT4s_14_port, 
                           IR_IN2(13) => IR_OUT4s_13_port, IR_IN2(12) => 
                           IR_OUT4s_12_port, IR_IN2(11) => IR_OUT4s_11_port, 
                           IR_IN2(10) => IR_OUT4s_10_port, IR_IN2(9) => 
                           IR_OUT4s_9_port, IR_IN2(8) => IR_OUT4s_8_port, 
                           IR_IN2(7) => IR_OUT4s_7_port, IR_IN2(6) => 
                           IR_OUT4s_6_port, IR_IN2(5) => IR_OUT4s_5_port, 
                           IR_IN2(4) => IR_OUT4s_4_port, IR_IN2(3) => 
                           IR_OUT4s_3_port, IR_IN2(2) => IR_OUT4s_2_port, 
                           IR_IN2(1) => IR_OUT4s_1_port, IR_IN2(0) => 
                           IR_OUT4s_0_port, IR_OUT2(31) => IR_OUT2s_31_port, 
                           IR_OUT2(30) => IR_OUT2s_30_port, IR_OUT2(29) => 
                           IR_OUT2s_29_port, IR_OUT2(28) => IR_OUT2s_28_port, 
                           IR_OUT2(27) => IR_OUT2s_27_port, IR_OUT2(26) => 
                           IR_OUT2s_26_port, IR_OUT2(25) => IR_OUT2s_25_port, 
                           IR_OUT2(24) => IR_OUT2s_24_port, IR_OUT2(23) => 
                           IR_OUT2s_23_port, IR_OUT2(22) => IR_OUT2s_22_port, 
                           IR_OUT2(21) => IR_OUT2s_21_port, IR_OUT2(20) => 
                           IR_OUT2s_20_port, IR_OUT2(19) => IR_OUT2s_19_port, 
                           IR_OUT2(18) => IR_OUT2s_18_port, IR_OUT2(17) => 
                           IR_OUT2s_17_port, IR_OUT2(16) => IR_OUT2s_16_port, 
                           IR_OUT2(15) => IR_OUT2s_15_port, IR_OUT2(14) => 
                           IR_OUT2s_14_port, IR_OUT2(13) => IR_OUT2s_13_port, 
                           IR_OUT2(12) => IR_OUT2s_12_port, IR_OUT2(11) => 
                           IR_OUT2s_11_port, IR_OUT2(10) => IR_OUT2s_10_port, 
                           IR_OUT2(9) => IR_OUT2s_9_port, IR_OUT2(8) => 
                           IR_OUT2s_8_port, IR_OUT2(7) => IR_OUT2s_7_port, 
                           IR_OUT2(6) => IR_OUT2s_6_port, IR_OUT2(5) => 
                           IR_OUT2s_5_port, IR_OUT2(4) => IR_OUT2s_4_port, 
                           IR_OUT2(3) => IR_OUT2s_3_port, IR_OUT2(2) => 
                           IR_OUT2s_2_port, IR_OUT2(1) => IR_OUT2s_1_port, 
                           IR_OUT2(0) => IR_OUT2s_0_port, NPC_IN(31) => 
                           NPC_OUTs_31_port, NPC_IN(30) => NPC_OUTs_30_port, 
                           NPC_IN(29) => NPC_OUTs_29_port, NPC_IN(28) => 
                           NPC_OUTs_28_port, NPC_IN(27) => NPC_OUTs_27_port, 
                           NPC_IN(26) => NPC_OUTs_26_port, NPC_IN(25) => 
                           NPC_OUTs_25_port, NPC_IN(24) => NPC_OUTs_24_port, 
                           NPC_IN(23) => NPC_OUTs_23_port, NPC_IN(22) => 
                           NPC_OUTs_22_port, NPC_IN(21) => NPC_OUTs_21_port, 
                           NPC_IN(20) => NPC_OUTs_20_port, NPC_IN(19) => 
                           NPC_OUTs_19_port, NPC_IN(18) => NPC_OUTs_18_port, 
                           NPC_IN(17) => NPC_OUTs_17_port, NPC_IN(16) => 
                           NPC_OUTs_16_port, NPC_IN(15) => NPC_OUTs_15_port, 
                           NPC_IN(14) => NPC_OUTs_14_port, NPC_IN(13) => 
                           NPC_OUTs_13_port, NPC_IN(12) => NPC_OUTs_12_port, 
                           NPC_IN(11) => NPC_OUTs_11_port, NPC_IN(10) => 
                           NPC_OUTs_10_port, NPC_IN(9) => NPC_OUTs_9_port, 
                           NPC_IN(8) => NPC_OUTs_8_port, NPC_IN(7) => 
                           NPC_OUTs_7_port, NPC_IN(6) => NPC_OUTs_6_port, 
                           NPC_IN(5) => NPC_OUTs_5_port, NPC_IN(4) => 
                           NPC_OUTs_4_port, NPC_IN(3) => NPC_OUTs_3_port, 
                           NPC_IN(2) => NPC_OUTs_2_port, NPC_IN(1) => 
                           NPC_OUTs_1_port, NPC_IN(0) => NPC_OUTs_0_port, 
                           NPC2_OUT(31) => NPC2_OUTs_31_port, NPC2_OUT(30) => 
                           NPC2_OUTs_30_port, NPC2_OUT(29) => NPC2_OUTs_29_port
                           , NPC2_OUT(28) => NPC2_OUTs_28_port, NPC2_OUT(27) =>
                           NPC2_OUTs_27_port, NPC2_OUT(26) => NPC2_OUTs_26_port
                           , NPC2_OUT(25) => NPC2_OUTs_25_port, NPC2_OUT(24) =>
                           NPC2_OUTs_24_port, NPC2_OUT(23) => NPC2_OUTs_23_port
                           , NPC2_OUT(22) => NPC2_OUTs_22_port, NPC2_OUT(21) =>
                           NPC2_OUTs_21_port, NPC2_OUT(20) => NPC2_OUTs_20_port
                           , NPC2_OUT(19) => NPC2_OUTs_19_port, NPC2_OUT(18) =>
                           NPC2_OUTs_18_port, NPC2_OUT(17) => NPC2_OUTs_17_port
                           , NPC2_OUT(16) => NPC2_OUTs_16_port, NPC2_OUT(15) =>
                           NPC2_OUTs_15_port, NPC2_OUT(14) => NPC2_OUTs_14_port
                           , NPC2_OUT(13) => NPC2_OUTs_13_port, NPC2_OUT(12) =>
                           NPC2_OUTs_12_port, NPC2_OUT(11) => NPC2_OUTs_11_port
                           , NPC2_OUT(10) => NPC2_OUTs_10_port, NPC2_OUT(9) => 
                           NPC2_OUTs_9_port, NPC2_OUT(8) => NPC2_OUTs_8_port, 
                           NPC2_OUT(7) => NPC2_OUTs_7_port, NPC2_OUT(6) => 
                           NPC2_OUTs_6_port, NPC2_OUT(5) => NPC2_OUTs_5_port, 
                           NPC2_OUT(4) => NPC2_OUTs_4_port, NPC2_OUT(3) => 
                           NPC2_OUTs_3_port, NPC2_OUT(2) => NPC2_OUTs_2_port, 
                           NPC2_OUT(1) => NPC2_OUTs_1_port, NPC2_OUT(0) => 
                           NPC2_OUTs_0_port);
   EXECUTE : executionUnit_nbits32 port map( clk => n2, rst => n1, 
                           ALU_OUTREG_ENABLE => ALU_OUTREG_EN, MUXA_SEL => 
                           MUXA_SEL, MUXB_SEL => MUXB_SEL, COND_ENABLE => 
                           EQ_COND, ALU_BITS(0) => ALU_OPCODE(0), ALU_BITS(1) 
                           => ALU_OPCODE(1), ALU_BITS(2) => ALU_OPCODE(2), 
                           ALU_BITS(3) => ALU_OPCODE(3), NPC_OUT(31) => 
                           NPC2_OUTs_31_port, NPC_OUT(30) => NPC2_OUTs_30_port,
                           NPC_OUT(29) => NPC2_OUTs_29_port, NPC_OUT(28) => 
                           NPC2_OUTs_28_port, NPC_OUT(27) => NPC2_OUTs_27_port,
                           NPC_OUT(26) => NPC2_OUTs_26_port, NPC_OUT(25) => 
                           NPC2_OUTs_25_port, NPC_OUT(24) => NPC2_OUTs_24_port,
                           NPC_OUT(23) => NPC2_OUTs_23_port, NPC_OUT(22) => 
                           NPC2_OUTs_22_port, NPC_OUT(21) => NPC2_OUTs_21_port,
                           NPC_OUT(20) => NPC2_OUTs_20_port, NPC_OUT(19) => 
                           NPC2_OUTs_19_port, NPC_OUT(18) => NPC2_OUTs_18_port,
                           NPC_OUT(17) => NPC2_OUTs_17_port, NPC_OUT(16) => 
                           NPC2_OUTs_16_port, NPC_OUT(15) => NPC2_OUTs_15_port,
                           NPC_OUT(14) => NPC2_OUTs_14_port, NPC_OUT(13) => 
                           NPC2_OUTs_13_port, NPC_OUT(12) => NPC2_OUTs_12_port,
                           NPC_OUT(11) => NPC2_OUTs_11_port, NPC_OUT(10) => 
                           NPC2_OUTs_10_port, NPC_OUT(9) => NPC2_OUTs_9_port, 
                           NPC_OUT(8) => NPC2_OUTs_8_port, NPC_OUT(7) => 
                           NPC2_OUTs_7_port, NPC_OUT(6) => NPC2_OUTs_6_port, 
                           NPC_OUT(5) => NPC2_OUTs_5_port, NPC_OUT(4) => 
                           NPC2_OUTs_4_port, NPC_OUT(3) => NPC2_OUTs_3_port, 
                           NPC_OUT(2) => NPC2_OUTs_2_port, NPC_OUT(1) => 
                           NPC2_OUTs_1_port, NPC_OUT(0) => NPC2_OUTs_0_port, 
                           A_out(31) => A_outs_31_port, A_out(30) => 
                           A_outs_30_port, A_out(29) => A_outs_29_port, 
                           A_out(28) => A_outs_28_port, A_out(27) => 
                           A_outs_27_port, A_out(26) => A_outs_26_port, 
                           A_out(25) => A_outs_25_port, A_out(24) => 
                           A_outs_24_port, A_out(23) => A_outs_23_port, 
                           A_out(22) => A_outs_22_port, A_out(21) => 
                           A_outs_21_port, A_out(20) => A_outs_20_port, 
                           A_out(19) => A_outs_19_port, A_out(18) => 
                           A_outs_18_port, A_out(17) => A_outs_17_port, 
                           A_out(16) => A_outs_16_port, A_out(15) => 
                           A_outs_15_port, A_out(14) => A_outs_14_port, 
                           A_out(13) => A_outs_13_port, A_out(12) => 
                           A_outs_12_port, A_out(11) => A_outs_11_port, 
                           A_out(10) => A_outs_10_port, A_out(9) => 
                           A_outs_9_port, A_out(8) => A_outs_8_port, A_out(7) 
                           => A_outs_7_port, A_out(6) => A_outs_6_port, 
                           A_out(5) => A_outs_5_port, A_out(4) => A_outs_4_port
                           , A_out(3) => A_outs_3_port, A_out(2) => 
                           A_outs_2_port, A_out(1) => A_outs_1_port, A_out(0) 
                           => A_outs_0_port, B_out(31) => B_outs_31_port, 
                           B_out(30) => B_outs_30_port, B_out(29) => 
                           B_outs_29_port, B_out(28) => B_outs_28_port, 
                           B_out(27) => B_outs_27_port, B_out(26) => 
                           B_outs_26_port, B_out(25) => B_outs_25_port, 
                           B_out(24) => B_outs_24_port, B_out(23) => 
                           B_outs_23_port, B_out(22) => B_outs_22_port, 
                           B_out(21) => B_outs_21_port, B_out(20) => 
                           B_outs_20_port, B_out(19) => B_outs_19_port, 
                           B_out(18) => B_outs_18_port, B_out(17) => 
                           B_outs_17_port, B_out(16) => B_outs_16_port, 
                           B_out(15) => B_outs_15_port, B_out(14) => 
                           B_outs_14_port, B_out(13) => B_outs_13_port, 
                           B_out(12) => B_outs_12_port, B_out(11) => 
                           B_outs_11_port, B_out(10) => B_outs_10_port, 
                           B_out(9) => B_outs_9_port, B_out(8) => B_outs_8_port
                           , B_out(7) => B_outs_7_port, B_out(6) => 
                           B_outs_6_port, B_out(5) => B_outs_5_port, B_out(4) 
                           => B_outs_4_port, B_out(3) => B_outs_3_port, 
                           B_out(2) => B_outs_2_port, B_out(1) => B_outs_1_port
                           , B_out(0) => B_outs_0_port, Imm_out(31) => 
                           Imm_outs_31_port, Imm_out(30) => Imm_outs_30_port, 
                           Imm_out(29) => Imm_outs_29_port, Imm_out(28) => 
                           Imm_outs_28_port, Imm_out(27) => Imm_outs_27_port, 
                           Imm_out(26) => Imm_outs_26_port, Imm_out(25) => 
                           Imm_outs_25_port, Imm_out(24) => Imm_outs_24_port, 
                           Imm_out(23) => Imm_outs_23_port, Imm_out(22) => 
                           Imm_outs_22_port, Imm_out(21) => Imm_outs_21_port, 
                           Imm_out(20) => Imm_outs_20_port, Imm_out(19) => 
                           Imm_outs_19_port, Imm_out(18) => Imm_outs_18_port, 
                           Imm_out(17) => Imm_outs_17_port, Imm_out(16) => 
                           Imm_outs_16_port, Imm_out(15) => Imm_outs_15_port, 
                           Imm_out(14) => Imm_outs_14_port, Imm_out(13) => 
                           Imm_outs_13_port, Imm_out(12) => Imm_outs_12_port, 
                           Imm_out(11) => Imm_outs_11_port, Imm_out(10) => 
                           Imm_outs_10_port, Imm_out(9) => Imm_outs_9_port, 
                           Imm_out(8) => Imm_outs_8_port, Imm_out(7) => 
                           Imm_outs_7_port, Imm_out(6) => Imm_outs_6_port, 
                           Imm_out(5) => Imm_outs_5_port, Imm_out(4) => 
                           Imm_outs_4_port, Imm_out(3) => Imm_outs_3_port, 
                           Imm_out(2) => Imm_outs_2_port, Imm_out(1) => 
                           Imm_outs_1_port, Imm_out(0) => Imm_outs_0_port, 
                           ALUREG_OUTPUT(31) => ALU_OUT_31_port, 
                           ALUREG_OUTPUT(30) => ALU_OUT_30_port, 
                           ALUREG_OUTPUT(29) => ALU_OUT_29_port, 
                           ALUREG_OUTPUT(28) => ALU_OUT_28_port, 
                           ALUREG_OUTPUT(27) => ALU_OUT_27_port, 
                           ALUREG_OUTPUT(26) => ALU_OUT_26_port, 
                           ALUREG_OUTPUT(25) => ALU_OUT_25_port, 
                           ALUREG_OUTPUT(24) => ALU_OUT_24_port, 
                           ALUREG_OUTPUT(23) => ALU_OUT_23_port, 
                           ALUREG_OUTPUT(22) => ALU_OUT_22_port, 
                           ALUREG_OUTPUT(21) => ALU_OUT_21_port, 
                           ALUREG_OUTPUT(20) => ALU_OUT_20_port, 
                           ALUREG_OUTPUT(19) => ALU_OUT_19_port, 
                           ALUREG_OUTPUT(18) => ALU_OUT_18_port, 
                           ALUREG_OUTPUT(17) => ALU_OUT_17_port, 
                           ALUREG_OUTPUT(16) => ALU_OUT_16_port, 
                           ALUREG_OUTPUT(15) => ALU_OUT_15_port, 
                           ALUREG_OUTPUT(14) => ALU_OUT_14_port, 
                           ALUREG_OUTPUT(13) => ALU_OUT_13_port, 
                           ALUREG_OUTPUT(12) => ALU_OUT_12_port, 
                           ALUREG_OUTPUT(11) => ALU_OUT_11_port, 
                           ALUREG_OUTPUT(10) => ALU_OUT_10_port, 
                           ALUREG_OUTPUT(9) => ALU_OUT_9_port, ALUREG_OUTPUT(8)
                           => ALU_OUT_8_port, ALUREG_OUTPUT(7) => 
                           ALU_OUT_7_port, ALUREG_OUTPUT(6) => ALU_OUT_6_port, 
                           ALUREG_OUTPUT(5) => ALU_OUT_5_port, ALUREG_OUTPUT(4)
                           => ALU_OUT_4_port, ALUREG_OUTPUT(3) => 
                           ALU_OUT_3_port, ALUREG_OUTPUT(2) => ALU_OUT_2_port, 
                           ALUREG_OUTPUT(1) => ALU_OUT_1_port, ALUREG_OUTPUT(0)
                           => ALU_OUT_0_port, COND_OUT => COND_OUTs, IR_IN3(31)
                           => IR_OUT2s_31_port, IR_IN3(30) => IR_OUT2s_30_port,
                           IR_IN3(29) => IR_OUT2s_29_port, IR_IN3(28) => 
                           IR_OUT2s_28_port, IR_IN3(27) => IR_OUT2s_27_port, 
                           IR_IN3(26) => IR_OUT2s_26_port, IR_IN3(25) => 
                           IR_OUT2s_25_port, IR_IN3(24) => IR_OUT2s_24_port, 
                           IR_IN3(23) => IR_OUT2s_23_port, IR_IN3(22) => 
                           IR_OUT2s_22_port, IR_IN3(21) => IR_OUT2s_21_port, 
                           IR_IN3(20) => IR_OUT2s_20_port, IR_IN3(19) => 
                           IR_OUT2s_19_port, IR_IN3(18) => IR_OUT2s_18_port, 
                           IR_IN3(17) => IR_OUT2s_17_port, IR_IN3(16) => 
                           IR_OUT2s_16_port, IR_IN3(15) => IR_OUT2s_15_port, 
                           IR_IN3(14) => IR_OUT2s_14_port, IR_IN3(13) => 
                           IR_OUT2s_13_port, IR_IN3(12) => IR_OUT2s_12_port, 
                           IR_IN3(11) => IR_OUT2s_11_port, IR_IN3(10) => 
                           IR_OUT2s_10_port, IR_IN3(9) => IR_OUT2s_9_port, 
                           IR_IN3(8) => IR_OUT2s_8_port, IR_IN3(7) => 
                           IR_OUT2s_7_port, IR_IN3(6) => IR_OUT2s_6_port, 
                           IR_IN3(5) => IR_OUT2s_5_port, IR_IN3(4) => 
                           IR_OUT2s_4_port, IR_IN3(3) => IR_OUT2s_3_port, 
                           IR_IN3(2) => IR_OUT2s_2_port, IR_IN3(1) => 
                           IR_OUT2s_1_port, IR_IN3(0) => IR_OUT2s_0_port, 
                           IR_OUT3(31) => IR_OUT3s_31_port, IR_OUT3(30) => 
                           IR_OUT3s_30_port, IR_OUT3(29) => IR_OUT3s_29_port, 
                           IR_OUT3(28) => IR_OUT3s_28_port, IR_OUT3(27) => 
                           IR_OUT3s_27_port, IR_OUT3(26) => IR_OUT3s_26_port, 
                           IR_OUT3(25) => IR_OUT3s_25_port, IR_OUT3(24) => 
                           IR_OUT3s_24_port, IR_OUT3(23) => IR_OUT3s_23_port, 
                           IR_OUT3(22) => IR_OUT3s_22_port, IR_OUT3(21) => 
                           IR_OUT3s_21_port, IR_OUT3(20) => IR_OUT3s_20_port, 
                           IR_OUT3(19) => IR_OUT3s_19_port, IR_OUT3(18) => 
                           IR_OUT3s_18_port, IR_OUT3(17) => IR_OUT3s_17_port, 
                           IR_OUT3(16) => IR_OUT3s_16_port, IR_OUT3(15) => 
                           IR_OUT3s_15_port, IR_OUT3(14) => IR_OUT3s_14_port, 
                           IR_OUT3(13) => IR_OUT3s_13_port, IR_OUT3(12) => 
                           IR_OUT3s_12_port, IR_OUT3(11) => IR_OUT3s_11_port, 
                           IR_OUT3(10) => IR_OUT3s_10_port, IR_OUT3(9) => 
                           IR_OUT3s_9_port, IR_OUT3(8) => IR_OUT3s_8_port, 
                           IR_OUT3(7) => IR_OUT3s_7_port, IR_OUT3(6) => 
                           IR_OUT3s_6_port, IR_OUT3(5) => IR_OUT3s_5_port, 
                           IR_OUT3(4) => IR_OUT3s_4_port, IR_OUT3(3) => 
                           IR_OUT3s_3_port, IR_OUT3(2) => IR_OUT3s_2_port, 
                           IR_OUT3(1) => IR_OUT3s_1_port, IR_OUT3(0) => 
                           IR_OUT3s_0_port, B_outreg(31) => B(31), B_outreg(30)
                           => B(30), B_outreg(29) => B(29), B_outreg(28) => 
                           B(28), B_outreg(27) => B(27), B_outreg(26) => B(26),
                           B_outreg(25) => B(25), B_outreg(24) => B(24), 
                           B_outreg(23) => B(23), B_outreg(22) => B(22), 
                           B_outreg(21) => B(21), B_outreg(20) => B(20), 
                           B_outreg(19) => B(19), B_outreg(18) => B(18), 
                           B_outreg(17) => B(17), B_outreg(16) => B(16), 
                           B_outreg(15) => B(15), B_outreg(14) => B(14), 
                           B_outreg(13) => B(13), B_outreg(12) => B(12), 
                           B_outreg(11) => B(11), B_outreg(10) => B(10), 
                           B_outreg(9) => B(9), B_outreg(8) => B(8), 
                           B_outreg(7) => B(7), B_outreg(6) => B(6), 
                           B_outreg(5) => B(5), B_outreg(4) => B(4), 
                           B_outreg(3) => B(3), B_outreg(2) => B(2), 
                           B_outreg(1) => B(1), B_outreg(0) => B(0));
   MEMORY : memoryUnit_nbits32 port map( clk => n2, rst => n1, LMD_LATCH_EN => 
                           LMD_LATCH_EN, JUMP_EN => JUMP_EN, DRAM_DATA(31) => 
                           DRAM_DATA(31), DRAM_DATA(30) => DRAM_DATA(30), 
                           DRAM_DATA(29) => DRAM_DATA(29), DRAM_DATA(28) => 
                           DRAM_DATA(28), DRAM_DATA(27) => DRAM_DATA(27), 
                           DRAM_DATA(26) => DRAM_DATA(26), DRAM_DATA(25) => 
                           DRAM_DATA(25), DRAM_DATA(24) => DRAM_DATA(24), 
                           DRAM_DATA(23) => DRAM_DATA(23), DRAM_DATA(22) => 
                           DRAM_DATA(22), DRAM_DATA(21) => DRAM_DATA(21), 
                           DRAM_DATA(20) => DRAM_DATA(20), DRAM_DATA(19) => 
                           DRAM_DATA(19), DRAM_DATA(18) => DRAM_DATA(18), 
                           DRAM_DATA(17) => DRAM_DATA(17), DRAM_DATA(16) => 
                           DRAM_DATA(16), DRAM_DATA(15) => DRAM_DATA(15), 
                           DRAM_DATA(14) => DRAM_DATA(14), DRAM_DATA(13) => 
                           DRAM_DATA(13), DRAM_DATA(12) => DRAM_DATA(12), 
                           DRAM_DATA(11) => DRAM_DATA(11), DRAM_DATA(10) => 
                           DRAM_DATA(10), DRAM_DATA(9) => DRAM_DATA(9), 
                           DRAM_DATA(8) => DRAM_DATA(8), DRAM_DATA(7) => 
                           DRAM_DATA(7), DRAM_DATA(6) => DRAM_DATA(6), 
                           DRAM_DATA(5) => DRAM_DATA(5), DRAM_DATA(4) => 
                           DRAM_DATA(4), DRAM_DATA(3) => DRAM_DATA(3), 
                           DRAM_DATA(2) => DRAM_DATA(2), DRAM_DATA(1) => 
                           DRAM_DATA(1), DRAM_DATA(0) => DRAM_DATA(0), 
                           ALUREG_OUTPUT(31) => ALU_OUT_31_port, 
                           ALUREG_OUTPUT(30) => ALU_OUT_30_port, 
                           ALUREG_OUTPUT(29) => ALU_OUT_29_port, 
                           ALUREG_OUTPUT(28) => ALU_OUT_28_port, 
                           ALUREG_OUTPUT(27) => ALU_OUT_27_port, 
                           ALUREG_OUTPUT(26) => ALU_OUT_26_port, 
                           ALUREG_OUTPUT(25) => ALU_OUT_25_port, 
                           ALUREG_OUTPUT(24) => ALU_OUT_24_port, 
                           ALUREG_OUTPUT(23) => ALU_OUT_23_port, 
                           ALUREG_OUTPUT(22) => ALU_OUT_22_port, 
                           ALUREG_OUTPUT(21) => ALU_OUT_21_port, 
                           ALUREG_OUTPUT(20) => ALU_OUT_20_port, 
                           ALUREG_OUTPUT(19) => ALU_OUT_19_port, 
                           ALUREG_OUTPUT(18) => ALU_OUT_18_port, 
                           ALUREG_OUTPUT(17) => ALU_OUT_17_port, 
                           ALUREG_OUTPUT(16) => ALU_OUT_16_port, 
                           ALUREG_OUTPUT(15) => ALU_OUT_15_port, 
                           ALUREG_OUTPUT(14) => ALU_OUT_14_port, 
                           ALUREG_OUTPUT(13) => ALU_OUT_13_port, 
                           ALUREG_OUTPUT(12) => ALU_OUT_12_port, 
                           ALUREG_OUTPUT(11) => ALU_OUT_11_port, 
                           ALUREG_OUTPUT(10) => ALU_OUT_10_port, 
                           ALUREG_OUTPUT(9) => ALU_OUT_9_port, ALUREG_OUTPUT(8)
                           => ALU_OUT_8_port, ALUREG_OUTPUT(7) => 
                           ALU_OUT_7_port, ALUREG_OUTPUT(6) => ALU_OUT_6_port, 
                           ALUREG_OUTPUT(5) => ALU_OUT_5_port, ALUREG_OUTPUT(4)
                           => ALU_OUT_4_port, ALUREG_OUTPUT(3) => 
                           ALU_OUT_3_port, ALUREG_OUTPUT(2) => ALU_OUT_2_port, 
                           ALUREG_OUTPUT(1) => ALU_OUT_1_port, ALUREG_OUTPUT(0)
                           => ALU_OUT_0_port, NPC_OUT(31) => 
                           ADDERPC_OUTs_31_port, NPC_OUT(30) => 
                           ADDERPC_OUTs_30_port, NPC_OUT(29) => 
                           ADDERPC_OUTs_29_port, NPC_OUT(28) => 
                           ADDERPC_OUTs_28_port, NPC_OUT(27) => 
                           ADDERPC_OUTs_27_port, NPC_OUT(26) => 
                           ADDERPC_OUTs_26_port, NPC_OUT(25) => 
                           ADDERPC_OUTs_25_port, NPC_OUT(24) => 
                           ADDERPC_OUTs_24_port, NPC_OUT(23) => 
                           ADDERPC_OUTs_23_port, NPC_OUT(22) => 
                           ADDERPC_OUTs_22_port, NPC_OUT(21) => 
                           ADDERPC_OUTs_21_port, NPC_OUT(20) => 
                           ADDERPC_OUTs_20_port, NPC_OUT(19) => 
                           ADDERPC_OUTs_19_port, NPC_OUT(18) => 
                           ADDERPC_OUTs_18_port, NPC_OUT(17) => 
                           ADDERPC_OUTs_17_port, NPC_OUT(16) => 
                           ADDERPC_OUTs_16_port, NPC_OUT(15) => 
                           ADDERPC_OUTs_15_port, NPC_OUT(14) => 
                           ADDERPC_OUTs_14_port, NPC_OUT(13) => 
                           ADDERPC_OUTs_13_port, NPC_OUT(12) => 
                           ADDERPC_OUTs_12_port, NPC_OUT(11) => 
                           ADDERPC_OUTs_11_port, NPC_OUT(10) => 
                           ADDERPC_OUTs_10_port, NPC_OUT(9) => 
                           ADDERPC_OUTs_9_port, NPC_OUT(8) => 
                           ADDERPC_OUTs_8_port, NPC_OUT(7) => 
                           ADDERPC_OUTs_7_port, NPC_OUT(6) => 
                           ADDERPC_OUTs_6_port, NPC_OUT(5) => 
                           ADDERPC_OUTs_5_port, NPC_OUT(4) => 
                           ADDERPC_OUTs_4_port, NPC_OUT(3) => 
                           ADDERPC_OUTs_3_port, NPC_OUT(2) => 
                           ADDERPC_OUTs_2_port, NPC_OUT(1) => 
                           ADDERPC_OUTs_1_port, NPC_OUT(0) => 
                           ADDERPC_OUTs_0_port, COND_OUT => COND_OUTs, 
                           DRAM_DATAout(31) => LMD_OUTs_31_port, 
                           DRAM_DATAout(30) => LMD_OUTs_30_port, 
                           DRAM_DATAout(29) => LMD_OUTs_29_port, 
                           DRAM_DATAout(28) => LMD_OUTs_28_port, 
                           DRAM_DATAout(27) => LMD_OUTs_27_port, 
                           DRAM_DATAout(26) => LMD_OUTs_26_port, 
                           DRAM_DATAout(25) => LMD_OUTs_25_port, 
                           DRAM_DATAout(24) => LMD_OUTs_24_port, 
                           DRAM_DATAout(23) => LMD_OUTs_23_port, 
                           DRAM_DATAout(22) => LMD_OUTs_22_port, 
                           DRAM_DATAout(21) => LMD_OUTs_21_port, 
                           DRAM_DATAout(20) => LMD_OUTs_20_port, 
                           DRAM_DATAout(19) => LMD_OUTs_19_port, 
                           DRAM_DATAout(18) => LMD_OUTs_18_port, 
                           DRAM_DATAout(17) => LMD_OUTs_17_port, 
                           DRAM_DATAout(16) => LMD_OUTs_16_port, 
                           DRAM_DATAout(15) => LMD_OUTs_15_port, 
                           DRAM_DATAout(14) => LMD_OUTs_14_port, 
                           DRAM_DATAout(13) => LMD_OUTs_13_port, 
                           DRAM_DATAout(12) => LMD_OUTs_12_port, 
                           DRAM_DATAout(11) => LMD_OUTs_11_port, 
                           DRAM_DATAout(10) => LMD_OUTs_10_port, 
                           DRAM_DATAout(9) => LMD_OUTs_9_port, DRAM_DATAout(8) 
                           => LMD_OUTs_8_port, DRAM_DATAout(7) => 
                           LMD_OUTs_7_port, DRAM_DATAout(6) => LMD_OUTs_6_port,
                           DRAM_DATAout(5) => LMD_OUTs_5_port, DRAM_DATAout(4) 
                           => LMD_OUTs_4_port, DRAM_DATAout(3) => 
                           LMD_OUTs_3_port, DRAM_DATAout(2) => LMD_OUTs_2_port,
                           DRAM_DATAout(1) => LMD_OUTs_1_port, DRAM_DATAout(0) 
                           => LMD_OUTs_0_port, TO_PC_OUT(31) => 
                           TO_PC_OUTs_31_port, TO_PC_OUT(30) => 
                           TO_PC_OUTs_30_port, TO_PC_OUT(29) => 
                           TO_PC_OUTs_29_port, TO_PC_OUT(28) => 
                           TO_PC_OUTs_28_port, TO_PC_OUT(27) => 
                           TO_PC_OUTs_27_port, TO_PC_OUT(26) => 
                           TO_PC_OUTs_26_port, TO_PC_OUT(25) => 
                           TO_PC_OUTs_25_port, TO_PC_OUT(24) => 
                           TO_PC_OUTs_24_port, TO_PC_OUT(23) => 
                           TO_PC_OUTs_23_port, TO_PC_OUT(22) => 
                           TO_PC_OUTs_22_port, TO_PC_OUT(21) => 
                           TO_PC_OUTs_21_port, TO_PC_OUT(20) => 
                           TO_PC_OUTs_20_port, TO_PC_OUT(19) => 
                           TO_PC_OUTs_19_port, TO_PC_OUT(18) => 
                           TO_PC_OUTs_18_port, TO_PC_OUT(17) => 
                           TO_PC_OUTs_17_port, TO_PC_OUT(16) => 
                           TO_PC_OUTs_16_port, TO_PC_OUT(15) => 
                           TO_PC_OUTs_15_port, TO_PC_OUT(14) => 
                           TO_PC_OUTs_14_port, TO_PC_OUT(13) => 
                           TO_PC_OUTs_13_port, TO_PC_OUT(12) => 
                           TO_PC_OUTs_12_port, TO_PC_OUT(11) => 
                           TO_PC_OUTs_11_port, TO_PC_OUT(10) => 
                           TO_PC_OUTs_10_port, TO_PC_OUT(9) => 
                           TO_PC_OUTs_9_port, TO_PC_OUT(8) => TO_PC_OUTs_8_port
                           , TO_PC_OUT(7) => TO_PC_OUTs_7_port, TO_PC_OUT(6) =>
                           TO_PC_OUTs_6_port, TO_PC_OUT(5) => TO_PC_OUTs_5_port
                           , TO_PC_OUT(4) => TO_PC_OUTs_4_port, TO_PC_OUT(3) =>
                           TO_PC_OUTs_3_port, TO_PC_OUT(2) => TO_PC_OUTs_2_port
                           , TO_PC_OUT(1) => TO_PC_OUTs_1_port, TO_PC_OUT(0) =>
                           TO_PC_OUTs_0_port, ALU_OUT2(31) => ALU_OUT2s_31_port
                           , ALU_OUT2(30) => ALU_OUT2s_30_port, ALU_OUT2(29) =>
                           ALU_OUT2s_29_port, ALU_OUT2(28) => ALU_OUT2s_28_port
                           , ALU_OUT2(27) => ALU_OUT2s_27_port, ALU_OUT2(26) =>
                           ALU_OUT2s_26_port, ALU_OUT2(25) => ALU_OUT2s_25_port
                           , ALU_OUT2(24) => ALU_OUT2s_24_port, ALU_OUT2(23) =>
                           ALU_OUT2s_23_port, ALU_OUT2(22) => ALU_OUT2s_22_port
                           , ALU_OUT2(21) => ALU_OUT2s_21_port, ALU_OUT2(20) =>
                           ALU_OUT2s_20_port, ALU_OUT2(19) => ALU_OUT2s_19_port
                           , ALU_OUT2(18) => ALU_OUT2s_18_port, ALU_OUT2(17) =>
                           ALU_OUT2s_17_port, ALU_OUT2(16) => ALU_OUT2s_16_port
                           , ALU_OUT2(15) => ALU_OUT2s_15_port, ALU_OUT2(14) =>
                           ALU_OUT2s_14_port, ALU_OUT2(13) => ALU_OUT2s_13_port
                           , ALU_OUT2(12) => ALU_OUT2s_12_port, ALU_OUT2(11) =>
                           ALU_OUT2s_11_port, ALU_OUT2(10) => ALU_OUT2s_10_port
                           , ALU_OUT2(9) => ALU_OUT2s_9_port, ALU_OUT2(8) => 
                           ALU_OUT2s_8_port, ALU_OUT2(7) => ALU_OUT2s_7_port, 
                           ALU_OUT2(6) => ALU_OUT2s_6_port, ALU_OUT2(5) => 
                           ALU_OUT2s_5_port, ALU_OUT2(4) => ALU_OUT2s_4_port, 
                           ALU_OUT2(3) => ALU_OUT2s_3_port, ALU_OUT2(2) => 
                           ALU_OUT2s_2_port, ALU_OUT2(1) => ALU_OUT2s_1_port, 
                           ALU_OUT2(0) => ALU_OUT2s_0_port, IR_IN4(31) => 
                           IR_OUT3s_31_port, IR_IN4(30) => IR_OUT3s_30_port, 
                           IR_IN4(29) => IR_OUT3s_29_port, IR_IN4(28) => 
                           IR_OUT3s_28_port, IR_IN4(27) => IR_OUT3s_27_port, 
                           IR_IN4(26) => IR_OUT3s_26_port, IR_IN4(25) => 
                           IR_OUT3s_25_port, IR_IN4(24) => IR_OUT3s_24_port, 
                           IR_IN4(23) => IR_OUT3s_23_port, IR_IN4(22) => 
                           IR_OUT3s_22_port, IR_IN4(21) => IR_OUT3s_21_port, 
                           IR_IN4(20) => IR_OUT3s_20_port, IR_IN4(19) => 
                           IR_OUT3s_19_port, IR_IN4(18) => IR_OUT3s_18_port, 
                           IR_IN4(17) => IR_OUT3s_17_port, IR_IN4(16) => 
                           IR_OUT3s_16_port, IR_IN4(15) => IR_OUT3s_15_port, 
                           IR_IN4(14) => IR_OUT3s_14_port, IR_IN4(13) => 
                           IR_OUT3s_13_port, IR_IN4(12) => IR_OUT3s_12_port, 
                           IR_IN4(11) => IR_OUT3s_11_port, IR_IN4(10) => 
                           IR_OUT3s_10_port, IR_IN4(9) => IR_OUT3s_9_port, 
                           IR_IN4(8) => IR_OUT3s_8_port, IR_IN4(7) => 
                           IR_OUT3s_7_port, IR_IN4(6) => IR_OUT3s_6_port, 
                           IR_IN4(5) => IR_OUT3s_5_port, IR_IN4(4) => 
                           IR_OUT3s_4_port, IR_IN4(3) => IR_OUT3s_3_port, 
                           IR_IN4(2) => IR_OUT3s_2_port, IR_IN4(1) => 
                           IR_OUT3s_1_port, IR_IN4(0) => IR_OUT3s_0_port, 
                           IR_OUT4(31) => IR_OUT4s_31_port, IR_OUT4(30) => 
                           IR_OUT4s_30_port, IR_OUT4(29) => IR_OUT4s_29_port, 
                           IR_OUT4(28) => IR_OUT4s_28_port, IR_OUT4(27) => 
                           IR_OUT4s_27_port, IR_OUT4(26) => IR_OUT4s_26_port, 
                           IR_OUT4(25) => IR_OUT4s_25_port, IR_OUT4(24) => 
                           IR_OUT4s_24_port, IR_OUT4(23) => IR_OUT4s_23_port, 
                           IR_OUT4(22) => IR_OUT4s_22_port, IR_OUT4(21) => 
                           IR_OUT4s_21_port, IR_OUT4(20) => IR_OUT4s_20_port, 
                           IR_OUT4(19) => IR_OUT4s_19_port, IR_OUT4(18) => 
                           IR_OUT4s_18_port, IR_OUT4(17) => IR_OUT4s_17_port, 
                           IR_OUT4(16) => IR_OUT4s_16_port, IR_OUT4(15) => 
                           IR_OUT4s_15_port, IR_OUT4(14) => IR_OUT4s_14_port, 
                           IR_OUT4(13) => IR_OUT4s_13_port, IR_OUT4(12) => 
                           IR_OUT4s_12_port, IR_OUT4(11) => IR_OUT4s_11_port, 
                           IR_OUT4(10) => IR_OUT4s_10_port, IR_OUT4(9) => 
                           IR_OUT4s_9_port, IR_OUT4(8) => IR_OUT4s_8_port, 
                           IR_OUT4(7) => IR_OUT4s_7_port, IR_OUT4(6) => 
                           IR_OUT4s_6_port, IR_OUT4(5) => IR_OUT4s_5_port, 
                           IR_OUT4(4) => IR_OUT4s_4_port, IR_OUT4(3) => 
                           IR_OUT4s_3_port, IR_OUT4(2) => IR_OUT4s_2_port, 
                           IR_OUT4(1) => IR_OUT4s_1_port, IR_OUT4(0) => 
                           IR_OUT4s_0_port);
   WB : writeBack_nbits32 port map( LMD_OUT(31) => LMD_OUTs_31_port, 
                           LMD_OUT(30) => LMD_OUTs_30_port, LMD_OUT(29) => 
                           LMD_OUTs_29_port, LMD_OUT(28) => LMD_OUTs_28_port, 
                           LMD_OUT(27) => LMD_OUTs_27_port, LMD_OUT(26) => 
                           LMD_OUTs_26_port, LMD_OUT(25) => LMD_OUTs_25_port, 
                           LMD_OUT(24) => LMD_OUTs_24_port, LMD_OUT(23) => 
                           LMD_OUTs_23_port, LMD_OUT(22) => LMD_OUTs_22_port, 
                           LMD_OUT(21) => LMD_OUTs_21_port, LMD_OUT(20) => 
                           LMD_OUTs_20_port, LMD_OUT(19) => LMD_OUTs_19_port, 
                           LMD_OUT(18) => LMD_OUTs_18_port, LMD_OUT(17) => 
                           LMD_OUTs_17_port, LMD_OUT(16) => LMD_OUTs_16_port, 
                           LMD_OUT(15) => LMD_OUTs_15_port, LMD_OUT(14) => 
                           LMD_OUTs_14_port, LMD_OUT(13) => LMD_OUTs_13_port, 
                           LMD_OUT(12) => LMD_OUTs_12_port, LMD_OUT(11) => 
                           LMD_OUTs_11_port, LMD_OUT(10) => LMD_OUTs_10_port, 
                           LMD_OUT(9) => LMD_OUTs_9_port, LMD_OUT(8) => 
                           LMD_OUTs_8_port, LMD_OUT(7) => LMD_OUTs_7_port, 
                           LMD_OUT(6) => LMD_OUTs_6_port, LMD_OUT(5) => 
                           LMD_OUTs_5_port, LMD_OUT(4) => LMD_OUTs_4_port, 
                           LMD_OUT(3) => LMD_OUTs_3_port, LMD_OUT(2) => 
                           LMD_OUTs_2_port, LMD_OUT(1) => LMD_OUTs_1_port, 
                           LMD_OUT(0) => LMD_OUTs_0_port, ALUREG_OUTPUT(31) => 
                           ALU_OUT2s_31_port, ALUREG_OUTPUT(30) => 
                           ALU_OUT2s_30_port, ALUREG_OUTPUT(29) => 
                           ALU_OUT2s_29_port, ALUREG_OUTPUT(28) => 
                           ALU_OUT2s_28_port, ALUREG_OUTPUT(27) => 
                           ALU_OUT2s_27_port, ALUREG_OUTPUT(26) => 
                           ALU_OUT2s_26_port, ALUREG_OUTPUT(25) => 
                           ALU_OUT2s_25_port, ALUREG_OUTPUT(24) => 
                           ALU_OUT2s_24_port, ALUREG_OUTPUT(23) => 
                           ALU_OUT2s_23_port, ALUREG_OUTPUT(22) => 
                           ALU_OUT2s_22_port, ALUREG_OUTPUT(21) => 
                           ALU_OUT2s_21_port, ALUREG_OUTPUT(20) => 
                           ALU_OUT2s_20_port, ALUREG_OUTPUT(19) => 
                           ALU_OUT2s_19_port, ALUREG_OUTPUT(18) => 
                           ALU_OUT2s_18_port, ALUREG_OUTPUT(17) => 
                           ALU_OUT2s_17_port, ALUREG_OUTPUT(16) => 
                           ALU_OUT2s_16_port, ALUREG_OUTPUT(15) => 
                           ALU_OUT2s_15_port, ALUREG_OUTPUT(14) => 
                           ALU_OUT2s_14_port, ALUREG_OUTPUT(13) => 
                           ALU_OUT2s_13_port, ALUREG_OUTPUT(12) => 
                           ALU_OUT2s_12_port, ALUREG_OUTPUT(11) => 
                           ALU_OUT2s_11_port, ALUREG_OUTPUT(10) => 
                           ALU_OUT2s_10_port, ALUREG_OUTPUT(9) => 
                           ALU_OUT2s_9_port, ALUREG_OUTPUT(8) => 
                           ALU_OUT2s_8_port, ALUREG_OUTPUT(7) => 
                           ALU_OUT2s_7_port, ALUREG_OUTPUT(6) => 
                           ALU_OUT2s_6_port, ALUREG_OUTPUT(5) => 
                           ALU_OUT2s_5_port, ALUREG_OUTPUT(4) => 
                           ALU_OUT2s_4_port, ALUREG_OUTPUT(3) => 
                           ALU_OUT2s_3_port, ALUREG_OUTPUT(2) => 
                           ALU_OUT2s_2_port, ALUREG_OUTPUT(1) => 
                           ALU_OUT2s_1_port, ALUREG_OUTPUT(0) => 
                           ALU_OUT2s_0_port, WB_MUX_SEL => WB_MUX_SEL, 
                           DATAIN_RF(31) => DATAIN_RFs_31_port, DATAIN_RF(30) 
                           => DATAIN_RFs_30_port, DATAIN_RF(29) => 
                           DATAIN_RFs_29_port, DATAIN_RF(28) => 
                           DATAIN_RFs_28_port, DATAIN_RF(27) => 
                           DATAIN_RFs_27_port, DATAIN_RF(26) => 
                           DATAIN_RFs_26_port, DATAIN_RF(25) => 
                           DATAIN_RFs_25_port, DATAIN_RF(24) => 
                           DATAIN_RFs_24_port, DATAIN_RF(23) => 
                           DATAIN_RFs_23_port, DATAIN_RF(22) => 
                           DATAIN_RFs_22_port, DATAIN_RF(21) => 
                           DATAIN_RFs_21_port, DATAIN_RF(20) => 
                           DATAIN_RFs_20_port, DATAIN_RF(19) => 
                           DATAIN_RFs_19_port, DATAIN_RF(18) => 
                           DATAIN_RFs_18_port, DATAIN_RF(17) => 
                           DATAIN_RFs_17_port, DATAIN_RF(16) => 
                           DATAIN_RFs_16_port, DATAIN_RF(15) => 
                           DATAIN_RFs_15_port, DATAIN_RF(14) => 
                           DATAIN_RFs_14_port, DATAIN_RF(13) => 
                           DATAIN_RFs_13_port, DATAIN_RF(12) => 
                           DATAIN_RFs_12_port, DATAIN_RF(11) => 
                           DATAIN_RFs_11_port, DATAIN_RF(10) => 
                           DATAIN_RFs_10_port, DATAIN_RF(9) => 
                           DATAIN_RFs_9_port, DATAIN_RF(8) => DATAIN_RFs_8_port
                           , DATAIN_RF(7) => DATAIN_RFs_7_port, DATAIN_RF(6) =>
                           DATAIN_RFs_6_port, DATAIN_RF(5) => DATAIN_RFs_5_port
                           , DATAIN_RF(4) => DATAIN_RFs_4_port, DATAIN_RF(3) =>
                           DATAIN_RFs_3_port, DATAIN_RF(2) => DATAIN_RFs_2_port
                           , DATAIN_RF(1) => DATAIN_RFs_1_port, DATAIN_RF(0) =>
                           DATAIN_RFs_0_port);
   U1 : BUF_X1 port map( A => clk, Z => n2);
   U2 : BUF_X1 port map( A => rst, Z => n1);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
         std_logic;  ALU_OPCODE : out std_logic_vector (0 to 3);  DRAM_WE, 
         LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, WB_MUX_SEL, RF_WE : out std_logic
         );

end dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, aluOpcode_i_3_port, aluOpcode_i_2_port, 
      aluOpcode_i_1_port, aluOpcode_i_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n_1405, n_1406, n_1407, n_1408 : std_logic;

begin
   IR_LATCH_EN <= X_Logic1_port;
   NPC_LATCH_EN <= X_Logic1_port;
   PC_LATCH_EN <= X_Logic1_port;
   
   X_Logic1_port <= '1';
   RegIMM_LATCH_EN <= '0';
   RegB_LATCH_EN <= '0';
   RegA_LATCH_EN <= '0';
   aluOpcode1_reg_3_inst : DFFS_X1 port map( D => aluOpcode_i_3_port, CK => Clk
                           , SN => n2, Q => ALU_OPCODE(0), QN => n_1405);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => aluOpcode_i_2_port, CK => Clk
                           , RN => n2, Q => ALU_OPCODE(1), QN => n_1406);
   aluOpcode1_reg_1_inst : DFFS_X1 port map( D => aluOpcode_i_1_port, CK => Clk
                           , SN => n2, Q => ALU_OPCODE(2), QN => n_1407);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => aluOpcode_i_0_port, CK => Clk
                           , RN => n2, Q => ALU_OPCODE(3), QN => n_1408);
   RF_WE <= '0';
   WB_MUX_SEL <= '0';
   JUMP_EN <= '0';
   LMD_LATCH_EN <= '0';
   DRAM_WE <= '0';
   EQ_COND <= '0';
   ALU_OUTREG_EN <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   U3 : XNOR2_X1 port map( A => n16, B => IR_IN(3), ZN => n1);
   U13 : INV_X1 port map( A => Rst, ZN => n2);
   U14 : NAND3_X1 port map( A1 => n3, A2 => n4, A3 => n5, ZN => 
                           aluOpcode_i_3_port);
   U15 : NAND3_X1 port map( A1 => n6, A2 => IR_IN(3), A3 => IR_IN(2), ZN => n3)
                           ;
   U16 : OAI211_X1 port map( C1 => n7, C2 => n8, A => n9, B => n10, ZN => 
                           aluOpcode_i_2_port);
   U17 : NAND3_X1 port map( A1 => n6, A2 => n11, A3 => n12, ZN => n9);
   U18 : MUX2_X1 port map( A => n13, B => n14, S => IR_IN(3), Z => n12);
   U19 : NOR3_X1 port map( A1 => n15, A2 => IR_IN(2), A3 => n16, ZN => n14);
   U20 : AOI21_X1 port map( B1 => n15, B2 => n17, A => n18, ZN => n13);
   U21 : NAND2_X1 port map( A1 => IR_IN(5), A2 => n16, ZN => n17);
   U22 : NAND3_X1 port map( A1 => n19, A2 => n5, A3 => n20, ZN => 
                           aluOpcode_i_1_port);
   U23 : NOR4_X1 port map( A1 => n7, A2 => n21, A3 => n22, A4 => n23, ZN => n20
                           );
   U24 : AOI211_X1 port map( C1 => IR_IN(2), C2 => n24, A => n25, B => n26, ZN 
                           => n23);
   U25 : INV_X1 port map( A => n10, ZN => n22);
   U26 : INV_X1 port map( A => n27, ZN => n5);
   U27 : OAI211_X1 port map( C1 => n28, C2 => n25, A => n29, B => n30, ZN => 
                           n27);
   U28 : MUX2_X1 port map( A => n31, B => n32, S => IR_IN(30), Z => n30);
   U29 : AOI21_X1 port map( B1 => n33, B2 => n34, A => n35, ZN => n32);
   U30 : MUX2_X1 port map( A => IR_IN(26), B => IR_IN(27), S => IR_IN(29), Z =>
                           n35);
   U31 : NAND3_X1 port map( A1 => n36, A2 => n34, A3 => IR_IN(26), ZN => n31);
   U32 : MUX2_X1 port map( A => n37, B => n38, S => n7, Z => n29);
   U33 : NOR2_X1 port map( A1 => n36, A2 => n33, ZN => n7);
   U34 : NOR2_X1 port map( A1 => IR_IN(28), A2 => n39, ZN => n38);
   U35 : AOI21_X1 port map( B1 => IR_IN(27), B2 => n40, A => IR_IN(31), ZN => 
                           n37);
   U36 : AND3_X1 port map( A1 => n11, A2 => n41, A3 => n42, ZN => n28);
   U37 : OAI21_X1 port map( B1 => n1, B2 => n26, A => n18, ZN => n42);
   U38 : INV_X1 port map( A => IR_IN(5), ZN => n26);
   U39 : INV_X1 port map( A => IR_IN(0), ZN => n16);
   U40 : OAI21_X1 port map( B1 => IR_IN(3), B2 => IR_IN(0), A => n15, ZN => n41
                           );
   U41 : AOI22_X1 port map( A1 => n40, A2 => IR_IN(28), B1 => n43, B2 => 
                           IR_IN(27), ZN => n19);
   U42 : NAND3_X1 port map( A1 => n44, A2 => n10, A3 => n45, ZN => 
                           aluOpcode_i_0_port);
   U43 : MUX2_X1 port map( A => n46, B => n47, S => IR_IN(26), Z => n45);
   U44 : OAI21_X1 port map( B1 => n48, B2 => n43, A => n36, ZN => n47);
   U45 : INV_X1 port map( A => n8, ZN => n43);
   U46 : NAND4_X1 port map( A1 => IR_IN(29), A2 => IR_IN(28), A3 => n49, A4 => 
                           n39, ZN => n8);
   U47 : INV_X1 port map( A => n4, ZN => n48);
   U48 : NAND4_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), A3 => IR_IN(28), 
                           A4 => n39, ZN => n4);
   U49 : OAI211_X1 port map( C1 => n50, C2 => n21, A => n39, B => IR_IN(27), ZN
                           => n46);
   U50 : INV_X1 port map( A => IR_IN(31), ZN => n39);
   U51 : AND3_X1 port map( A1 => n34, A2 => n49, A3 => IR_IN(29), ZN => n21);
   U52 : NOR3_X1 port map( A1 => n49, A2 => IR_IN(29), A3 => n34, ZN => n50);
   U53 : INV_X1 port map( A => IR_IN(28), ZN => n34);
   U54 : INV_X1 port map( A => IR_IN(30), ZN => n49);
   U55 : NAND4_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), A3 => IR_IN(26), 
                           A4 => n51, ZN => n10);
   U56 : NOR3_X1 port map( A1 => IR_IN(27), A2 => IR_IN(31), A3 => IR_IN(28), 
                           ZN => n51);
   U57 : NAND3_X1 port map( A1 => n6, A2 => n11, A3 => n52, ZN => n44);
   U58 : MUX2_X1 port map( A => n53, B => n54, S => IR_IN(0), Z => n52);
   U59 : AOI21_X1 port map( B1 => n55, B2 => n18, A => n15, ZN => n54);
   U60 : NAND2_X1 port map( A1 => IR_IN(5), A2 => n24, ZN => n15);
   U61 : INV_X1 port map( A => IR_IN(3), ZN => n55);
   U62 : NOR3_X1 port map( A1 => n24, A2 => IR_IN(3), A3 => n56, ZN => n53);
   U63 : XOR2_X1 port map( A => IR_IN(5), B => n18, Z => n56);
   U64 : INV_X1 port map( A => IR_IN(2), ZN => n18);
   U65 : INV_X1 port map( A => IR_IN(1), ZN => n24);
   U66 : NOR4_X1 port map( A1 => IR_IN(6), A2 => IR_IN(4), A3 => IR_IN(10), A4 
                           => n57, ZN => n11);
   U67 : OR3_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), ZN =>
                           n57);
   U68 : INV_X1 port map( A => n25, ZN => n6);
   U69 : NAND4_X1 port map( A1 => n40, A2 => n33, A3 => n58, A4 => n36, ZN => 
                           n25);
   U70 : INV_X1 port map( A => IR_IN(27), ZN => n36);
   U71 : NOR2_X1 port map( A1 => IR_IN(31), A2 => IR_IN(28), ZN => n58);
   U72 : INV_X1 port map( A => IR_IN(26), ZN => n33);
   U73 : NOR2_X1 port map( A1 => IR_IN(29), A2 => IR_IN(30), ZN => n40);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity dlx is

   port( Clk_port, Rst_port : in std_logic;  DATA_IRAM_port, DATAread_DRAM_port
         : in std_logic_vector (31 downto 0);  WE_DRAM_port : out std_logic;  
         ADDRESS_DRAM_port, DATAwrite_DRAM_port, ADDRESS_IRAM_port : out 
         std_logic_vector (31 downto 0));

end dlx;

architecture SYN_STRUCTURAL of dlx is

   component datapath_nbits32
      port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 
            downto 0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN, RegA_LATCH_EN, 
            RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE, MUXA_SEL, MUXB_SEL, 
            ALU_OUTREG_EN, EQ_COND : in std_logic;  ALU_OPCODE : in 
            std_logic_vector (0 to 3);  DRAM_DATA : in std_logic_vector (31 
            downto 0);  LMD_LATCH_EN, JUMP_EN, WB_MUX_SEL : in std_logic;  B, 
            ALU_OUT, ADDRESS_IRAM, IR_OUT : out std_logic_vector (31 downto 0)
            );
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
            std_logic;  ALU_OPCODE : out std_logic_vector (0 to 3);  DRAM_WE, 
            LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, WB_MUX_SEL, RF_WE : out 
            std_logic);
   end component;
   
   signal IR_OUT_signal_31_port, IR_OUT_signal_30_port, IR_OUT_signal_29_port, 
      IR_OUT_signal_28_port, IR_OUT_signal_27_port, IR_OUT_signal_26_port, 
      IR_OUT_signal_25_port, IR_OUT_signal_24_port, IR_OUT_signal_23_port, 
      IR_OUT_signal_22_port, IR_OUT_signal_21_port, IR_OUT_signal_20_port, 
      IR_OUT_signal_19_port, IR_OUT_signal_18_port, IR_OUT_signal_17_port, 
      IR_OUT_signal_16_port, IR_OUT_signal_15_port, IR_OUT_signal_14_port, 
      IR_OUT_signal_13_port, IR_OUT_signal_12_port, IR_OUT_signal_11_port, 
      IR_OUT_signal_10_port, IR_OUT_signal_9_port, IR_OUT_signal_8_port, 
      IR_OUT_signal_7_port, IR_OUT_signal_6_port, IR_OUT_signal_5_port, 
      IR_OUT_signal_4_port, IR_OUT_signal_3_port, IR_OUT_signal_2_port, 
      IR_OUT_signal_1_port, IR_OUT_signal_0_port, IR_LATCH_EN_signal, 
      NPC_LATCH_EN_signal, RegA_LATCH_EN_signal, RegB_LATCH_EN_signal, 
      RegIMM_LATCH_EN_signal, MUXA_SEL_signal, MUXB_SEL_signal, 
      ALU_OUTREG_EN_signal, EQ_COND_signal, ALU_OPCODE_signal_0_port, 
      ALU_OPCODE_signal_1_port, ALU_OPCODE_signal_2_port, 
      ALU_OPCODE_signal_3_port, LMD_LATCH_EN_signal, JUMP_EN_signal, 
      PC_LATCH_EN_signal, WB_MUX_SEL_signal, RF_WE_signal, n_1409, n_1410, 
      n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, 
      n_1420, n_1421, n_1422, n_1423 : std_logic;

begin
   
   CONTROL_UNIT : 
                           dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 
                           port map( Clk => Clk_port, Rst => Rst_port, 
                           IR_IN(31) => IR_OUT_signal_31_port, IR_IN(30) => 
                           IR_OUT_signal_30_port, IR_IN(29) => 
                           IR_OUT_signal_29_port, IR_IN(28) => 
                           IR_OUT_signal_28_port, IR_IN(27) => 
                           IR_OUT_signal_27_port, IR_IN(26) => 
                           IR_OUT_signal_26_port, IR_IN(25) => 
                           IR_OUT_signal_25_port, IR_IN(24) => 
                           IR_OUT_signal_24_port, IR_IN(23) => 
                           IR_OUT_signal_23_port, IR_IN(22) => 
                           IR_OUT_signal_22_port, IR_IN(21) => 
                           IR_OUT_signal_21_port, IR_IN(20) => 
                           IR_OUT_signal_20_port, IR_IN(19) => 
                           IR_OUT_signal_19_port, IR_IN(18) => 
                           IR_OUT_signal_18_port, IR_IN(17) => 
                           IR_OUT_signal_17_port, IR_IN(16) => 
                           IR_OUT_signal_16_port, IR_IN(15) => 
                           IR_OUT_signal_15_port, IR_IN(14) => 
                           IR_OUT_signal_14_port, IR_IN(13) => 
                           IR_OUT_signal_13_port, IR_IN(12) => 
                           IR_OUT_signal_12_port, IR_IN(11) => 
                           IR_OUT_signal_11_port, IR_IN(10) => 
                           IR_OUT_signal_10_port, IR_IN(9) => 
                           IR_OUT_signal_9_port, IR_IN(8) => 
                           IR_OUT_signal_8_port, IR_IN(7) => 
                           IR_OUT_signal_7_port, IR_IN(6) => 
                           IR_OUT_signal_6_port, IR_IN(5) => 
                           IR_OUT_signal_5_port, IR_IN(4) => 
                           IR_OUT_signal_4_port, IR_IN(3) => 
                           IR_OUT_signal_3_port, IR_IN(2) => 
                           IR_OUT_signal_2_port, IR_IN(1) => 
                           IR_OUT_signal_1_port, IR_IN(0) => 
                           IR_OUT_signal_0_port, IR_LATCH_EN => n_1409, 
                           NPC_LATCH_EN => n_1410, RegA_LATCH_EN => n_1411, 
                           RegB_LATCH_EN => n_1412, RegIMM_LATCH_EN => n_1413, 
                           MUXA_SEL => n_1414, MUXB_SEL => n_1415, 
                           ALU_OUTREG_EN => n_1416, EQ_COND => n_1417, 
                           ALU_OPCODE(0) => ALU_OPCODE_signal_0_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_signal_1_port, 
                           ALU_OPCODE(2) => ALU_OPCODE_signal_2_port, 
                           ALU_OPCODE(3) => ALU_OPCODE_signal_3_port, DRAM_WE 
                           => n_1418, LMD_LATCH_EN => n_1419, JUMP_EN => n_1420
                           , PC_LATCH_EN => n_1421, WB_MUX_SEL => n_1422, RF_WE
                           => n_1423);
   DATA_PATH : datapath_nbits32 port map( clk => Clk_port, rst => Rst_port, 
                           DATA_IRAM(31) => DATA_IRAM_port(31), DATA_IRAM(30) 
                           => DATA_IRAM_port(30), DATA_IRAM(29) => 
                           DATA_IRAM_port(29), DATA_IRAM(28) => 
                           DATA_IRAM_port(28), DATA_IRAM(27) => 
                           DATA_IRAM_port(27), DATA_IRAM(26) => 
                           DATA_IRAM_port(26), DATA_IRAM(25) => 
                           DATA_IRAM_port(25), DATA_IRAM(24) => 
                           DATA_IRAM_port(24), DATA_IRAM(23) => 
                           DATA_IRAM_port(23), DATA_IRAM(22) => 
                           DATA_IRAM_port(22), DATA_IRAM(21) => 
                           DATA_IRAM_port(21), DATA_IRAM(20) => 
                           DATA_IRAM_port(20), DATA_IRAM(19) => 
                           DATA_IRAM_port(19), DATA_IRAM(18) => 
                           DATA_IRAM_port(18), DATA_IRAM(17) => 
                           DATA_IRAM_port(17), DATA_IRAM(16) => 
                           DATA_IRAM_port(16), DATA_IRAM(15) => 
                           DATA_IRAM_port(15), DATA_IRAM(14) => 
                           DATA_IRAM_port(14), DATA_IRAM(13) => 
                           DATA_IRAM_port(13), DATA_IRAM(12) => 
                           DATA_IRAM_port(12), DATA_IRAM(11) => 
                           DATA_IRAM_port(11), DATA_IRAM(10) => 
                           DATA_IRAM_port(10), DATA_IRAM(9) => 
                           DATA_IRAM_port(9), DATA_IRAM(8) => DATA_IRAM_port(8)
                           , DATA_IRAM(7) => DATA_IRAM_port(7), DATA_IRAM(6) =>
                           DATA_IRAM_port(6), DATA_IRAM(5) => DATA_IRAM_port(5)
                           , DATA_IRAM(4) => DATA_IRAM_port(4), DATA_IRAM(3) =>
                           DATA_IRAM_port(3), DATA_IRAM(2) => DATA_IRAM_port(2)
                           , DATA_IRAM(1) => DATA_IRAM_port(1), DATA_IRAM(0) =>
                           DATA_IRAM_port(0), IR_LATCH_EN => IR_LATCH_EN_signal
                           , NPC_LATCH_EN => NPC_LATCH_EN_signal, PC_LATCH_EN 
                           => PC_LATCH_EN_signal, RegA_LATCH_EN => 
                           RegA_LATCH_EN_signal, RegB_LATCH_EN => 
                           RegB_LATCH_EN_signal, RegIMM_LATCH_EN => 
                           RegIMM_LATCH_EN_signal, RF_WE => RF_WE_signal, 
                           MUXA_SEL => MUXA_SEL_signal, MUXB_SEL => 
                           MUXB_SEL_signal, ALU_OUTREG_EN => 
                           ALU_OUTREG_EN_signal, EQ_COND => EQ_COND_signal, 
                           ALU_OPCODE(0) => ALU_OPCODE_signal_0_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_signal_1_port, 
                           ALU_OPCODE(2) => ALU_OPCODE_signal_2_port, 
                           ALU_OPCODE(3) => ALU_OPCODE_signal_3_port, 
                           DRAM_DATA(31) => DATAread_DRAM_port(31), 
                           DRAM_DATA(30) => DATAread_DRAM_port(30), 
                           DRAM_DATA(29) => DATAread_DRAM_port(29), 
                           DRAM_DATA(28) => DATAread_DRAM_port(28), 
                           DRAM_DATA(27) => DATAread_DRAM_port(27), 
                           DRAM_DATA(26) => DATAread_DRAM_port(26), 
                           DRAM_DATA(25) => DATAread_DRAM_port(25), 
                           DRAM_DATA(24) => DATAread_DRAM_port(24), 
                           DRAM_DATA(23) => DATAread_DRAM_port(23), 
                           DRAM_DATA(22) => DATAread_DRAM_port(22), 
                           DRAM_DATA(21) => DATAread_DRAM_port(21), 
                           DRAM_DATA(20) => DATAread_DRAM_port(20), 
                           DRAM_DATA(19) => DATAread_DRAM_port(19), 
                           DRAM_DATA(18) => DATAread_DRAM_port(18), 
                           DRAM_DATA(17) => DATAread_DRAM_port(17), 
                           DRAM_DATA(16) => DATAread_DRAM_port(16), 
                           DRAM_DATA(15) => DATAread_DRAM_port(15), 
                           DRAM_DATA(14) => DATAread_DRAM_port(14), 
                           DRAM_DATA(13) => DATAread_DRAM_port(13), 
                           DRAM_DATA(12) => DATAread_DRAM_port(12), 
                           DRAM_DATA(11) => DATAread_DRAM_port(11), 
                           DRAM_DATA(10) => DATAread_DRAM_port(10), 
                           DRAM_DATA(9) => DATAread_DRAM_port(9), DRAM_DATA(8) 
                           => DATAread_DRAM_port(8), DRAM_DATA(7) => 
                           DATAread_DRAM_port(7), DRAM_DATA(6) => 
                           DATAread_DRAM_port(6), DRAM_DATA(5) => 
                           DATAread_DRAM_port(5), DRAM_DATA(4) => 
                           DATAread_DRAM_port(4), DRAM_DATA(3) => 
                           DATAread_DRAM_port(3), DRAM_DATA(2) => 
                           DATAread_DRAM_port(2), DRAM_DATA(1) => 
                           DATAread_DRAM_port(1), DRAM_DATA(0) => 
                           DATAread_DRAM_port(0), LMD_LATCH_EN => 
                           LMD_LATCH_EN_signal, JUMP_EN => JUMP_EN_signal, 
                           WB_MUX_SEL => WB_MUX_SEL_signal, B(31) => 
                           DATAwrite_DRAM_port(31), B(30) => 
                           DATAwrite_DRAM_port(30), B(29) => 
                           DATAwrite_DRAM_port(29), B(28) => 
                           DATAwrite_DRAM_port(28), B(27) => 
                           DATAwrite_DRAM_port(27), B(26) => 
                           DATAwrite_DRAM_port(26), B(25) => 
                           DATAwrite_DRAM_port(25), B(24) => 
                           DATAwrite_DRAM_port(24), B(23) => 
                           DATAwrite_DRAM_port(23), B(22) => 
                           DATAwrite_DRAM_port(22), B(21) => 
                           DATAwrite_DRAM_port(21), B(20) => 
                           DATAwrite_DRAM_port(20), B(19) => 
                           DATAwrite_DRAM_port(19), B(18) => 
                           DATAwrite_DRAM_port(18), B(17) => 
                           DATAwrite_DRAM_port(17), B(16) => 
                           DATAwrite_DRAM_port(16), B(15) => 
                           DATAwrite_DRAM_port(15), B(14) => 
                           DATAwrite_DRAM_port(14), B(13) => 
                           DATAwrite_DRAM_port(13), B(12) => 
                           DATAwrite_DRAM_port(12), B(11) => 
                           DATAwrite_DRAM_port(11), B(10) => 
                           DATAwrite_DRAM_port(10), B(9) => 
                           DATAwrite_DRAM_port(9), B(8) => 
                           DATAwrite_DRAM_port(8), B(7) => 
                           DATAwrite_DRAM_port(7), B(6) => 
                           DATAwrite_DRAM_port(6), B(5) => 
                           DATAwrite_DRAM_port(5), B(4) => 
                           DATAwrite_DRAM_port(4), B(3) => 
                           DATAwrite_DRAM_port(3), B(2) => 
                           DATAwrite_DRAM_port(2), B(1) => 
                           DATAwrite_DRAM_port(1), B(0) => 
                           DATAwrite_DRAM_port(0), ALU_OUT(31) => 
                           ADDRESS_DRAM_port(31), ALU_OUT(30) => 
                           ADDRESS_DRAM_port(30), ALU_OUT(29) => 
                           ADDRESS_DRAM_port(29), ALU_OUT(28) => 
                           ADDRESS_DRAM_port(28), ALU_OUT(27) => 
                           ADDRESS_DRAM_port(27), ALU_OUT(26) => 
                           ADDRESS_DRAM_port(26), ALU_OUT(25) => 
                           ADDRESS_DRAM_port(25), ALU_OUT(24) => 
                           ADDRESS_DRAM_port(24), ALU_OUT(23) => 
                           ADDRESS_DRAM_port(23), ALU_OUT(22) => 
                           ADDRESS_DRAM_port(22), ALU_OUT(21) => 
                           ADDRESS_DRAM_port(21), ALU_OUT(20) => 
                           ADDRESS_DRAM_port(20), ALU_OUT(19) => 
                           ADDRESS_DRAM_port(19), ALU_OUT(18) => 
                           ADDRESS_DRAM_port(18), ALU_OUT(17) => 
                           ADDRESS_DRAM_port(17), ALU_OUT(16) => 
                           ADDRESS_DRAM_port(16), ALU_OUT(15) => 
                           ADDRESS_DRAM_port(15), ALU_OUT(14) => 
                           ADDRESS_DRAM_port(14), ALU_OUT(13) => 
                           ADDRESS_DRAM_port(13), ALU_OUT(12) => 
                           ADDRESS_DRAM_port(12), ALU_OUT(11) => 
                           ADDRESS_DRAM_port(11), ALU_OUT(10) => 
                           ADDRESS_DRAM_port(10), ALU_OUT(9) => 
                           ADDRESS_DRAM_port(9), ALU_OUT(8) => 
                           ADDRESS_DRAM_port(8), ALU_OUT(7) => 
                           ADDRESS_DRAM_port(7), ALU_OUT(6) => 
                           ADDRESS_DRAM_port(6), ALU_OUT(5) => 
                           ADDRESS_DRAM_port(5), ALU_OUT(4) => 
                           ADDRESS_DRAM_port(4), ALU_OUT(3) => 
                           ADDRESS_DRAM_port(3), ALU_OUT(2) => 
                           ADDRESS_DRAM_port(2), ALU_OUT(1) => 
                           ADDRESS_DRAM_port(1), ALU_OUT(0) => 
                           ADDRESS_DRAM_port(0), ADDRESS_IRAM(31) => 
                           ADDRESS_IRAM_port(31), ADDRESS_IRAM(30) => 
                           ADDRESS_IRAM_port(30), ADDRESS_IRAM(29) => 
                           ADDRESS_IRAM_port(29), ADDRESS_IRAM(28) => 
                           ADDRESS_IRAM_port(28), ADDRESS_IRAM(27) => 
                           ADDRESS_IRAM_port(27), ADDRESS_IRAM(26) => 
                           ADDRESS_IRAM_port(26), ADDRESS_IRAM(25) => 
                           ADDRESS_IRAM_port(25), ADDRESS_IRAM(24) => 
                           ADDRESS_IRAM_port(24), ADDRESS_IRAM(23) => 
                           ADDRESS_IRAM_port(23), ADDRESS_IRAM(22) => 
                           ADDRESS_IRAM_port(22), ADDRESS_IRAM(21) => 
                           ADDRESS_IRAM_port(21), ADDRESS_IRAM(20) => 
                           ADDRESS_IRAM_port(20), ADDRESS_IRAM(19) => 
                           ADDRESS_IRAM_port(19), ADDRESS_IRAM(18) => 
                           ADDRESS_IRAM_port(18), ADDRESS_IRAM(17) => 
                           ADDRESS_IRAM_port(17), ADDRESS_IRAM(16) => 
                           ADDRESS_IRAM_port(16), ADDRESS_IRAM(15) => 
                           ADDRESS_IRAM_port(15), ADDRESS_IRAM(14) => 
                           ADDRESS_IRAM_port(14), ADDRESS_IRAM(13) => 
                           ADDRESS_IRAM_port(13), ADDRESS_IRAM(12) => 
                           ADDRESS_IRAM_port(12), ADDRESS_IRAM(11) => 
                           ADDRESS_IRAM_port(11), ADDRESS_IRAM(10) => 
                           ADDRESS_IRAM_port(10), ADDRESS_IRAM(9) => 
                           ADDRESS_IRAM_port(9), ADDRESS_IRAM(8) => 
                           ADDRESS_IRAM_port(8), ADDRESS_IRAM(7) => 
                           ADDRESS_IRAM_port(7), ADDRESS_IRAM(6) => 
                           ADDRESS_IRAM_port(6), ADDRESS_IRAM(5) => 
                           ADDRESS_IRAM_port(5), ADDRESS_IRAM(4) => 
                           ADDRESS_IRAM_port(4), ADDRESS_IRAM(3) => 
                           ADDRESS_IRAM_port(3), ADDRESS_IRAM(2) => 
                           ADDRESS_IRAM_port(2), ADDRESS_IRAM(1) => 
                           ADDRESS_IRAM_port(1), ADDRESS_IRAM(0) => 
                           ADDRESS_IRAM_port(0), IR_OUT(31) => 
                           IR_OUT_signal_31_port, IR_OUT(30) => 
                           IR_OUT_signal_30_port, IR_OUT(29) => 
                           IR_OUT_signal_29_port, IR_OUT(28) => 
                           IR_OUT_signal_28_port, IR_OUT(27) => 
                           IR_OUT_signal_27_port, IR_OUT(26) => 
                           IR_OUT_signal_26_port, IR_OUT(25) => 
                           IR_OUT_signal_25_port, IR_OUT(24) => 
                           IR_OUT_signal_24_port, IR_OUT(23) => 
                           IR_OUT_signal_23_port, IR_OUT(22) => 
                           IR_OUT_signal_22_port, IR_OUT(21) => 
                           IR_OUT_signal_21_port, IR_OUT(20) => 
                           IR_OUT_signal_20_port, IR_OUT(19) => 
                           IR_OUT_signal_19_port, IR_OUT(18) => 
                           IR_OUT_signal_18_port, IR_OUT(17) => 
                           IR_OUT_signal_17_port, IR_OUT(16) => 
                           IR_OUT_signal_16_port, IR_OUT(15) => 
                           IR_OUT_signal_15_port, IR_OUT(14) => 
                           IR_OUT_signal_14_port, IR_OUT(13) => 
                           IR_OUT_signal_13_port, IR_OUT(12) => 
                           IR_OUT_signal_12_port, IR_OUT(11) => 
                           IR_OUT_signal_11_port, IR_OUT(10) => 
                           IR_OUT_signal_10_port, IR_OUT(9) => 
                           IR_OUT_signal_9_port, IR_OUT(8) => 
                           IR_OUT_signal_8_port, IR_OUT(7) => 
                           IR_OUT_signal_7_port, IR_OUT(6) => 
                           IR_OUT_signal_6_port, IR_OUT(5) => 
                           IR_OUT_signal_5_port, IR_OUT(4) => 
                           IR_OUT_signal_4_port, IR_OUT(3) => 
                           IR_OUT_signal_3_port, IR_OUT(2) => 
                           IR_OUT_signal_2_port, IR_OUT(1) => 
                           IR_OUT_signal_1_port, IR_OUT(0) => 
                           IR_OUT_signal_0_port);
   RF_WE_signal <= '0';
   WB_MUX_SEL_signal <= '0';
   PC_LATCH_EN_signal <= '1';
   JUMP_EN_signal <= '0';
   LMD_LATCH_EN_signal <= '0';
   WE_DRAM_port <= '0';
   EQ_COND_signal <= '0';
   ALU_OUTREG_EN_signal <= '0';
   MUXB_SEL_signal <= '0';
   MUXA_SEL_signal <= '0';
   RegIMM_LATCH_EN_signal <= '0';
   RegB_LATCH_EN_signal <= '0';
   RegA_LATCH_EN_signal <= '0';
   NPC_LATCH_EN_signal <= '1';
   IR_LATCH_EN_signal <= '1';

end SYN_STRUCTURAL;
