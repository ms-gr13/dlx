
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_top is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_top;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top.all;

entity top is

   port( Clk_port_top, Rst_port_top : in std_logic);

end top;

architecture SYN_STRUCTURAL of top is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component alu
      port( FUNC : in std_logic_vector (3 downto 0);  A, B : in 
            std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
            downto 0));
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component dram
      port( clk, w_r : in std_logic;  addr, data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component IRAM
      port( Rst : in std_logic;  Addr : in std_logic_vector (31 downto 0);  
            Dout : out std_logic_vector (31 downto 0));
   end component;
   
   signal DATA_IRAM_signal_31_port, DATA_IRAM_signal_30_port, 
      DATA_IRAM_signal_29_port, DATA_IRAM_signal_28_port, 
      DATA_IRAM_signal_27_port, DATA_IRAM_signal_26_port, 
      DATA_IRAM_signal_25_port, DATA_IRAM_signal_24_port, 
      DATA_IRAM_signal_23_port, DATA_IRAM_signal_22_port, 
      DATA_IRAM_signal_21_port, DATA_IRAM_signal_20_port, 
      DATA_IRAM_signal_19_port, DATA_IRAM_signal_18_port, 
      DATA_IRAM_signal_17_port, DATA_IRAM_signal_16_port, 
      DATA_IRAM_signal_15_port, DATA_IRAM_signal_14_port, 
      DATA_IRAM_signal_13_port, DATA_IRAM_signal_12_port, 
      DATA_IRAM_signal_11_port, DATA_IRAM_signal_10_port, 
      DATA_IRAM_signal_9_port, DATA_IRAM_signal_8_port, DATA_IRAM_signal_7_port
      , DATA_IRAM_signal_6_port, DATA_IRAM_signal_5_port, 
      DATA_IRAM_signal_4_port, DATA_IRAM_signal_3_port, DATA_IRAM_signal_2_port
      , DATA_IRAM_signal_1_port, DATA_IRAM_signal_0_port, 
      ADDRESS_DRAM_signal_31_port, ADDRESS_DRAM_signal_30_port, 
      ADDRESS_DRAM_signal_29_port, ADDRESS_DRAM_signal_28_port, 
      ADDRESS_DRAM_signal_27_port, ADDRESS_DRAM_signal_26_port, 
      ADDRESS_DRAM_signal_25_port, ADDRESS_DRAM_signal_24_port, 
      ADDRESS_DRAM_signal_23_port, ADDRESS_DRAM_signal_22_port, 
      ADDRESS_DRAM_signal_21_port, ADDRESS_DRAM_signal_20_port, 
      ADDRESS_DRAM_signal_19_port, ADDRESS_DRAM_signal_18_port, 
      ADDRESS_DRAM_signal_17_port, ADDRESS_DRAM_signal_16_port, 
      ADDRESS_DRAM_signal_15_port, ADDRESS_DRAM_signal_14_port, 
      ADDRESS_DRAM_signal_13_port, ADDRESS_DRAM_signal_12_port, 
      ADDRESS_DRAM_signal_11_port, ADDRESS_DRAM_signal_10_port, 
      ADDRESS_DRAM_signal_9_port, ADDRESS_DRAM_signal_8_port, 
      ADDRESS_DRAM_signal_7_port, ADDRESS_DRAM_signal_6_port, 
      ADDRESS_DRAM_signal_5_port, ADDRESS_DRAM_signal_4_port, 
      ADDRESS_DRAM_signal_3_port, ADDRESS_DRAM_signal_2_port, 
      ADDRESS_DRAM_signal_1_port, ADDRESS_DRAM_signal_0_port, 
      DATAwrite_DRAM_signal_31_port, DATAwrite_DRAM_signal_30_port, 
      DATAwrite_DRAM_signal_29_port, DATAwrite_DRAM_signal_28_port, 
      DATAwrite_DRAM_signal_27_port, DATAwrite_DRAM_signal_26_port, 
      DATAwrite_DRAM_signal_25_port, DATAwrite_DRAM_signal_24_port, 
      DATAwrite_DRAM_signal_23_port, DATAwrite_DRAM_signal_22_port, 
      DATAwrite_DRAM_signal_21_port, DATAwrite_DRAM_signal_20_port, 
      DATAwrite_DRAM_signal_19_port, DATAwrite_DRAM_signal_18_port, 
      DATAwrite_DRAM_signal_17_port, DATAwrite_DRAM_signal_16_port, 
      DATAwrite_DRAM_signal_15_port, DATAwrite_DRAM_signal_14_port, 
      DATAwrite_DRAM_signal_13_port, DATAwrite_DRAM_signal_12_port, 
      DATAwrite_DRAM_signal_11_port, DATAwrite_DRAM_signal_10_port, 
      DATAwrite_DRAM_signal_9_port, DATAwrite_DRAM_signal_8_port, 
      DATAwrite_DRAM_signal_7_port, DATAwrite_DRAM_signal_6_port, 
      DATAwrite_DRAM_signal_5_port, DATAwrite_DRAM_signal_4_port, 
      DATAwrite_DRAM_signal_3_port, DATAwrite_DRAM_signal_2_port, 
      DATAwrite_DRAM_signal_1_port, DATAwrite_DRAM_signal_0_port, 
      ADDRESS_IRAM_signal_31_port, ADDRESS_IRAM_signal_30_port, 
      ADDRESS_IRAM_signal_29_port, ADDRESS_IRAM_signal_28_port, 
      ADDRESS_IRAM_signal_27_port, ADDRESS_IRAM_signal_26_port, 
      ADDRESS_IRAM_signal_25_port, ADDRESS_IRAM_signal_24_port, 
      ADDRESS_IRAM_signal_23_port, ADDRESS_IRAM_signal_22_port, 
      ADDRESS_IRAM_signal_21_port, ADDRESS_IRAM_signal_20_port, 
      ADDRESS_IRAM_signal_19_port, ADDRESS_IRAM_signal_18_port, 
      ADDRESS_IRAM_signal_17_port, ADDRESS_IRAM_signal_16_port, 
      ADDRESS_IRAM_signal_15_port, ADDRESS_IRAM_signal_14_port, 
      ADDRESS_IRAM_signal_13_port, ADDRESS_IRAM_signal_12_port, 
      ADDRESS_IRAM_signal_11_port, ADDRESS_IRAM_signal_10_port, 
      ADDRESS_IRAM_signal_9_port, ADDRESS_IRAM_signal_8_port, 
      ADDRESS_IRAM_signal_7_port, ADDRESS_IRAM_signal_6_port, 
      ADDRESS_IRAM_signal_5_port, ADDRESS_IRAM_signal_4_port, 
      ADDRESS_IRAM_signal_3_port, ADDRESS_IRAM_signal_2_port, 
      ADDRESS_IRAM_signal_1_port, ADDRESS_IRAM_signal_0_port, n1, DLX_INST_n2, 
      DLX_INST_RF_WE_signal, DLX_INST_WB_MUX_SEL_signal, 
      DLX_INST_PC_LATCH_EN_signal, DLX_INST_JUMP_EN_signal, 
      DLX_INST_LMD_LATCH_EN_signal, DLX_INST_ALU_OPCODE_signal_3_port, 
      DLX_INST_ALU_OPCODE_signal_2_port, DLX_INST_ALU_OPCODE_signal_1_port, 
      DLX_INST_ALU_OPCODE_signal_0_port, DLX_INST_EQ_COND_signal, 
      DLX_INST_ALU_OUTREG_EN_signal, DLX_INST_MUXB_SEL_signal, 
      DLX_INST_MUXA_SEL_signal, DLX_INST_RegIMM_LATCH_EN_signal, 
      DLX_INST_RegB_LATCH_EN_signal, DLX_INST_RegA_LATCH_EN_signal, 
      DLX_INST_NPC_LATCH_EN_signal, DLX_INST_IR_LATCH_EN_signal, 
      DLX_INST_IR_OUT_signal_16_port, DLX_INST_IR_OUT_signal_17_port, 
      DLX_INST_IR_OUT_signal_18_port, DLX_INST_IR_OUT_signal_19_port, 
      DLX_INST_IR_OUT_signal_20_port, DLX_INST_IR_OUT_signal_21_port, 
      DLX_INST_IR_OUT_signal_22_port, DLX_INST_IR_OUT_signal_23_port, 
      DLX_INST_IR_OUT_signal_24_port, DLX_INST_IR_OUT_signal_25_port, 
      DLX_INST_IR_OUT_signal_26_port, DLX_INST_IR_OUT_signal_27_port, 
      DLX_INST_IR_OUT_signal_28_port, DLX_INST_IR_OUT_signal_29_port, 
      DLX_INST_IR_OUT_signal_30_port, DLX_INST_IR_OUT_signal_31_port, 
      DLX_INST_WE_DRAM_port, DLX_INST_CONTROL_UNIT_n117, 
      DLX_INST_CONTROL_UNIT_n116, DLX_INST_CONTROL_UNIT_n115, 
      DLX_INST_CONTROL_UNIT_n114, DLX_INST_CONTROL_UNIT_n113, 
      DLX_INST_CONTROL_UNIT_n112, DLX_INST_CONTROL_UNIT_n111, 
      DLX_INST_CONTROL_UNIT_n110, DLX_INST_CONTROL_UNIT_n109, 
      DLX_INST_CONTROL_UNIT_n108, DLX_INST_CONTROL_UNIT_n107, 
      DLX_INST_CONTROL_UNIT_n106, DLX_INST_CONTROL_UNIT_n105, 
      DLX_INST_CONTROL_UNIT_n104, DLX_INST_CONTROL_UNIT_n103, 
      DLX_INST_CONTROL_UNIT_n102, DLX_INST_CONTROL_UNIT_n101, 
      DLX_INST_CONTROL_UNIT_n100, DLX_INST_CONTROL_UNIT_n99, 
      DLX_INST_CONTROL_UNIT_n98, DLX_INST_CONTROL_UNIT_n97, 
      DLX_INST_CONTROL_UNIT_n96, DLX_INST_CONTROL_UNIT_n95, 
      DLX_INST_CONTROL_UNIT_n94, DLX_INST_CONTROL_UNIT_n93, 
      DLX_INST_CONTROL_UNIT_n92, DLX_INST_CONTROL_UNIT_n91, 
      DLX_INST_CONTROL_UNIT_n90, DLX_INST_CONTROL_UNIT_n89, 
      DLX_INST_CONTROL_UNIT_n88, DLX_INST_CONTROL_UNIT_n87, 
      DLX_INST_CONTROL_UNIT_n86, DLX_INST_CONTROL_UNIT_n85, 
      DLX_INST_CONTROL_UNIT_n84, DLX_INST_CONTROL_UNIT_n83, 
      DLX_INST_CONTROL_UNIT_n82, DLX_INST_CONTROL_UNIT_n81, 
      DLX_INST_CONTROL_UNIT_n80, DLX_INST_CONTROL_UNIT_n79, 
      DLX_INST_CONTROL_UNIT_n78, DLX_INST_CONTROL_UNIT_n77, 
      DLX_INST_CONTROL_UNIT_n76, DLX_INST_CONTROL_UNIT_n75, 
      DLX_INST_CONTROL_UNIT_n74, DLX_INST_CONTROL_UNIT_n73, 
      DLX_INST_CONTROL_UNIT_n72, DLX_INST_CONTROL_UNIT_n71, 
      DLX_INST_CONTROL_UNIT_n70, DLX_INST_CONTROL_UNIT_n69, 
      DLX_INST_CONTROL_UNIT_n68, DLX_INST_CONTROL_UNIT_n67, 
      DLX_INST_CONTROL_UNIT_n66, DLX_INST_CONTROL_UNIT_n65, 
      DLX_INST_CONTROL_UNIT_n64, DLX_INST_CONTROL_UNIT_n63, 
      DLX_INST_CONTROL_UNIT_n62, DLX_INST_CONTROL_UNIT_n61, 
      DLX_INST_CONTROL_UNIT_n60, DLX_INST_CONTROL_UNIT_n59, 
      DLX_INST_CONTROL_UNIT_net1651, DLX_INST_CONTROL_UNIT_net1650, 
      DLX_INST_CONTROL_UNIT_net1649, DLX_INST_CONTROL_UNIT_aluOpcode_i_0_port, 
      DLX_INST_CONTROL_UNIT_aluOpcode_i_1_port, 
      DLX_INST_CONTROL_UNIT_aluOpcode_i_2_port, 
      DLX_INST_CONTROL_UNIT_aluOpcode_i_3_port, DLX_INST_CONTROL_UNIT_RF_WE, 
      DLX_INST_CONTROL_UNIT_WB_MUX_SEL, DLX_INST_CONTROL_UNIT_JUMP_EN, 
      DLX_INST_CONTROL_UNIT_LMD_LATCH_EN, DLX_INST_CONTROL_UNIT_DRAM_WE, 
      DLX_INST_CONTROL_UNIT_EQ_COND, DLX_INST_CONTROL_UNIT_ALU_OUTREG_EN, 
      DLX_INST_CONTROL_UNIT_MUXB_SEL, DLX_INST_CONTROL_UNIT_MUXA_SEL, 
      DLX_INST_CONTROL_UNIT_Logic1_port, DLX_INST_DATA_PATH_n4, 
      DLX_INST_DATA_PATH_n3, DLX_INST_DATA_PATH_ALU_OUT2s_0_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_1_port, DLX_INST_DATA_PATH_ALU_OUT2s_2_port,
      DLX_INST_DATA_PATH_ALU_OUT2s_3_port, DLX_INST_DATA_PATH_ALU_OUT2s_4_port,
      DLX_INST_DATA_PATH_ALU_OUT2s_5_port, DLX_INST_DATA_PATH_ALU_OUT2s_6_port,
      DLX_INST_DATA_PATH_ALU_OUT2s_7_port, DLX_INST_DATA_PATH_ALU_OUT2s_8_port,
      DLX_INST_DATA_PATH_ALU_OUT2s_9_port, DLX_INST_DATA_PATH_ALU_OUT2s_10_port
      , DLX_INST_DATA_PATH_ALU_OUT2s_11_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_12_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_13_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_14_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_15_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_16_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_17_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_18_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_19_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_20_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_21_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_22_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_23_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_24_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_25_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_26_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_27_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_28_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_29_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_30_port, 
      DLX_INST_DATA_PATH_ALU_OUT2s_31_port, DLX_INST_DATA_PATH_LMD_OUTs_0_port,
      DLX_INST_DATA_PATH_LMD_OUTs_1_port, DLX_INST_DATA_PATH_LMD_OUTs_2_port, 
      DLX_INST_DATA_PATH_LMD_OUTs_3_port, DLX_INST_DATA_PATH_LMD_OUTs_4_port, 
      DLX_INST_DATA_PATH_LMD_OUTs_5_port, DLX_INST_DATA_PATH_LMD_OUTs_6_port, 
      DLX_INST_DATA_PATH_LMD_OUTs_7_port, DLX_INST_DATA_PATH_LMD_OUTs_8_port, 
      DLX_INST_DATA_PATH_LMD_OUTs_9_port, DLX_INST_DATA_PATH_LMD_OUTs_10_port, 
      DLX_INST_DATA_PATH_LMD_OUTs_11_port, DLX_INST_DATA_PATH_LMD_OUTs_12_port,
      DLX_INST_DATA_PATH_LMD_OUTs_13_port, DLX_INST_DATA_PATH_LMD_OUTs_14_port,
      DLX_INST_DATA_PATH_LMD_OUTs_15_port, DLX_INST_DATA_PATH_LMD_OUTs_16_port,
      DLX_INST_DATA_PATH_LMD_OUTs_17_port, DLX_INST_DATA_PATH_LMD_OUTs_18_port,
      DLX_INST_DATA_PATH_LMD_OUTs_19_port, DLX_INST_DATA_PATH_LMD_OUTs_20_port,
      DLX_INST_DATA_PATH_LMD_OUTs_21_port, DLX_INST_DATA_PATH_LMD_OUTs_22_port,
      DLX_INST_DATA_PATH_LMD_OUTs_23_port, DLX_INST_DATA_PATH_LMD_OUTs_24_port,
      DLX_INST_DATA_PATH_LMD_OUTs_25_port, DLX_INST_DATA_PATH_LMD_OUTs_26_port,
      DLX_INST_DATA_PATH_LMD_OUTs_27_port, DLX_INST_DATA_PATH_LMD_OUTs_28_port,
      DLX_INST_DATA_PATH_LMD_OUTs_29_port, DLX_INST_DATA_PATH_LMD_OUTs_30_port,
      DLX_INST_DATA_PATH_LMD_OUTs_31_port, DLX_INST_DATA_PATH_IR_OUT3s_0_port, 
      DLX_INST_DATA_PATH_IR_OUT3s_1_port, DLX_INST_DATA_PATH_IR_OUT3s_2_port, 
      DLX_INST_DATA_PATH_IR_OUT3s_3_port, DLX_INST_DATA_PATH_IR_OUT3s_4_port, 
      DLX_INST_DATA_PATH_IR_OUT3s_5_port, DLX_INST_DATA_PATH_IR_OUT3s_6_port, 
      DLX_INST_DATA_PATH_IR_OUT3s_7_port, DLX_INST_DATA_PATH_IR_OUT3s_8_port, 
      DLX_INST_DATA_PATH_IR_OUT3s_9_port, DLX_INST_DATA_PATH_IR_OUT3s_10_port, 
      DLX_INST_DATA_PATH_IR_OUT3s_11_port, DLX_INST_DATA_PATH_IR_OUT3s_12_port,
      DLX_INST_DATA_PATH_IR_OUT3s_13_port, DLX_INST_DATA_PATH_IR_OUT3s_14_port,
      DLX_INST_DATA_PATH_IR_OUT3s_15_port, DLX_INST_DATA_PATH_IR_OUT3s_16_port,
      DLX_INST_DATA_PATH_IR_OUT3s_17_port, DLX_INST_DATA_PATH_IR_OUT3s_18_port,
      DLX_INST_DATA_PATH_IR_OUT3s_19_port, DLX_INST_DATA_PATH_IR_OUT3s_20_port,
      DLX_INST_DATA_PATH_IR_OUT3s_21_port, DLX_INST_DATA_PATH_IR_OUT3s_22_port,
      DLX_INST_DATA_PATH_IR_OUT3s_23_port, DLX_INST_DATA_PATH_IR_OUT3s_24_port,
      DLX_INST_DATA_PATH_IR_OUT3s_25_port, DLX_INST_DATA_PATH_IR_OUT3s_26_port,
      DLX_INST_DATA_PATH_IR_OUT3s_27_port, DLX_INST_DATA_PATH_IR_OUT3s_28_port,
      DLX_INST_DATA_PATH_IR_OUT3s_29_port, DLX_INST_DATA_PATH_IR_OUT3s_30_port,
      DLX_INST_DATA_PATH_IR_OUT3s_31_port, DLX_INST_DATA_PATH_COND_OUTs, 
      DLX_INST_DATA_PATH_NPC2_OUTs_0_port, DLX_INST_DATA_PATH_NPC2_OUTs_1_port,
      DLX_INST_DATA_PATH_NPC2_OUTs_2_port, DLX_INST_DATA_PATH_NPC2_OUTs_3_port,
      DLX_INST_DATA_PATH_NPC2_OUTs_4_port, DLX_INST_DATA_PATH_NPC2_OUTs_5_port,
      DLX_INST_DATA_PATH_NPC2_OUTs_6_port, DLX_INST_DATA_PATH_NPC2_OUTs_7_port,
      DLX_INST_DATA_PATH_NPC2_OUTs_8_port, DLX_INST_DATA_PATH_NPC2_OUTs_9_port,
      DLX_INST_DATA_PATH_NPC2_OUTs_10_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_11_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_12_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_13_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_14_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_15_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_16_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_17_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_18_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_19_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_20_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_21_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_22_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_23_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_24_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_25_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_26_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_27_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_28_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_29_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_30_port, 
      DLX_INST_DATA_PATH_NPC2_OUTs_31_port, DLX_INST_DATA_PATH_IR_OUT2s_0_port,
      DLX_INST_DATA_PATH_IR_OUT2s_1_port, DLX_INST_DATA_PATH_IR_OUT2s_2_port, 
      DLX_INST_DATA_PATH_IR_OUT2s_3_port, DLX_INST_DATA_PATH_IR_OUT2s_4_port, 
      DLX_INST_DATA_PATH_IR_OUT2s_5_port, DLX_INST_DATA_PATH_IR_OUT2s_6_port, 
      DLX_INST_DATA_PATH_IR_OUT2s_7_port, DLX_INST_DATA_PATH_IR_OUT2s_8_port, 
      DLX_INST_DATA_PATH_IR_OUT2s_9_port, DLX_INST_DATA_PATH_IR_OUT2s_10_port, 
      DLX_INST_DATA_PATH_IR_OUT2s_11_port, DLX_INST_DATA_PATH_IR_OUT2s_12_port,
      DLX_INST_DATA_PATH_IR_OUT2s_13_port, DLX_INST_DATA_PATH_IR_OUT2s_14_port,
      DLX_INST_DATA_PATH_IR_OUT2s_15_port, DLX_INST_DATA_PATH_IR_OUT2s_16_port,
      DLX_INST_DATA_PATH_IR_OUT2s_17_port, DLX_INST_DATA_PATH_IR_OUT2s_18_port,
      DLX_INST_DATA_PATH_IR_OUT2s_19_port, DLX_INST_DATA_PATH_IR_OUT2s_20_port,
      DLX_INST_DATA_PATH_IR_OUT2s_21_port, DLX_INST_DATA_PATH_IR_OUT2s_22_port,
      DLX_INST_DATA_PATH_IR_OUT2s_23_port, DLX_INST_DATA_PATH_IR_OUT2s_24_port,
      DLX_INST_DATA_PATH_IR_OUT2s_25_port, DLX_INST_DATA_PATH_IR_OUT2s_26_port,
      DLX_INST_DATA_PATH_IR_OUT2s_27_port, DLX_INST_DATA_PATH_IR_OUT2s_28_port,
      DLX_INST_DATA_PATH_IR_OUT2s_29_port, DLX_INST_DATA_PATH_IR_OUT2s_30_port,
      DLX_INST_DATA_PATH_IR_OUT2s_31_port, DLX_INST_DATA_PATH_IR_OUT4s_0_port, 
      DLX_INST_DATA_PATH_IR_OUT4s_1_port, DLX_INST_DATA_PATH_IR_OUT4s_2_port, 
      DLX_INST_DATA_PATH_IR_OUT4s_3_port, DLX_INST_DATA_PATH_IR_OUT4s_4_port, 
      DLX_INST_DATA_PATH_IR_OUT4s_5_port, DLX_INST_DATA_PATH_IR_OUT4s_6_port, 
      DLX_INST_DATA_PATH_IR_OUT4s_7_port, DLX_INST_DATA_PATH_IR_OUT4s_8_port, 
      DLX_INST_DATA_PATH_IR_OUT4s_9_port, DLX_INST_DATA_PATH_IR_OUT4s_10_port, 
      DLX_INST_DATA_PATH_IR_OUT4s_11_port, DLX_INST_DATA_PATH_IR_OUT4s_12_port,
      DLX_INST_DATA_PATH_IR_OUT4s_13_port, DLX_INST_DATA_PATH_IR_OUT4s_14_port,
      DLX_INST_DATA_PATH_IR_OUT4s_15_port, DLX_INST_DATA_PATH_IR_OUT4s_16_port,
      DLX_INST_DATA_PATH_IR_OUT4s_17_port, DLX_INST_DATA_PATH_IR_OUT4s_18_port,
      DLX_INST_DATA_PATH_IR_OUT4s_19_port, DLX_INST_DATA_PATH_IR_OUT4s_20_port,
      DLX_INST_DATA_PATH_IR_OUT4s_21_port, DLX_INST_DATA_PATH_IR_OUT4s_22_port,
      DLX_INST_DATA_PATH_IR_OUT4s_23_port, DLX_INST_DATA_PATH_IR_OUT4s_24_port,
      DLX_INST_DATA_PATH_IR_OUT4s_25_port, DLX_INST_DATA_PATH_IR_OUT4s_26_port,
      DLX_INST_DATA_PATH_IR_OUT4s_27_port, DLX_INST_DATA_PATH_IR_OUT4s_28_port,
      DLX_INST_DATA_PATH_IR_OUT4s_29_port, DLX_INST_DATA_PATH_IR_OUT4s_30_port,
      DLX_INST_DATA_PATH_IR_OUT4s_31_port, DLX_INST_DATA_PATH_Imm_outs_0_port, 
      DLX_INST_DATA_PATH_Imm_outs_1_port, DLX_INST_DATA_PATH_Imm_outs_2_port, 
      DLX_INST_DATA_PATH_Imm_outs_3_port, DLX_INST_DATA_PATH_Imm_outs_4_port, 
      DLX_INST_DATA_PATH_Imm_outs_5_port, DLX_INST_DATA_PATH_Imm_outs_6_port, 
      DLX_INST_DATA_PATH_Imm_outs_7_port, DLX_INST_DATA_PATH_Imm_outs_8_port, 
      DLX_INST_DATA_PATH_Imm_outs_9_port, DLX_INST_DATA_PATH_Imm_outs_10_port, 
      DLX_INST_DATA_PATH_Imm_outs_11_port, DLX_INST_DATA_PATH_Imm_outs_12_port,
      DLX_INST_DATA_PATH_Imm_outs_13_port, DLX_INST_DATA_PATH_Imm_outs_14_port,
      DLX_INST_DATA_PATH_Imm_outs_15_port, DLX_INST_DATA_PATH_Imm_outs_16_port,
      DLX_INST_DATA_PATH_Imm_outs_17_port, DLX_INST_DATA_PATH_Imm_outs_18_port,
      DLX_INST_DATA_PATH_Imm_outs_19_port, DLX_INST_DATA_PATH_Imm_outs_20_port,
      DLX_INST_DATA_PATH_Imm_outs_21_port, DLX_INST_DATA_PATH_Imm_outs_22_port,
      DLX_INST_DATA_PATH_Imm_outs_23_port, DLX_INST_DATA_PATH_Imm_outs_24_port,
      DLX_INST_DATA_PATH_Imm_outs_25_port, DLX_INST_DATA_PATH_Imm_outs_26_port,
      DLX_INST_DATA_PATH_Imm_outs_27_port, DLX_INST_DATA_PATH_Imm_outs_28_port,
      DLX_INST_DATA_PATH_Imm_outs_29_port, DLX_INST_DATA_PATH_Imm_outs_30_port,
      DLX_INST_DATA_PATH_Imm_outs_31_port, DLX_INST_DATA_PATH_B_outs_0_port, 
      DLX_INST_DATA_PATH_B_outs_1_port, DLX_INST_DATA_PATH_B_outs_2_port, 
      DLX_INST_DATA_PATH_B_outs_3_port, DLX_INST_DATA_PATH_B_outs_4_port, 
      DLX_INST_DATA_PATH_B_outs_5_port, DLX_INST_DATA_PATH_B_outs_6_port, 
      DLX_INST_DATA_PATH_B_outs_7_port, DLX_INST_DATA_PATH_B_outs_8_port, 
      DLX_INST_DATA_PATH_B_outs_9_port, DLX_INST_DATA_PATH_B_outs_10_port, 
      DLX_INST_DATA_PATH_B_outs_11_port, DLX_INST_DATA_PATH_B_outs_12_port, 
      DLX_INST_DATA_PATH_B_outs_13_port, DLX_INST_DATA_PATH_B_outs_14_port, 
      DLX_INST_DATA_PATH_B_outs_15_port, DLX_INST_DATA_PATH_B_outs_16_port, 
      DLX_INST_DATA_PATH_B_outs_17_port, DLX_INST_DATA_PATH_B_outs_18_port, 
      DLX_INST_DATA_PATH_B_outs_19_port, DLX_INST_DATA_PATH_B_outs_20_port, 
      DLX_INST_DATA_PATH_B_outs_21_port, DLX_INST_DATA_PATH_B_outs_22_port, 
      DLX_INST_DATA_PATH_B_outs_23_port, DLX_INST_DATA_PATH_B_outs_24_port, 
      DLX_INST_DATA_PATH_B_outs_25_port, DLX_INST_DATA_PATH_B_outs_26_port, 
      DLX_INST_DATA_PATH_B_outs_27_port, DLX_INST_DATA_PATH_B_outs_28_port, 
      DLX_INST_DATA_PATH_B_outs_29_port, DLX_INST_DATA_PATH_B_outs_30_port, 
      DLX_INST_DATA_PATH_B_outs_31_port, DLX_INST_DATA_PATH_A_outs_0_port, 
      DLX_INST_DATA_PATH_A_outs_1_port, DLX_INST_DATA_PATH_A_outs_2_port, 
      DLX_INST_DATA_PATH_A_outs_3_port, DLX_INST_DATA_PATH_A_outs_4_port, 
      DLX_INST_DATA_PATH_A_outs_5_port, DLX_INST_DATA_PATH_A_outs_6_port, 
      DLX_INST_DATA_PATH_A_outs_7_port, DLX_INST_DATA_PATH_A_outs_8_port, 
      DLX_INST_DATA_PATH_A_outs_9_port, DLX_INST_DATA_PATH_A_outs_10_port, 
      DLX_INST_DATA_PATH_A_outs_11_port, DLX_INST_DATA_PATH_A_outs_12_port, 
      DLX_INST_DATA_PATH_A_outs_13_port, DLX_INST_DATA_PATH_A_outs_14_port, 
      DLX_INST_DATA_PATH_A_outs_15_port, DLX_INST_DATA_PATH_A_outs_16_port, 
      DLX_INST_DATA_PATH_A_outs_17_port, DLX_INST_DATA_PATH_A_outs_18_port, 
      DLX_INST_DATA_PATH_A_outs_19_port, DLX_INST_DATA_PATH_A_outs_20_port, 
      DLX_INST_DATA_PATH_A_outs_21_port, DLX_INST_DATA_PATH_A_outs_22_port, 
      DLX_INST_DATA_PATH_A_outs_23_port, DLX_INST_DATA_PATH_A_outs_24_port, 
      DLX_INST_DATA_PATH_A_outs_25_port, DLX_INST_DATA_PATH_A_outs_26_port, 
      DLX_INST_DATA_PATH_A_outs_27_port, DLX_INST_DATA_PATH_A_outs_28_port, 
      DLX_INST_DATA_PATH_A_outs_29_port, DLX_INST_DATA_PATH_A_outs_30_port, 
      DLX_INST_DATA_PATH_A_outs_31_port, DLX_INST_DATA_PATH_DATAIN_RFs_0_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_1_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_2_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_3_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_4_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_5_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_6_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_7_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_8_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_9_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_10_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_11_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_12_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_13_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_14_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_15_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_16_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_17_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_18_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_19_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_20_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_21_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_22_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_23_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_24_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_25_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_26_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_27_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_28_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_29_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_30_port, 
      DLX_INST_DATA_PATH_DATAIN_RFs_31_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_0_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_1_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_2_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_3_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_4_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_5_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_6_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_7_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_8_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_9_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_10_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_11_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_12_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_13_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_14_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_15_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_16_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_17_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_18_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_19_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_20_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_21_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_22_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_23_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_24_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_25_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_26_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_27_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_28_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_29_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_30_port, 
      DLX_INST_DATA_PATH_ADDERPC_OUTs_31_port, 
      DLX_INST_DATA_PATH_NPC_OUTs_0_port, DLX_INST_DATA_PATH_NPC_OUTs_1_port, 
      DLX_INST_DATA_PATH_NPC_OUTs_2_port, DLX_INST_DATA_PATH_NPC_OUTs_3_port, 
      DLX_INST_DATA_PATH_NPC_OUTs_4_port, DLX_INST_DATA_PATH_NPC_OUTs_5_port, 
      DLX_INST_DATA_PATH_NPC_OUTs_6_port, DLX_INST_DATA_PATH_NPC_OUTs_7_port, 
      DLX_INST_DATA_PATH_NPC_OUTs_8_port, DLX_INST_DATA_PATH_NPC_OUTs_9_port, 
      DLX_INST_DATA_PATH_NPC_OUTs_10_port, DLX_INST_DATA_PATH_NPC_OUTs_11_port,
      DLX_INST_DATA_PATH_NPC_OUTs_12_port, DLX_INST_DATA_PATH_NPC_OUTs_13_port,
      DLX_INST_DATA_PATH_NPC_OUTs_14_port, DLX_INST_DATA_PATH_NPC_OUTs_15_port,
      DLX_INST_DATA_PATH_NPC_OUTs_16_port, DLX_INST_DATA_PATH_NPC_OUTs_17_port,
      DLX_INST_DATA_PATH_NPC_OUTs_18_port, DLX_INST_DATA_PATH_NPC_OUTs_19_port,
      DLX_INST_DATA_PATH_NPC_OUTs_20_port, DLX_INST_DATA_PATH_NPC_OUTs_21_port,
      DLX_INST_DATA_PATH_NPC_OUTs_22_port, DLX_INST_DATA_PATH_NPC_OUTs_23_port,
      DLX_INST_DATA_PATH_NPC_OUTs_24_port, DLX_INST_DATA_PATH_NPC_OUTs_25_port,
      DLX_INST_DATA_PATH_NPC_OUTs_26_port, DLX_INST_DATA_PATH_NPC_OUTs_27_port,
      DLX_INST_DATA_PATH_NPC_OUTs_28_port, DLX_INST_DATA_PATH_NPC_OUTs_29_port,
      DLX_INST_DATA_PATH_NPC_OUTs_30_port, DLX_INST_DATA_PATH_NPC_OUTs_31_port,
      DLX_INST_DATA_PATH_TO_PC_OUTs_0_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_1_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_2_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_3_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_4_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_5_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_6_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_7_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_8_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_9_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_10_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_11_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_12_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_13_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_14_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_15_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_16_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_17_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_18_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_19_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_20_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_21_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_22_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_23_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_24_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_25_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_26_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_27_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_28_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_29_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_30_port, 
      DLX_INST_DATA_PATH_TO_PC_OUTs_31_port, DLX_INST_DATA_PATH_FETCH_n4, 
      DLX_INST_DATA_PATH_FETCH_n3, DLX_INST_DATA_PATH_FETCH_Logic0_port, 
      DLX_INST_DATA_PATH_FETCH_Logic1_port, DLX_INST_DATA_PATH_FETCH_ADD_n346, 
      DLX_INST_DATA_PATH_FETCH_ADD_n345, DLX_INST_DATA_PATH_FETCH_ADD_n344, 
      DLX_INST_DATA_PATH_FETCH_ADD_n343, DLX_INST_DATA_PATH_FETCH_ADD_n342, 
      DLX_INST_DATA_PATH_FETCH_ADD_n341, DLX_INST_DATA_PATH_FETCH_ADD_n340, 
      DLX_INST_DATA_PATH_FETCH_ADD_n339, DLX_INST_DATA_PATH_FETCH_ADD_n338, 
      DLX_INST_DATA_PATH_FETCH_ADD_n337, DLX_INST_DATA_PATH_FETCH_ADD_n336, 
      DLX_INST_DATA_PATH_FETCH_ADD_n335, DLX_INST_DATA_PATH_FETCH_ADD_n334, 
      DLX_INST_DATA_PATH_FETCH_ADD_n333, DLX_INST_DATA_PATH_FETCH_ADD_n332, 
      DLX_INST_DATA_PATH_FETCH_ADD_n331, DLX_INST_DATA_PATH_FETCH_ADD_n330, 
      DLX_INST_DATA_PATH_FETCH_ADD_n329, DLX_INST_DATA_PATH_FETCH_ADD_n328, 
      DLX_INST_DATA_PATH_FETCH_ADD_n327, DLX_INST_DATA_PATH_FETCH_ADD_n326, 
      DLX_INST_DATA_PATH_FETCH_ADD_n325, DLX_INST_DATA_PATH_FETCH_ADD_n324, 
      DLX_INST_DATA_PATH_FETCH_ADD_n323, DLX_INST_DATA_PATH_FETCH_ADD_n322, 
      DLX_INST_DATA_PATH_FETCH_ADD_n321, DLX_INST_DATA_PATH_FETCH_ADD_n320, 
      DLX_INST_DATA_PATH_FETCH_ADD_n319, DLX_INST_DATA_PATH_FETCH_ADD_n318, 
      DLX_INST_DATA_PATH_FETCH_ADD_n317, DLX_INST_DATA_PATH_FETCH_ADD_n316, 
      DLX_INST_DATA_PATH_FETCH_ADD_n315, DLX_INST_DATA_PATH_FETCH_ADD_n314, 
      DLX_INST_DATA_PATH_FETCH_ADD_n313, DLX_INST_DATA_PATH_FETCH_ADD_n312, 
      DLX_INST_DATA_PATH_FETCH_ADD_n311, DLX_INST_DATA_PATH_FETCH_ADD_n310, 
      DLX_INST_DATA_PATH_FETCH_ADD_n309, DLX_INST_DATA_PATH_FETCH_ADD_n308, 
      DLX_INST_DATA_PATH_FETCH_ADD_n307, DLX_INST_DATA_PATH_FETCH_ADD_n306, 
      DLX_INST_DATA_PATH_FETCH_ADD_n305, DLX_INST_DATA_PATH_FETCH_ADD_n304, 
      DLX_INST_DATA_PATH_FETCH_ADD_n303, DLX_INST_DATA_PATH_FETCH_ADD_n302, 
      DLX_INST_DATA_PATH_FETCH_ADD_n301, DLX_INST_DATA_PATH_FETCH_ADD_n300, 
      DLX_INST_DATA_PATH_FETCH_ADD_n299, DLX_INST_DATA_PATH_FETCH_ADD_n298, 
      DLX_INST_DATA_PATH_FETCH_ADD_n297, DLX_INST_DATA_PATH_FETCH_ADD_n296, 
      DLX_INST_DATA_PATH_FETCH_ADD_n295, DLX_INST_DATA_PATH_FETCH_ADD_n294, 
      DLX_INST_DATA_PATH_FETCH_ADD_n293, DLX_INST_DATA_PATH_FETCH_ADD_n292, 
      DLX_INST_DATA_PATH_FETCH_ADD_n291, DLX_INST_DATA_PATH_FETCH_ADD_n290, 
      DLX_INST_DATA_PATH_FETCH_ADD_n289, DLX_INST_DATA_PATH_FETCH_ADD_n288, 
      DLX_INST_DATA_PATH_FETCH_ADD_n287, DLX_INST_DATA_PATH_FETCH_ADD_n286, 
      DLX_INST_DATA_PATH_FETCH_ADD_n285, DLX_INST_DATA_PATH_FETCH_ADD_n284, 
      DLX_INST_DATA_PATH_FETCH_ADD_n283, DLX_INST_DATA_PATH_FETCH_ADD_n282, 
      DLX_INST_DATA_PATH_FETCH_ADD_n281, DLX_INST_DATA_PATH_FETCH_ADD_n280, 
      DLX_INST_DATA_PATH_FETCH_ADD_n279, DLX_INST_DATA_PATH_FETCH_ADD_n278, 
      DLX_INST_DATA_PATH_FETCH_ADD_n277, DLX_INST_DATA_PATH_FETCH_ADD_n276, 
      DLX_INST_DATA_PATH_FETCH_ADD_n275, DLX_INST_DATA_PATH_FETCH_ADD_n274, 
      DLX_INST_DATA_PATH_FETCH_ADD_n273, DLX_INST_DATA_PATH_FETCH_ADD_n272, 
      DLX_INST_DATA_PATH_FETCH_ADD_n271, DLX_INST_DATA_PATH_FETCH_ADD_n270, 
      DLX_INST_DATA_PATH_FETCH_ADD_n269, DLX_INST_DATA_PATH_FETCH_ADD_n268, 
      DLX_INST_DATA_PATH_FETCH_ADD_n267, DLX_INST_DATA_PATH_FETCH_ADD_n266, 
      DLX_INST_DATA_PATH_FETCH_ADD_n265, DLX_INST_DATA_PATH_FETCH_ADD_n264, 
      DLX_INST_DATA_PATH_FETCH_ADD_n263, DLX_INST_DATA_PATH_FETCH_ADD_n262, 
      DLX_INST_DATA_PATH_FETCH_ADD_n261, DLX_INST_DATA_PATH_FETCH_ADD_n260, 
      DLX_INST_DATA_PATH_FETCH_ADD_n259, DLX_INST_DATA_PATH_FETCH_ADD_n258, 
      DLX_INST_DATA_PATH_FETCH_ADD_n257, DLX_INST_DATA_PATH_FETCH_ADD_n256, 
      DLX_INST_DATA_PATH_FETCH_ADD_n255, DLX_INST_DATA_PATH_FETCH_ADD_n254, 
      DLX_INST_DATA_PATH_FETCH_ADD_n253, DLX_INST_DATA_PATH_FETCH_ADD_n252, 
      DLX_INST_DATA_PATH_FETCH_ADD_n251, DLX_INST_DATA_PATH_FETCH_ADD_n250, 
      DLX_INST_DATA_PATH_FETCH_ADD_n249, DLX_INST_DATA_PATH_FETCH_ADD_n248, 
      DLX_INST_DATA_PATH_FETCH_ADD_n247, DLX_INST_DATA_PATH_FETCH_ADD_n246, 
      DLX_INST_DATA_PATH_FETCH_ADD_n245, DLX_INST_DATA_PATH_FETCH_ADD_n244, 
      DLX_INST_DATA_PATH_FETCH_ADD_n243, DLX_INST_DATA_PATH_FETCH_ADD_n242, 
      DLX_INST_DATA_PATH_FETCH_ADD_n241, DLX_INST_DATA_PATH_FETCH_ADD_n240, 
      DLX_INST_DATA_PATH_FETCH_ADD_n239, DLX_INST_DATA_PATH_FETCH_ADD_n238, 
      DLX_INST_DATA_PATH_FETCH_ADD_n237, DLX_INST_DATA_PATH_FETCH_ADD_n236, 
      DLX_INST_DATA_PATH_FETCH_ADD_n235, DLX_INST_DATA_PATH_FETCH_ADD_n234, 
      DLX_INST_DATA_PATH_FETCH_ADD_n233, DLX_INST_DATA_PATH_FETCH_ADD_n232, 
      DLX_INST_DATA_PATH_FETCH_ADD_n231, DLX_INST_DATA_PATH_FETCH_ADD_n230, 
      DLX_INST_DATA_PATH_FETCH_ADD_n229, DLX_INST_DATA_PATH_FETCH_ADD_n228, 
      DLX_INST_DATA_PATH_FETCH_ADD_n227, DLX_INST_DATA_PATH_FETCH_ADD_n226, 
      DLX_INST_DATA_PATH_FETCH_ADD_n225, DLX_INST_DATA_PATH_FETCH_ADD_n224, 
      DLX_INST_DATA_PATH_FETCH_ADD_n223, DLX_INST_DATA_PATH_FETCH_ADD_n222, 
      DLX_INST_DATA_PATH_FETCH_ADD_n221, DLX_INST_DATA_PATH_FETCH_ADD_n220, 
      DLX_INST_DATA_PATH_FETCH_ADD_n219, DLX_INST_DATA_PATH_FETCH_ADD_n218, 
      DLX_INST_DATA_PATH_FETCH_ADD_n217, DLX_INST_DATA_PATH_FETCH_ADD_n216, 
      DLX_INST_DATA_PATH_FETCH_ADD_n215, DLX_INST_DATA_PATH_FETCH_ADD_n214, 
      DLX_INST_DATA_PATH_FETCH_ADD_n213, DLX_INST_DATA_PATH_FETCH_ADD_n212, 
      DLX_INST_DATA_PATH_FETCH_ADD_n211, DLX_INST_DATA_PATH_FETCH_ADD_n210, 
      DLX_INST_DATA_PATH_FETCH_ADD_n209, DLX_INST_DATA_PATH_FETCH_ADD_n208, 
      DLX_INST_DATA_PATH_FETCH_ADD_n207, DLX_INST_DATA_PATH_FETCH_ADD_n206, 
      DLX_INST_DATA_PATH_FETCH_ADD_n205, DLX_INST_DATA_PATH_FETCH_ADD_n204, 
      DLX_INST_DATA_PATH_FETCH_ADD_n203, DLX_INST_DATA_PATH_FETCH_ADD_n202, 
      DLX_INST_DATA_PATH_FETCH_ADD_n201, DLX_INST_DATA_PATH_FETCH_ADD_n200, 
      DLX_INST_DATA_PATH_FETCH_ADD_n199, DLX_INST_DATA_PATH_FETCH_ADD_n198, 
      DLX_INST_DATA_PATH_FETCH_ADD_n197, DLX_INST_DATA_PATH_FETCH_ADD_n196, 
      DLX_INST_DATA_PATH_FETCH_ADD_n195, DLX_INST_DATA_PATH_FETCH_ADD_n194, 
      DLX_INST_DATA_PATH_FETCH_ADD_n193, DLX_INST_DATA_PATH_FETCH_ADD_n192, 
      DLX_INST_DATA_PATH_FETCH_ADD_n191, DLX_INST_DATA_PATH_FETCH_ADD_n190, 
      DLX_INST_DATA_PATH_FETCH_ADD_n189, DLX_INST_DATA_PATH_FETCH_ADD_n188, 
      DLX_INST_DATA_PATH_FETCH_ADD_n187, DLX_INST_DATA_PATH_FETCH_ADD_n186, 
      DLX_INST_DATA_PATH_FETCH_ADD_n185, DLX_INST_DATA_PATH_FETCH_ADD_n184, 
      DLX_INST_DATA_PATH_FETCH_ADD_n183, DLX_INST_DATA_PATH_FETCH_ADD_n182, 
      DLX_INST_DATA_PATH_FETCH_ADD_n181, DLX_INST_DATA_PATH_FETCH_ADD_n180, 
      DLX_INST_DATA_PATH_FETCH_ADD_n179, DLX_INST_DATA_PATH_FETCH_ADD_n178, 
      DLX_INST_DATA_PATH_FETCH_ADD_n177, DLX_INST_DATA_PATH_FETCH_ADD_n176, 
      DLX_INST_DATA_PATH_FETCH_ADD_n175, DLX_INST_DATA_PATH_FETCH_ADD_Co, 
      DLX_INST_DATA_PATH_FETCH_PC_n16, DLX_INST_DATA_PATH_FETCH_PC_n15, 
      DLX_INST_DATA_PATH_FETCH_PC_n14, DLX_INST_DATA_PATH_FETCH_PC_n13, 
      DLX_INST_DATA_PATH_FETCH_PC_n12, DLX_INST_DATA_PATH_FETCH_PC_n11, 
      DLX_INST_DATA_PATH_FETCH_PC_n10, DLX_INST_DATA_PATH_FETCH_PC_n9, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_0_n2, DLX_INST_DATA_PATH_FETCH_PC_FF_0_n1,
      DLX_INST_DATA_PATH_FETCH_PC_FF_1_n2, DLX_INST_DATA_PATH_FETCH_PC_FF_1_n1,
      DLX_INST_DATA_PATH_FETCH_PC_FF_2_n2, DLX_INST_DATA_PATH_FETCH_PC_FF_2_n1,
      DLX_INST_DATA_PATH_FETCH_PC_FF_3_n2, DLX_INST_DATA_PATH_FETCH_PC_FF_3_n1,
      DLX_INST_DATA_PATH_FETCH_PC_FF_4_n2, DLX_INST_DATA_PATH_FETCH_PC_FF_4_n1,
      DLX_INST_DATA_PATH_FETCH_PC_FF_5_n2, DLX_INST_DATA_PATH_FETCH_PC_FF_5_n1,
      DLX_INST_DATA_PATH_FETCH_PC_FF_6_n2, DLX_INST_DATA_PATH_FETCH_PC_FF_6_n1,
      DLX_INST_DATA_PATH_FETCH_PC_FF_7_n2, DLX_INST_DATA_PATH_FETCH_PC_FF_7_n1,
      DLX_INST_DATA_PATH_FETCH_PC_FF_8_n2, DLX_INST_DATA_PATH_FETCH_PC_FF_8_n1,
      DLX_INST_DATA_PATH_FETCH_PC_FF_9_n2, DLX_INST_DATA_PATH_FETCH_PC_FF_9_n1,
      DLX_INST_DATA_PATH_FETCH_PC_FF_10_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_10_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_11_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_11_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_12_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_12_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_13_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_13_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_14_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_14_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_15_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_15_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_16_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_16_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_17_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_17_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_18_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_18_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_19_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_19_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_20_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_20_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_21_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_21_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_22_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_22_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_23_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_23_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_24_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_24_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_25_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_25_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_26_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_26_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_27_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_27_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_28_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_28_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_29_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_29_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_30_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_30_n1, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_31_n2, 
      DLX_INST_DATA_PATH_FETCH_PC_FF_31_n1, DLX_INST_DATA_PATH_FETCH_IR_n16, 
      DLX_INST_DATA_PATH_FETCH_IR_n15, DLX_INST_DATA_PATH_FETCH_IR_n14, 
      DLX_INST_DATA_PATH_FETCH_IR_n13, DLX_INST_DATA_PATH_FETCH_IR_n12, 
      DLX_INST_DATA_PATH_FETCH_IR_n11, DLX_INST_DATA_PATH_FETCH_IR_n10, 
      DLX_INST_DATA_PATH_FETCH_IR_n9, DLX_INST_DATA_PATH_FETCH_IR_FF_0_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_0_n1, DLX_INST_DATA_PATH_FETCH_IR_FF_1_n2,
      DLX_INST_DATA_PATH_FETCH_IR_FF_1_n1, DLX_INST_DATA_PATH_FETCH_IR_FF_2_n2,
      DLX_INST_DATA_PATH_FETCH_IR_FF_2_n1, DLX_INST_DATA_PATH_FETCH_IR_FF_3_n2,
      DLX_INST_DATA_PATH_FETCH_IR_FF_3_n1, DLX_INST_DATA_PATH_FETCH_IR_FF_4_n2,
      DLX_INST_DATA_PATH_FETCH_IR_FF_4_n1, DLX_INST_DATA_PATH_FETCH_IR_FF_5_n2,
      DLX_INST_DATA_PATH_FETCH_IR_FF_5_n1, DLX_INST_DATA_PATH_FETCH_IR_FF_6_n2,
      DLX_INST_DATA_PATH_FETCH_IR_FF_6_n1, DLX_INST_DATA_PATH_FETCH_IR_FF_7_n2,
      DLX_INST_DATA_PATH_FETCH_IR_FF_7_n1, DLX_INST_DATA_PATH_FETCH_IR_FF_8_n2,
      DLX_INST_DATA_PATH_FETCH_IR_FF_8_n1, DLX_INST_DATA_PATH_FETCH_IR_FF_9_n2,
      DLX_INST_DATA_PATH_FETCH_IR_FF_9_n1, DLX_INST_DATA_PATH_FETCH_IR_FF_10_n2
      , DLX_INST_DATA_PATH_FETCH_IR_FF_10_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_11_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_11_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_12_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_12_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_13_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_13_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_14_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_14_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_15_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_15_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_16_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_16_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_17_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_17_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_18_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_18_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_19_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_19_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_20_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_20_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_21_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_21_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_22_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_22_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_23_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_23_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_24_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_24_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_25_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_25_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_26_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_26_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_27_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_27_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_28_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_28_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_29_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_29_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_30_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_30_n1, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_31_n2, 
      DLX_INST_DATA_PATH_FETCH_IR_FF_31_n1, DLX_INST_DATA_PATH_FETCH_NPC_n16, 
      DLX_INST_DATA_PATH_FETCH_NPC_n15, DLX_INST_DATA_PATH_FETCH_NPC_n14, 
      DLX_INST_DATA_PATH_FETCH_NPC_n13, DLX_INST_DATA_PATH_FETCH_NPC_n12, 
      DLX_INST_DATA_PATH_FETCH_NPC_n11, DLX_INST_DATA_PATH_FETCH_NPC_n10, 
      DLX_INST_DATA_PATH_FETCH_NPC_n9, DLX_INST_DATA_PATH_FETCH_NPC_FF_0_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_0_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_1_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_1_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_2_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_2_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_3_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_3_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_4_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_4_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_5_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_5_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_6_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_6_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_7_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_7_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_8_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_8_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_9_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_9_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_10_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_10_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_11_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_11_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_12_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_12_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_13_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_13_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_14_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_14_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_15_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_15_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_16_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_16_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_17_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_17_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_18_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_18_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_19_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_19_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_20_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_20_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_21_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_21_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_22_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_22_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_23_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_23_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_24_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_24_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_25_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_25_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_26_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_26_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_27_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_27_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_28_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_28_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_29_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_29_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_30_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_30_n1, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_31_n2, 
      DLX_INST_DATA_PATH_FETCH_NPC_FF_31_n1, DLX_INST_DATA_PATH_DECODE_n13, 
      DLX_INST_DATA_PATH_DECODE_n12, DLX_INST_DATA_PATH_DECODE_n11, 
      DLX_INST_DATA_PATH_DECODE_n10, DLX_INST_DATA_PATH_DECODE_n5, 
      DLX_INST_DATA_PATH_DECODE_n4, DLX_INST_DATA_PATH_DECODE_n3, 
      DLX_INST_DATA_PATH_DECODE_n2, DLX_INST_DATA_PATH_DECODE_n1, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_0_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_1_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_2_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_3_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_4_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_5_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_6_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_7_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_8_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_9_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_10_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_11_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_12_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_13_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_14_port, 
      DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, 
      DLX_INST_DATA_PATH_DECODE_Logic1_port, DLX_INST_DATA_PATH_DECODE_NPC2_n16
      , DLX_INST_DATA_PATH_DECODE_NPC2_n15, DLX_INST_DATA_PATH_DECODE_NPC2_n14,
      DLX_INST_DATA_PATH_DECODE_NPC2_n13, DLX_INST_DATA_PATH_DECODE_NPC2_n12, 
      DLX_INST_DATA_PATH_DECODE_NPC2_n11, DLX_INST_DATA_PATH_DECODE_NPC2_n10, 
      DLX_INST_DATA_PATH_DECODE_NPC2_n9, DLX_INST_DATA_PATH_DECODE_NPC2_FF_0_n2
      , DLX_INST_DATA_PATH_DECODE_NPC2_FF_0_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_1_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_1_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_2_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_2_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_3_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_3_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_4_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_4_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_5_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_5_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_6_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_6_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_7_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_7_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_8_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_8_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_9_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_9_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_10_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_10_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_11_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_11_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_12_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_12_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_13_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_13_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_14_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_14_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_15_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_15_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_16_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_16_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_17_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_17_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_18_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_18_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_19_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_19_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_20_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_20_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_21_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_21_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_22_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_22_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_23_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_23_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_24_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_24_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_25_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_25_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_26_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_26_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_27_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_27_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_28_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_28_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_29_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_29_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_30_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_30_n1, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_31_n2, 
      DLX_INST_DATA_PATH_DECODE_NPC2_FF_31_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_n16, DLX_INST_DATA_PATH_DECODE_Imm_n15, 
      DLX_INST_DATA_PATH_DECODE_Imm_n14, DLX_INST_DATA_PATH_DECODE_Imm_n13, 
      DLX_INST_DATA_PATH_DECODE_Imm_n12, DLX_INST_DATA_PATH_DECODE_Imm_n11, 
      DLX_INST_DATA_PATH_DECODE_Imm_n10, DLX_INST_DATA_PATH_DECODE_Imm_n9, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_0_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_0_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_1_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_1_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_2_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_2_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_3_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_3_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_4_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_4_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_5_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_5_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_6_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_6_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_7_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_7_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_8_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_8_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_9_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_9_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_10_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_10_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_11_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_11_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_12_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_12_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_13_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_13_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_14_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_14_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_15_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_15_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_16_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_16_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_17_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_17_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_18_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_18_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_19_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_19_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_20_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_20_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_21_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_21_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_22_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_22_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_23_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_23_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_24_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_24_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_25_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_25_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_26_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_26_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_27_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_27_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_28_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_28_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_29_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_29_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_30_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_30_n1, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_31_n2, 
      DLX_INST_DATA_PATH_DECODE_Imm_FF_31_n1, DLX_INST_DATA_PATH_DECODE_IR2_n16
      , DLX_INST_DATA_PATH_DECODE_IR2_n15, DLX_INST_DATA_PATH_DECODE_IR2_n14, 
      DLX_INST_DATA_PATH_DECODE_IR2_n13, DLX_INST_DATA_PATH_DECODE_IR2_n12, 
      DLX_INST_DATA_PATH_DECODE_IR2_n11, DLX_INST_DATA_PATH_DECODE_IR2_n10, 
      DLX_INST_DATA_PATH_DECODE_IR2_n9, DLX_INST_DATA_PATH_DECODE_IR2_FF_0_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_0_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_1_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_1_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_2_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_2_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_3_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_3_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_4_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_4_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_5_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_5_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_6_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_6_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_7_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_7_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_8_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_8_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_9_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_9_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_10_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_10_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_11_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_11_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_12_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_12_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_13_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_13_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_14_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_14_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_15_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_15_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_16_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_16_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_17_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_17_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_18_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_18_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_19_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_19_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_20_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_20_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_21_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_21_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_22_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_22_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_23_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_23_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_24_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_24_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_25_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_25_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_26_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_26_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_27_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_27_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_28_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_28_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_29_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_29_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_30_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_30_n1, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_31_n2, 
      DLX_INST_DATA_PATH_DECODE_IR2_FF_31_n1, 
      DLX_INST_DATA_PATH_DECODE_RF_n7087, DLX_INST_DATA_PATH_DECODE_RF_n7086, 
      DLX_INST_DATA_PATH_DECODE_RF_n7085, DLX_INST_DATA_PATH_DECODE_RF_n7084, 
      DLX_INST_DATA_PATH_DECODE_RF_n7083, DLX_INST_DATA_PATH_DECODE_RF_n7082, 
      DLX_INST_DATA_PATH_DECODE_RF_n7081, DLX_INST_DATA_PATH_DECODE_RF_n7080, 
      DLX_INST_DATA_PATH_DECODE_RF_n7079, DLX_INST_DATA_PATH_DECODE_RF_n7078, 
      DLX_INST_DATA_PATH_DECODE_RF_n7077, DLX_INST_DATA_PATH_DECODE_RF_n7076, 
      DLX_INST_DATA_PATH_DECODE_RF_n7075, DLX_INST_DATA_PATH_DECODE_RF_n7074, 
      DLX_INST_DATA_PATH_DECODE_RF_n7073, DLX_INST_DATA_PATH_DECODE_RF_n7072, 
      DLX_INST_DATA_PATH_DECODE_RF_n7071, DLX_INST_DATA_PATH_DECODE_RF_n7070, 
      DLX_INST_DATA_PATH_DECODE_RF_n7069, DLX_INST_DATA_PATH_DECODE_RF_n7068, 
      DLX_INST_DATA_PATH_DECODE_RF_n7067, DLX_INST_DATA_PATH_DECODE_RF_n7066, 
      DLX_INST_DATA_PATH_DECODE_RF_n7065, DLX_INST_DATA_PATH_DECODE_RF_n7064, 
      DLX_INST_DATA_PATH_DECODE_RF_n7063, DLX_INST_DATA_PATH_DECODE_RF_n7062, 
      DLX_INST_DATA_PATH_DECODE_RF_n7061, DLX_INST_DATA_PATH_DECODE_RF_n7060, 
      DLX_INST_DATA_PATH_DECODE_RF_n7059, DLX_INST_DATA_PATH_DECODE_RF_n7058, 
      DLX_INST_DATA_PATH_DECODE_RF_n7057, DLX_INST_DATA_PATH_DECODE_RF_n7056, 
      DLX_INST_DATA_PATH_DECODE_RF_n7055, DLX_INST_DATA_PATH_DECODE_RF_n7054, 
      DLX_INST_DATA_PATH_DECODE_RF_n7053, DLX_INST_DATA_PATH_DECODE_RF_n7052, 
      DLX_INST_DATA_PATH_DECODE_RF_n7051, DLX_INST_DATA_PATH_DECODE_RF_n7050, 
      DLX_INST_DATA_PATH_DECODE_RF_n7049, DLX_INST_DATA_PATH_DECODE_RF_n7048, 
      DLX_INST_DATA_PATH_DECODE_RF_n7047, DLX_INST_DATA_PATH_DECODE_RF_n7046, 
      DLX_INST_DATA_PATH_DECODE_RF_n7045, DLX_INST_DATA_PATH_DECODE_RF_n7044, 
      DLX_INST_DATA_PATH_DECODE_RF_n7043, DLX_INST_DATA_PATH_DECODE_RF_n7042, 
      DLX_INST_DATA_PATH_DECODE_RF_n7041, DLX_INST_DATA_PATH_DECODE_RF_n7040, 
      DLX_INST_DATA_PATH_DECODE_RF_n7039, DLX_INST_DATA_PATH_DECODE_RF_n7038, 
      DLX_INST_DATA_PATH_DECODE_RF_n7037, DLX_INST_DATA_PATH_DECODE_RF_n7036, 
      DLX_INST_DATA_PATH_DECODE_RF_n7035, DLX_INST_DATA_PATH_DECODE_RF_n7034, 
      DLX_INST_DATA_PATH_DECODE_RF_n7033, DLX_INST_DATA_PATH_DECODE_RF_n7032, 
      DLX_INST_DATA_PATH_DECODE_RF_n7031, DLX_INST_DATA_PATH_DECODE_RF_n7030, 
      DLX_INST_DATA_PATH_DECODE_RF_n7029, DLX_INST_DATA_PATH_DECODE_RF_n7028, 
      DLX_INST_DATA_PATH_DECODE_RF_n7027, DLX_INST_DATA_PATH_DECODE_RF_n7026, 
      DLX_INST_DATA_PATH_DECODE_RF_n7025, DLX_INST_DATA_PATH_DECODE_RF_n7024, 
      DLX_INST_DATA_PATH_DECODE_RF_n7023, DLX_INST_DATA_PATH_DECODE_RF_n7022, 
      DLX_INST_DATA_PATH_DECODE_RF_n7021, DLX_INST_DATA_PATH_DECODE_RF_n7020, 
      DLX_INST_DATA_PATH_DECODE_RF_n7019, DLX_INST_DATA_PATH_DECODE_RF_n7018, 
      DLX_INST_DATA_PATH_DECODE_RF_n7017, DLX_INST_DATA_PATH_DECODE_RF_n7016, 
      DLX_INST_DATA_PATH_DECODE_RF_n7015, DLX_INST_DATA_PATH_DECODE_RF_n7014, 
      DLX_INST_DATA_PATH_DECODE_RF_n7013, DLX_INST_DATA_PATH_DECODE_RF_n7012, 
      DLX_INST_DATA_PATH_DECODE_RF_n7011, DLX_INST_DATA_PATH_DECODE_RF_n7010, 
      DLX_INST_DATA_PATH_DECODE_RF_n7009, DLX_INST_DATA_PATH_DECODE_RF_n7008, 
      DLX_INST_DATA_PATH_DECODE_RF_n7007, DLX_INST_DATA_PATH_DECODE_RF_n7006, 
      DLX_INST_DATA_PATH_DECODE_RF_n7005, DLX_INST_DATA_PATH_DECODE_RF_n7004, 
      DLX_INST_DATA_PATH_DECODE_RF_n7003, DLX_INST_DATA_PATH_DECODE_RF_n7002, 
      DLX_INST_DATA_PATH_DECODE_RF_n7001, DLX_INST_DATA_PATH_DECODE_RF_n7000, 
      DLX_INST_DATA_PATH_DECODE_RF_n6999, DLX_INST_DATA_PATH_DECODE_RF_n6998, 
      DLX_INST_DATA_PATH_DECODE_RF_n6997, DLX_INST_DATA_PATH_DECODE_RF_n6996, 
      DLX_INST_DATA_PATH_DECODE_RF_n6995, DLX_INST_DATA_PATH_DECODE_RF_n6994, 
      DLX_INST_DATA_PATH_DECODE_RF_n6993, DLX_INST_DATA_PATH_DECODE_RF_n6992, 
      DLX_INST_DATA_PATH_DECODE_RF_n6991, DLX_INST_DATA_PATH_DECODE_RF_n6990, 
      DLX_INST_DATA_PATH_DECODE_RF_n6989, DLX_INST_DATA_PATH_DECODE_RF_n6988, 
      DLX_INST_DATA_PATH_DECODE_RF_n6987, DLX_INST_DATA_PATH_DECODE_RF_n6986, 
      DLX_INST_DATA_PATH_DECODE_RF_n6985, DLX_INST_DATA_PATH_DECODE_RF_n6984, 
      DLX_INST_DATA_PATH_DECODE_RF_n6983, DLX_INST_DATA_PATH_DECODE_RF_n6982, 
      DLX_INST_DATA_PATH_DECODE_RF_n6981, DLX_INST_DATA_PATH_DECODE_RF_n6980, 
      DLX_INST_DATA_PATH_DECODE_RF_n6979, DLX_INST_DATA_PATH_DECODE_RF_n6978, 
      DLX_INST_DATA_PATH_DECODE_RF_n6977, DLX_INST_DATA_PATH_DECODE_RF_n6976, 
      DLX_INST_DATA_PATH_DECODE_RF_n6975, DLX_INST_DATA_PATH_DECODE_RF_n6974, 
      DLX_INST_DATA_PATH_DECODE_RF_n6973, DLX_INST_DATA_PATH_DECODE_RF_n6972, 
      DLX_INST_DATA_PATH_DECODE_RF_n6971, DLX_INST_DATA_PATH_DECODE_RF_n6970, 
      DLX_INST_DATA_PATH_DECODE_RF_n6969, DLX_INST_DATA_PATH_DECODE_RF_n6968, 
      DLX_INST_DATA_PATH_DECODE_RF_n6967, DLX_INST_DATA_PATH_DECODE_RF_n6966, 
      DLX_INST_DATA_PATH_DECODE_RF_n6965, DLX_INST_DATA_PATH_DECODE_RF_n6964, 
      DLX_INST_DATA_PATH_DECODE_RF_n6963, DLX_INST_DATA_PATH_DECODE_RF_n6962, 
      DLX_INST_DATA_PATH_DECODE_RF_n6961, DLX_INST_DATA_PATH_DECODE_RF_n6960, 
      DLX_INST_DATA_PATH_DECODE_RF_n6959, DLX_INST_DATA_PATH_DECODE_RF_n6958, 
      DLX_INST_DATA_PATH_DECODE_RF_n6957, DLX_INST_DATA_PATH_DECODE_RF_n6956, 
      DLX_INST_DATA_PATH_DECODE_RF_n6955, DLX_INST_DATA_PATH_DECODE_RF_n6954, 
      DLX_INST_DATA_PATH_DECODE_RF_n6953, DLX_INST_DATA_PATH_DECODE_RF_n6952, 
      DLX_INST_DATA_PATH_DECODE_RF_n6951, DLX_INST_DATA_PATH_DECODE_RF_n6950, 
      DLX_INST_DATA_PATH_DECODE_RF_n6949, DLX_INST_DATA_PATH_DECODE_RF_n6948, 
      DLX_INST_DATA_PATH_DECODE_RF_n6947, DLX_INST_DATA_PATH_DECODE_RF_n6946, 
      DLX_INST_DATA_PATH_DECODE_RF_n6945, DLX_INST_DATA_PATH_DECODE_RF_n6944, 
      DLX_INST_DATA_PATH_DECODE_RF_n6943, DLX_INST_DATA_PATH_DECODE_RF_n6942, 
      DLX_INST_DATA_PATH_DECODE_RF_n6941, DLX_INST_DATA_PATH_DECODE_RF_n6940, 
      DLX_INST_DATA_PATH_DECODE_RF_n6939, DLX_INST_DATA_PATH_DECODE_RF_n6938, 
      DLX_INST_DATA_PATH_DECODE_RF_n6937, DLX_INST_DATA_PATH_DECODE_RF_n6936, 
      DLX_INST_DATA_PATH_DECODE_RF_n6935, DLX_INST_DATA_PATH_DECODE_RF_n6934, 
      DLX_INST_DATA_PATH_DECODE_RF_n6933, DLX_INST_DATA_PATH_DECODE_RF_n6932, 
      DLX_INST_DATA_PATH_DECODE_RF_n6931, DLX_INST_DATA_PATH_DECODE_RF_n6930, 
      DLX_INST_DATA_PATH_DECODE_RF_n6929, DLX_INST_DATA_PATH_DECODE_RF_n6928, 
      DLX_INST_DATA_PATH_DECODE_RF_n6927, DLX_INST_DATA_PATH_DECODE_RF_n6926, 
      DLX_INST_DATA_PATH_DECODE_RF_n6925, DLX_INST_DATA_PATH_DECODE_RF_n6924, 
      DLX_INST_DATA_PATH_DECODE_RF_n6923, DLX_INST_DATA_PATH_DECODE_RF_n6922, 
      DLX_INST_DATA_PATH_DECODE_RF_n6921, DLX_INST_DATA_PATH_DECODE_RF_n6920, 
      DLX_INST_DATA_PATH_DECODE_RF_n6919, DLX_INST_DATA_PATH_DECODE_RF_n6918, 
      DLX_INST_DATA_PATH_DECODE_RF_n6917, DLX_INST_DATA_PATH_DECODE_RF_n6916, 
      DLX_INST_DATA_PATH_DECODE_RF_n6915, DLX_INST_DATA_PATH_DECODE_RF_n6914, 
      DLX_INST_DATA_PATH_DECODE_RF_n6913, DLX_INST_DATA_PATH_DECODE_RF_n6912, 
      DLX_INST_DATA_PATH_DECODE_RF_n6911, DLX_INST_DATA_PATH_DECODE_RF_n6910, 
      DLX_INST_DATA_PATH_DECODE_RF_n6909, DLX_INST_DATA_PATH_DECODE_RF_n6908, 
      DLX_INST_DATA_PATH_DECODE_RF_n6907, DLX_INST_DATA_PATH_DECODE_RF_n6906, 
      DLX_INST_DATA_PATH_DECODE_RF_n6905, DLX_INST_DATA_PATH_DECODE_RF_n6904, 
      DLX_INST_DATA_PATH_DECODE_RF_n6903, DLX_INST_DATA_PATH_DECODE_RF_n6902, 
      DLX_INST_DATA_PATH_DECODE_RF_n6901, DLX_INST_DATA_PATH_DECODE_RF_n6900, 
      DLX_INST_DATA_PATH_DECODE_RF_n6899, DLX_INST_DATA_PATH_DECODE_RF_n6898, 
      DLX_INST_DATA_PATH_DECODE_RF_n6897, DLX_INST_DATA_PATH_DECODE_RF_n6896, 
      DLX_INST_DATA_PATH_DECODE_RF_n6895, DLX_INST_DATA_PATH_DECODE_RF_n6894, 
      DLX_INST_DATA_PATH_DECODE_RF_n6893, DLX_INST_DATA_PATH_DECODE_RF_n6892, 
      DLX_INST_DATA_PATH_DECODE_RF_n6891, DLX_INST_DATA_PATH_DECODE_RF_n6890, 
      DLX_INST_DATA_PATH_DECODE_RF_n6889, DLX_INST_DATA_PATH_DECODE_RF_n6888, 
      DLX_INST_DATA_PATH_DECODE_RF_n6887, DLX_INST_DATA_PATH_DECODE_RF_n6886, 
      DLX_INST_DATA_PATH_DECODE_RF_n6885, DLX_INST_DATA_PATH_DECODE_RF_n6884, 
      DLX_INST_DATA_PATH_DECODE_RF_n6883, DLX_INST_DATA_PATH_DECODE_RF_n6882, 
      DLX_INST_DATA_PATH_DECODE_RF_n6881, DLX_INST_DATA_PATH_DECODE_RF_n6880, 
      DLX_INST_DATA_PATH_DECODE_RF_n6879, DLX_INST_DATA_PATH_DECODE_RF_n6878, 
      DLX_INST_DATA_PATH_DECODE_RF_n6877, DLX_INST_DATA_PATH_DECODE_RF_n6876, 
      DLX_INST_DATA_PATH_DECODE_RF_n6875, DLX_INST_DATA_PATH_DECODE_RF_n6874, 
      DLX_INST_DATA_PATH_DECODE_RF_n6873, DLX_INST_DATA_PATH_DECODE_RF_n6872, 
      DLX_INST_DATA_PATH_DECODE_RF_n6871, DLX_INST_DATA_PATH_DECODE_RF_n6870, 
      DLX_INST_DATA_PATH_DECODE_RF_n6869, DLX_INST_DATA_PATH_DECODE_RF_n6868, 
      DLX_INST_DATA_PATH_DECODE_RF_n6867, DLX_INST_DATA_PATH_DECODE_RF_n6866, 
      DLX_INST_DATA_PATH_DECODE_RF_n6865, DLX_INST_DATA_PATH_DECODE_RF_n6864, 
      DLX_INST_DATA_PATH_DECODE_RF_n6863, DLX_INST_DATA_PATH_DECODE_RF_n6862, 
      DLX_INST_DATA_PATH_DECODE_RF_n6861, DLX_INST_DATA_PATH_DECODE_RF_n6860, 
      DLX_INST_DATA_PATH_DECODE_RF_n6859, DLX_INST_DATA_PATH_DECODE_RF_n6858, 
      DLX_INST_DATA_PATH_DECODE_RF_n6857, DLX_INST_DATA_PATH_DECODE_RF_n6856, 
      DLX_INST_DATA_PATH_DECODE_RF_n6855, DLX_INST_DATA_PATH_DECODE_RF_n6854, 
      DLX_INST_DATA_PATH_DECODE_RF_n6853, DLX_INST_DATA_PATH_DECODE_RF_n6852, 
      DLX_INST_DATA_PATH_DECODE_RF_n6851, DLX_INST_DATA_PATH_DECODE_RF_n6850, 
      DLX_INST_DATA_PATH_DECODE_RF_n6849, DLX_INST_DATA_PATH_DECODE_RF_n6848, 
      DLX_INST_DATA_PATH_DECODE_RF_n6847, DLX_INST_DATA_PATH_DECODE_RF_n6846, 
      DLX_INST_DATA_PATH_DECODE_RF_n6845, DLX_INST_DATA_PATH_DECODE_RF_n6844, 
      DLX_INST_DATA_PATH_DECODE_RF_n6843, DLX_INST_DATA_PATH_DECODE_RF_n6842, 
      DLX_INST_DATA_PATH_DECODE_RF_n6841, DLX_INST_DATA_PATH_DECODE_RF_n6840, 
      DLX_INST_DATA_PATH_DECODE_RF_n6839, DLX_INST_DATA_PATH_DECODE_RF_n6838, 
      DLX_INST_DATA_PATH_DECODE_RF_n6837, DLX_INST_DATA_PATH_DECODE_RF_n6836, 
      DLX_INST_DATA_PATH_DECODE_RF_n6835, DLX_INST_DATA_PATH_DECODE_RF_n6834, 
      DLX_INST_DATA_PATH_DECODE_RF_n6833, DLX_INST_DATA_PATH_DECODE_RF_n6832, 
      DLX_INST_DATA_PATH_DECODE_RF_n6831, DLX_INST_DATA_PATH_DECODE_RF_n6830, 
      DLX_INST_DATA_PATH_DECODE_RF_n6829, DLX_INST_DATA_PATH_DECODE_RF_n6828, 
      DLX_INST_DATA_PATH_DECODE_RF_n6827, DLX_INST_DATA_PATH_DECODE_RF_n6826, 
      DLX_INST_DATA_PATH_DECODE_RF_n6825, DLX_INST_DATA_PATH_DECODE_RF_n6824, 
      DLX_INST_DATA_PATH_DECODE_RF_n6823, DLX_INST_DATA_PATH_DECODE_RF_n6822, 
      DLX_INST_DATA_PATH_DECODE_RF_n6821, DLX_INST_DATA_PATH_DECODE_RF_n6820, 
      DLX_INST_DATA_PATH_DECODE_RF_n6819, DLX_INST_DATA_PATH_DECODE_RF_n6818, 
      DLX_INST_DATA_PATH_DECODE_RF_n6817, DLX_INST_DATA_PATH_DECODE_RF_n6816, 
      DLX_INST_DATA_PATH_DECODE_RF_n6815, DLX_INST_DATA_PATH_DECODE_RF_n6814, 
      DLX_INST_DATA_PATH_DECODE_RF_n6813, DLX_INST_DATA_PATH_DECODE_RF_n6812, 
      DLX_INST_DATA_PATH_DECODE_RF_n6811, DLX_INST_DATA_PATH_DECODE_RF_n6810, 
      DLX_INST_DATA_PATH_DECODE_RF_n6809, DLX_INST_DATA_PATH_DECODE_RF_n6808, 
      DLX_INST_DATA_PATH_DECODE_RF_n6807, DLX_INST_DATA_PATH_DECODE_RF_n6806, 
      DLX_INST_DATA_PATH_DECODE_RF_n6805, DLX_INST_DATA_PATH_DECODE_RF_n6804, 
      DLX_INST_DATA_PATH_DECODE_RF_n6803, DLX_INST_DATA_PATH_DECODE_RF_n6802, 
      DLX_INST_DATA_PATH_DECODE_RF_n6801, DLX_INST_DATA_PATH_DECODE_RF_n6800, 
      DLX_INST_DATA_PATH_DECODE_RF_n6799, DLX_INST_DATA_PATH_DECODE_RF_n6798, 
      DLX_INST_DATA_PATH_DECODE_RF_n6797, DLX_INST_DATA_PATH_DECODE_RF_n6796, 
      DLX_INST_DATA_PATH_DECODE_RF_n6795, DLX_INST_DATA_PATH_DECODE_RF_n6794, 
      DLX_INST_DATA_PATH_DECODE_RF_n6793, DLX_INST_DATA_PATH_DECODE_RF_n6792, 
      DLX_INST_DATA_PATH_DECODE_RF_n6791, DLX_INST_DATA_PATH_DECODE_RF_n6790, 
      DLX_INST_DATA_PATH_DECODE_RF_n6789, DLX_INST_DATA_PATH_DECODE_RF_n6788, 
      DLX_INST_DATA_PATH_DECODE_RF_n6787, DLX_INST_DATA_PATH_DECODE_RF_n6786, 
      DLX_INST_DATA_PATH_DECODE_RF_n6785, DLX_INST_DATA_PATH_DECODE_RF_n6784, 
      DLX_INST_DATA_PATH_DECODE_RF_n6783, DLX_INST_DATA_PATH_DECODE_RF_n6782, 
      DLX_INST_DATA_PATH_DECODE_RF_n6781, DLX_INST_DATA_PATH_DECODE_RF_n6780, 
      DLX_INST_DATA_PATH_DECODE_RF_n6779, DLX_INST_DATA_PATH_DECODE_RF_n6778, 
      DLX_INST_DATA_PATH_DECODE_RF_n6777, DLX_INST_DATA_PATH_DECODE_RF_n6776, 
      DLX_INST_DATA_PATH_DECODE_RF_n6775, DLX_INST_DATA_PATH_DECODE_RF_n6774, 
      DLX_INST_DATA_PATH_DECODE_RF_n6773, DLX_INST_DATA_PATH_DECODE_RF_n6772, 
      DLX_INST_DATA_PATH_DECODE_RF_n6771, DLX_INST_DATA_PATH_DECODE_RF_n6770, 
      DLX_INST_DATA_PATH_DECODE_RF_n6769, DLX_INST_DATA_PATH_DECODE_RF_n6768, 
      DLX_INST_DATA_PATH_DECODE_RF_n6767, DLX_INST_DATA_PATH_DECODE_RF_n6766, 
      DLX_INST_DATA_PATH_DECODE_RF_n6765, DLX_INST_DATA_PATH_DECODE_RF_n6764, 
      DLX_INST_DATA_PATH_DECODE_RF_n6763, DLX_INST_DATA_PATH_DECODE_RF_n6762, 
      DLX_INST_DATA_PATH_DECODE_RF_n6761, DLX_INST_DATA_PATH_DECODE_RF_n6760, 
      DLX_INST_DATA_PATH_DECODE_RF_n6759, DLX_INST_DATA_PATH_DECODE_RF_n6758, 
      DLX_INST_DATA_PATH_DECODE_RF_n6757, DLX_INST_DATA_PATH_DECODE_RF_n6756, 
      DLX_INST_DATA_PATH_DECODE_RF_n6755, DLX_INST_DATA_PATH_DECODE_RF_n6754, 
      DLX_INST_DATA_PATH_DECODE_RF_n6753, DLX_INST_DATA_PATH_DECODE_RF_n6752, 
      DLX_INST_DATA_PATH_DECODE_RF_n6751, DLX_INST_DATA_PATH_DECODE_RF_n6750, 
      DLX_INST_DATA_PATH_DECODE_RF_n6749, DLX_INST_DATA_PATH_DECODE_RF_n6748, 
      DLX_INST_DATA_PATH_DECODE_RF_n6747, DLX_INST_DATA_PATH_DECODE_RF_n6746, 
      DLX_INST_DATA_PATH_DECODE_RF_n6745, DLX_INST_DATA_PATH_DECODE_RF_n6744, 
      DLX_INST_DATA_PATH_DECODE_RF_n6743, DLX_INST_DATA_PATH_DECODE_RF_n6742, 
      DLX_INST_DATA_PATH_DECODE_RF_n6741, DLX_INST_DATA_PATH_DECODE_RF_n6740, 
      DLX_INST_DATA_PATH_DECODE_RF_n6739, DLX_INST_DATA_PATH_DECODE_RF_n6738, 
      DLX_INST_DATA_PATH_DECODE_RF_n6737, DLX_INST_DATA_PATH_DECODE_RF_n6736, 
      DLX_INST_DATA_PATH_DECODE_RF_n6735, DLX_INST_DATA_PATH_DECODE_RF_n6734, 
      DLX_INST_DATA_PATH_DECODE_RF_n6733, DLX_INST_DATA_PATH_DECODE_RF_n6732, 
      DLX_INST_DATA_PATH_DECODE_RF_n6731, DLX_INST_DATA_PATH_DECODE_RF_n6730, 
      DLX_INST_DATA_PATH_DECODE_RF_n6729, DLX_INST_DATA_PATH_DECODE_RF_n6728, 
      DLX_INST_DATA_PATH_DECODE_RF_n6727, DLX_INST_DATA_PATH_DECODE_RF_n6726, 
      DLX_INST_DATA_PATH_DECODE_RF_n6725, DLX_INST_DATA_PATH_DECODE_RF_n6724, 
      DLX_INST_DATA_PATH_DECODE_RF_n6723, DLX_INST_DATA_PATH_DECODE_RF_n6722, 
      DLX_INST_DATA_PATH_DECODE_RF_n6721, DLX_INST_DATA_PATH_DECODE_RF_n6720, 
      DLX_INST_DATA_PATH_DECODE_RF_n6719, DLX_INST_DATA_PATH_DECODE_RF_n6718, 
      DLX_INST_DATA_PATH_DECODE_RF_n6717, DLX_INST_DATA_PATH_DECODE_RF_n6716, 
      DLX_INST_DATA_PATH_DECODE_RF_n6715, DLX_INST_DATA_PATH_DECODE_RF_n6714, 
      DLX_INST_DATA_PATH_DECODE_RF_n6713, DLX_INST_DATA_PATH_DECODE_RF_n6712, 
      DLX_INST_DATA_PATH_DECODE_RF_n6711, DLX_INST_DATA_PATH_DECODE_RF_n6710, 
      DLX_INST_DATA_PATH_DECODE_RF_n6709, DLX_INST_DATA_PATH_DECODE_RF_n6708, 
      DLX_INST_DATA_PATH_DECODE_RF_n6707, DLX_INST_DATA_PATH_DECODE_RF_n6706, 
      DLX_INST_DATA_PATH_DECODE_RF_n6705, DLX_INST_DATA_PATH_DECODE_RF_n6704, 
      DLX_INST_DATA_PATH_DECODE_RF_n6703, DLX_INST_DATA_PATH_DECODE_RF_n6702, 
      DLX_INST_DATA_PATH_DECODE_RF_n6701, DLX_INST_DATA_PATH_DECODE_RF_n6700, 
      DLX_INST_DATA_PATH_DECODE_RF_n6699, DLX_INST_DATA_PATH_DECODE_RF_n6698, 
      DLX_INST_DATA_PATH_DECODE_RF_n6697, DLX_INST_DATA_PATH_DECODE_RF_n6696, 
      DLX_INST_DATA_PATH_DECODE_RF_n6695, DLX_INST_DATA_PATH_DECODE_RF_n6694, 
      DLX_INST_DATA_PATH_DECODE_RF_n6693, DLX_INST_DATA_PATH_DECODE_RF_n6692, 
      DLX_INST_DATA_PATH_DECODE_RF_n6691, DLX_INST_DATA_PATH_DECODE_RF_n6690, 
      DLX_INST_DATA_PATH_DECODE_RF_n6689, DLX_INST_DATA_PATH_DECODE_RF_n6688, 
      DLX_INST_DATA_PATH_DECODE_RF_n6687, DLX_INST_DATA_PATH_DECODE_RF_n6686, 
      DLX_INST_DATA_PATH_DECODE_RF_n6685, DLX_INST_DATA_PATH_DECODE_RF_n6684, 
      DLX_INST_DATA_PATH_DECODE_RF_n6683, DLX_INST_DATA_PATH_DECODE_RF_n6682, 
      DLX_INST_DATA_PATH_DECODE_RF_n6681, DLX_INST_DATA_PATH_DECODE_RF_n6680, 
      DLX_INST_DATA_PATH_DECODE_RF_n6679, DLX_INST_DATA_PATH_DECODE_RF_n6678, 
      DLX_INST_DATA_PATH_DECODE_RF_n6677, DLX_INST_DATA_PATH_DECODE_RF_n6676, 
      DLX_INST_DATA_PATH_DECODE_RF_n6675, DLX_INST_DATA_PATH_DECODE_RF_n6674, 
      DLX_INST_DATA_PATH_DECODE_RF_n6673, DLX_INST_DATA_PATH_DECODE_RF_n6672, 
      DLX_INST_DATA_PATH_DECODE_RF_n6671, DLX_INST_DATA_PATH_DECODE_RF_n6670, 
      DLX_INST_DATA_PATH_DECODE_RF_n6669, DLX_INST_DATA_PATH_DECODE_RF_n6668, 
      DLX_INST_DATA_PATH_DECODE_RF_n6667, DLX_INST_DATA_PATH_DECODE_RF_n6666, 
      DLX_INST_DATA_PATH_DECODE_RF_n6665, DLX_INST_DATA_PATH_DECODE_RF_n6664, 
      DLX_INST_DATA_PATH_DECODE_RF_n6663, DLX_INST_DATA_PATH_DECODE_RF_n6662, 
      DLX_INST_DATA_PATH_DECODE_RF_n6661, DLX_INST_DATA_PATH_DECODE_RF_n6660, 
      DLX_INST_DATA_PATH_DECODE_RF_n6659, DLX_INST_DATA_PATH_DECODE_RF_n6658, 
      DLX_INST_DATA_PATH_DECODE_RF_n6657, DLX_INST_DATA_PATH_DECODE_RF_n6656, 
      DLX_INST_DATA_PATH_DECODE_RF_n6655, DLX_INST_DATA_PATH_DECODE_RF_n6654, 
      DLX_INST_DATA_PATH_DECODE_RF_n6653, DLX_INST_DATA_PATH_DECODE_RF_n6652, 
      DLX_INST_DATA_PATH_DECODE_RF_n6651, DLX_INST_DATA_PATH_DECODE_RF_n6650, 
      DLX_INST_DATA_PATH_DECODE_RF_n6649, DLX_INST_DATA_PATH_DECODE_RF_n6648, 
      DLX_INST_DATA_PATH_DECODE_RF_n6647, DLX_INST_DATA_PATH_DECODE_RF_n6646, 
      DLX_INST_DATA_PATH_DECODE_RF_n6645, DLX_INST_DATA_PATH_DECODE_RF_n6644, 
      DLX_INST_DATA_PATH_DECODE_RF_n6643, DLX_INST_DATA_PATH_DECODE_RF_n6642, 
      DLX_INST_DATA_PATH_DECODE_RF_n6641, DLX_INST_DATA_PATH_DECODE_RF_n6640, 
      DLX_INST_DATA_PATH_DECODE_RF_n6639, DLX_INST_DATA_PATH_DECODE_RF_n6638, 
      DLX_INST_DATA_PATH_DECODE_RF_n6637, DLX_INST_DATA_PATH_DECODE_RF_n6636, 
      DLX_INST_DATA_PATH_DECODE_RF_n6635, DLX_INST_DATA_PATH_DECODE_RF_n6634, 
      DLX_INST_DATA_PATH_DECODE_RF_n6633, DLX_INST_DATA_PATH_DECODE_RF_n6632, 
      DLX_INST_DATA_PATH_DECODE_RF_n6631, DLX_INST_DATA_PATH_DECODE_RF_n6630, 
      DLX_INST_DATA_PATH_DECODE_RF_n6629, DLX_INST_DATA_PATH_DECODE_RF_n6628, 
      DLX_INST_DATA_PATH_DECODE_RF_n6627, DLX_INST_DATA_PATH_DECODE_RF_n6626, 
      DLX_INST_DATA_PATH_DECODE_RF_n6625, DLX_INST_DATA_PATH_DECODE_RF_n6624, 
      DLX_INST_DATA_PATH_DECODE_RF_n6623, DLX_INST_DATA_PATH_DECODE_RF_n6622, 
      DLX_INST_DATA_PATH_DECODE_RF_n6621, DLX_INST_DATA_PATH_DECODE_RF_n6620, 
      DLX_INST_DATA_PATH_DECODE_RF_n6619, DLX_INST_DATA_PATH_DECODE_RF_n6618, 
      DLX_INST_DATA_PATH_DECODE_RF_n6617, DLX_INST_DATA_PATH_DECODE_RF_n6616, 
      DLX_INST_DATA_PATH_DECODE_RF_n6615, DLX_INST_DATA_PATH_DECODE_RF_n6614, 
      DLX_INST_DATA_PATH_DECODE_RF_n6613, DLX_INST_DATA_PATH_DECODE_RF_n6612, 
      DLX_INST_DATA_PATH_DECODE_RF_n6611, DLX_INST_DATA_PATH_DECODE_RF_n6610, 
      DLX_INST_DATA_PATH_DECODE_RF_n6609, DLX_INST_DATA_PATH_DECODE_RF_n6608, 
      DLX_INST_DATA_PATH_DECODE_RF_n6607, DLX_INST_DATA_PATH_DECODE_RF_n6606, 
      DLX_INST_DATA_PATH_DECODE_RF_n6605, DLX_INST_DATA_PATH_DECODE_RF_n6604, 
      DLX_INST_DATA_PATH_DECODE_RF_n6603, DLX_INST_DATA_PATH_DECODE_RF_n6602, 
      DLX_INST_DATA_PATH_DECODE_RF_n6601, DLX_INST_DATA_PATH_DECODE_RF_n6600, 
      DLX_INST_DATA_PATH_DECODE_RF_n6599, DLX_INST_DATA_PATH_DECODE_RF_n6598, 
      DLX_INST_DATA_PATH_DECODE_RF_n6597, DLX_INST_DATA_PATH_DECODE_RF_n6596, 
      DLX_INST_DATA_PATH_DECODE_RF_n6595, DLX_INST_DATA_PATH_DECODE_RF_n6594, 
      DLX_INST_DATA_PATH_DECODE_RF_n6593, DLX_INST_DATA_PATH_DECODE_RF_n6592, 
      DLX_INST_DATA_PATH_DECODE_RF_n6591, DLX_INST_DATA_PATH_DECODE_RF_n6590, 
      DLX_INST_DATA_PATH_DECODE_RF_n6589, DLX_INST_DATA_PATH_DECODE_RF_n6588, 
      DLX_INST_DATA_PATH_DECODE_RF_n6587, DLX_INST_DATA_PATH_DECODE_RF_n6586, 
      DLX_INST_DATA_PATH_DECODE_RF_n6585, DLX_INST_DATA_PATH_DECODE_RF_n6584, 
      DLX_INST_DATA_PATH_DECODE_RF_n6583, DLX_INST_DATA_PATH_DECODE_RF_n6582, 
      DLX_INST_DATA_PATH_DECODE_RF_n6581, DLX_INST_DATA_PATH_DECODE_RF_n6580, 
      DLX_INST_DATA_PATH_DECODE_RF_n6579, DLX_INST_DATA_PATH_DECODE_RF_n6578, 
      DLX_INST_DATA_PATH_DECODE_RF_n6577, DLX_INST_DATA_PATH_DECODE_RF_n6576, 
      DLX_INST_DATA_PATH_DECODE_RF_n6575, DLX_INST_DATA_PATH_DECODE_RF_n6574, 
      DLX_INST_DATA_PATH_DECODE_RF_n6573, DLX_INST_DATA_PATH_DECODE_RF_n6572, 
      DLX_INST_DATA_PATH_DECODE_RF_n6571, DLX_INST_DATA_PATH_DECODE_RF_n6570, 
      DLX_INST_DATA_PATH_DECODE_RF_n6569, DLX_INST_DATA_PATH_DECODE_RF_n6568, 
      DLX_INST_DATA_PATH_DECODE_RF_n6567, DLX_INST_DATA_PATH_DECODE_RF_n6566, 
      DLX_INST_DATA_PATH_DECODE_RF_n6565, DLX_INST_DATA_PATH_DECODE_RF_n6564, 
      DLX_INST_DATA_PATH_DECODE_RF_n6563, DLX_INST_DATA_PATH_DECODE_RF_n6562, 
      DLX_INST_DATA_PATH_DECODE_RF_n6561, DLX_INST_DATA_PATH_DECODE_RF_n6560, 
      DLX_INST_DATA_PATH_DECODE_RF_n6559, DLX_INST_DATA_PATH_DECODE_RF_n6558, 
      DLX_INST_DATA_PATH_DECODE_RF_n6557, DLX_INST_DATA_PATH_DECODE_RF_n6556, 
      DLX_INST_DATA_PATH_DECODE_RF_n6555, DLX_INST_DATA_PATH_DECODE_RF_n6554, 
      DLX_INST_DATA_PATH_DECODE_RF_n6553, DLX_INST_DATA_PATH_DECODE_RF_n6552, 
      DLX_INST_DATA_PATH_DECODE_RF_n6551, DLX_INST_DATA_PATH_DECODE_RF_n6550, 
      DLX_INST_DATA_PATH_DECODE_RF_n6549, DLX_INST_DATA_PATH_DECODE_RF_n6548, 
      DLX_INST_DATA_PATH_DECODE_RF_n6547, DLX_INST_DATA_PATH_DECODE_RF_n6546, 
      DLX_INST_DATA_PATH_DECODE_RF_n6545, DLX_INST_DATA_PATH_DECODE_RF_n6544, 
      DLX_INST_DATA_PATH_DECODE_RF_n6543, DLX_INST_DATA_PATH_DECODE_RF_n6542, 
      DLX_INST_DATA_PATH_DECODE_RF_n6541, DLX_INST_DATA_PATH_DECODE_RF_n6540, 
      DLX_INST_DATA_PATH_DECODE_RF_n6539, DLX_INST_DATA_PATH_DECODE_RF_n6538, 
      DLX_INST_DATA_PATH_DECODE_RF_n6537, DLX_INST_DATA_PATH_DECODE_RF_n6536, 
      DLX_INST_DATA_PATH_DECODE_RF_n6535, DLX_INST_DATA_PATH_DECODE_RF_n6534, 
      DLX_INST_DATA_PATH_DECODE_RF_n6533, DLX_INST_DATA_PATH_DECODE_RF_n6532, 
      DLX_INST_DATA_PATH_DECODE_RF_n6531, DLX_INST_DATA_PATH_DECODE_RF_n6530, 
      DLX_INST_DATA_PATH_DECODE_RF_n6529, DLX_INST_DATA_PATH_DECODE_RF_n6528, 
      DLX_INST_DATA_PATH_DECODE_RF_n6527, DLX_INST_DATA_PATH_DECODE_RF_n6526, 
      DLX_INST_DATA_PATH_DECODE_RF_n6525, DLX_INST_DATA_PATH_DECODE_RF_n6524, 
      DLX_INST_DATA_PATH_DECODE_RF_n6523, DLX_INST_DATA_PATH_DECODE_RF_n6522, 
      DLX_INST_DATA_PATH_DECODE_RF_n6521, DLX_INST_DATA_PATH_DECODE_RF_n6520, 
      DLX_INST_DATA_PATH_DECODE_RF_n6519, DLX_INST_DATA_PATH_DECODE_RF_n6518, 
      DLX_INST_DATA_PATH_DECODE_RF_n6517, DLX_INST_DATA_PATH_DECODE_RF_n6516, 
      DLX_INST_DATA_PATH_DECODE_RF_n6515, DLX_INST_DATA_PATH_DECODE_RF_n6514, 
      DLX_INST_DATA_PATH_DECODE_RF_n6513, DLX_INST_DATA_PATH_DECODE_RF_n6512, 
      DLX_INST_DATA_PATH_DECODE_RF_n6511, DLX_INST_DATA_PATH_DECODE_RF_n6510, 
      DLX_INST_DATA_PATH_DECODE_RF_n6509, DLX_INST_DATA_PATH_DECODE_RF_n6508, 
      DLX_INST_DATA_PATH_DECODE_RF_n6507, DLX_INST_DATA_PATH_DECODE_RF_n6506, 
      DLX_INST_DATA_PATH_DECODE_RF_n6505, DLX_INST_DATA_PATH_DECODE_RF_n6504, 
      DLX_INST_DATA_PATH_DECODE_RF_n6503, DLX_INST_DATA_PATH_DECODE_RF_n6502, 
      DLX_INST_DATA_PATH_DECODE_RF_n6501, DLX_INST_DATA_PATH_DECODE_RF_n6500, 
      DLX_INST_DATA_PATH_DECODE_RF_n6499, DLX_INST_DATA_PATH_DECODE_RF_n6498, 
      DLX_INST_DATA_PATH_DECODE_RF_n6497, DLX_INST_DATA_PATH_DECODE_RF_n6496, 
      DLX_INST_DATA_PATH_DECODE_RF_n6495, DLX_INST_DATA_PATH_DECODE_RF_n6494, 
      DLX_INST_DATA_PATH_DECODE_RF_n6493, DLX_INST_DATA_PATH_DECODE_RF_n6492, 
      DLX_INST_DATA_PATH_DECODE_RF_n6491, DLX_INST_DATA_PATH_DECODE_RF_n6490, 
      DLX_INST_DATA_PATH_DECODE_RF_n6489, DLX_INST_DATA_PATH_DECODE_RF_n6488, 
      DLX_INST_DATA_PATH_DECODE_RF_n6487, DLX_INST_DATA_PATH_DECODE_RF_n6486, 
      DLX_INST_DATA_PATH_DECODE_RF_n6485, DLX_INST_DATA_PATH_DECODE_RF_n6484, 
      DLX_INST_DATA_PATH_DECODE_RF_n6483, DLX_INST_DATA_PATH_DECODE_RF_n6482, 
      DLX_INST_DATA_PATH_DECODE_RF_n6481, DLX_INST_DATA_PATH_DECODE_RF_n6480, 
      DLX_INST_DATA_PATH_DECODE_RF_n6479, DLX_INST_DATA_PATH_DECODE_RF_n6478, 
      DLX_INST_DATA_PATH_DECODE_RF_n6477, DLX_INST_DATA_PATH_DECODE_RF_n6476, 
      DLX_INST_DATA_PATH_DECODE_RF_n6475, DLX_INST_DATA_PATH_DECODE_RF_n6474, 
      DLX_INST_DATA_PATH_DECODE_RF_n6473, DLX_INST_DATA_PATH_DECODE_RF_n6472, 
      DLX_INST_DATA_PATH_DECODE_RF_n6471, DLX_INST_DATA_PATH_DECODE_RF_n6470, 
      DLX_INST_DATA_PATH_DECODE_RF_n6469, DLX_INST_DATA_PATH_DECODE_RF_n6468, 
      DLX_INST_DATA_PATH_DECODE_RF_n6467, DLX_INST_DATA_PATH_DECODE_RF_n6466, 
      DLX_INST_DATA_PATH_DECODE_RF_n6465, DLX_INST_DATA_PATH_DECODE_RF_n6464, 
      DLX_INST_DATA_PATH_DECODE_RF_n6463, DLX_INST_DATA_PATH_DECODE_RF_n6462, 
      DLX_INST_DATA_PATH_DECODE_RF_n6461, DLX_INST_DATA_PATH_DECODE_RF_n6460, 
      DLX_INST_DATA_PATH_DECODE_RF_n6459, DLX_INST_DATA_PATH_DECODE_RF_n6458, 
      DLX_INST_DATA_PATH_DECODE_RF_n6457, DLX_INST_DATA_PATH_DECODE_RF_n6456, 
      DLX_INST_DATA_PATH_DECODE_RF_n6455, DLX_INST_DATA_PATH_DECODE_RF_n6454, 
      DLX_INST_DATA_PATH_DECODE_RF_n6453, DLX_INST_DATA_PATH_DECODE_RF_n6452, 
      DLX_INST_DATA_PATH_DECODE_RF_n6451, DLX_INST_DATA_PATH_DECODE_RF_n6450, 
      DLX_INST_DATA_PATH_DECODE_RF_n6449, DLX_INST_DATA_PATH_DECODE_RF_n6448, 
      DLX_INST_DATA_PATH_DECODE_RF_n6447, DLX_INST_DATA_PATH_DECODE_RF_n6446, 
      DLX_INST_DATA_PATH_DECODE_RF_n6445, DLX_INST_DATA_PATH_DECODE_RF_n6444, 
      DLX_INST_DATA_PATH_DECODE_RF_n6443, DLX_INST_DATA_PATH_DECODE_RF_n6442, 
      DLX_INST_DATA_PATH_DECODE_RF_n6441, DLX_INST_DATA_PATH_DECODE_RF_n6440, 
      DLX_INST_DATA_PATH_DECODE_RF_n6439, DLX_INST_DATA_PATH_DECODE_RF_n6438, 
      DLX_INST_DATA_PATH_DECODE_RF_n6437, DLX_INST_DATA_PATH_DECODE_RF_n6436, 
      DLX_INST_DATA_PATH_DECODE_RF_n6435, DLX_INST_DATA_PATH_DECODE_RF_n6434, 
      DLX_INST_DATA_PATH_DECODE_RF_n6433, DLX_INST_DATA_PATH_DECODE_RF_n6432, 
      DLX_INST_DATA_PATH_DECODE_RF_n6431, DLX_INST_DATA_PATH_DECODE_RF_n6430, 
      DLX_INST_DATA_PATH_DECODE_RF_n6429, DLX_INST_DATA_PATH_DECODE_RF_n6428, 
      DLX_INST_DATA_PATH_DECODE_RF_n6427, DLX_INST_DATA_PATH_DECODE_RF_n6426, 
      DLX_INST_DATA_PATH_DECODE_RF_n6425, DLX_INST_DATA_PATH_DECODE_RF_n6424, 
      DLX_INST_DATA_PATH_DECODE_RF_n6423, DLX_INST_DATA_PATH_DECODE_RF_n6422, 
      DLX_INST_DATA_PATH_DECODE_RF_n6421, DLX_INST_DATA_PATH_DECODE_RF_n6420, 
      DLX_INST_DATA_PATH_DECODE_RF_n6419, DLX_INST_DATA_PATH_DECODE_RF_n6418, 
      DLX_INST_DATA_PATH_DECODE_RF_n6417, DLX_INST_DATA_PATH_DECODE_RF_n6416, 
      DLX_INST_DATA_PATH_DECODE_RF_n6415, DLX_INST_DATA_PATH_DECODE_RF_n6414, 
      DLX_INST_DATA_PATH_DECODE_RF_n6413, DLX_INST_DATA_PATH_DECODE_RF_n6412, 
      DLX_INST_DATA_PATH_DECODE_RF_n6411, DLX_INST_DATA_PATH_DECODE_RF_n6410, 
      DLX_INST_DATA_PATH_DECODE_RF_n6409, DLX_INST_DATA_PATH_DECODE_RF_n6408, 
      DLX_INST_DATA_PATH_DECODE_RF_n6407, DLX_INST_DATA_PATH_DECODE_RF_n6406, 
      DLX_INST_DATA_PATH_DECODE_RF_n6405, DLX_INST_DATA_PATH_DECODE_RF_n6404, 
      DLX_INST_DATA_PATH_DECODE_RF_n6403, DLX_INST_DATA_PATH_DECODE_RF_n6402, 
      DLX_INST_DATA_PATH_DECODE_RF_n6401, DLX_INST_DATA_PATH_DECODE_RF_n6400, 
      DLX_INST_DATA_PATH_DECODE_RF_n6399, DLX_INST_DATA_PATH_DECODE_RF_n6398, 
      DLX_INST_DATA_PATH_DECODE_RF_n6397, DLX_INST_DATA_PATH_DECODE_RF_n6396, 
      DLX_INST_DATA_PATH_DECODE_RF_n6395, DLX_INST_DATA_PATH_DECODE_RF_n6394, 
      DLX_INST_DATA_PATH_DECODE_RF_n6393, DLX_INST_DATA_PATH_DECODE_RF_n6392, 
      DLX_INST_DATA_PATH_DECODE_RF_n6391, DLX_INST_DATA_PATH_DECODE_RF_n6390, 
      DLX_INST_DATA_PATH_DECODE_RF_n6389, DLX_INST_DATA_PATH_DECODE_RF_n6388, 
      DLX_INST_DATA_PATH_DECODE_RF_n6387, DLX_INST_DATA_PATH_DECODE_RF_n6386, 
      DLX_INST_DATA_PATH_DECODE_RF_n6385, DLX_INST_DATA_PATH_DECODE_RF_n6384, 
      DLX_INST_DATA_PATH_DECODE_RF_n6383, DLX_INST_DATA_PATH_DECODE_RF_n6382, 
      DLX_INST_DATA_PATH_DECODE_RF_n6381, DLX_INST_DATA_PATH_DECODE_RF_n6380, 
      DLX_INST_DATA_PATH_DECODE_RF_n6379, DLX_INST_DATA_PATH_DECODE_RF_n6378, 
      DLX_INST_DATA_PATH_DECODE_RF_n6377, DLX_INST_DATA_PATH_DECODE_RF_n6376, 
      DLX_INST_DATA_PATH_DECODE_RF_n6375, DLX_INST_DATA_PATH_DECODE_RF_n6374, 
      DLX_INST_DATA_PATH_DECODE_RF_n6373, DLX_INST_DATA_PATH_DECODE_RF_n6372, 
      DLX_INST_DATA_PATH_DECODE_RF_n6371, DLX_INST_DATA_PATH_DECODE_RF_n6370, 
      DLX_INST_DATA_PATH_DECODE_RF_n6369, DLX_INST_DATA_PATH_DECODE_RF_n6368, 
      DLX_INST_DATA_PATH_DECODE_RF_n6367, DLX_INST_DATA_PATH_DECODE_RF_n6366, 
      DLX_INST_DATA_PATH_DECODE_RF_n6365, DLX_INST_DATA_PATH_DECODE_RF_n6364, 
      DLX_INST_DATA_PATH_DECODE_RF_n6363, DLX_INST_DATA_PATH_DECODE_RF_n6362, 
      DLX_INST_DATA_PATH_DECODE_RF_n6361, DLX_INST_DATA_PATH_DECODE_RF_n6360, 
      DLX_INST_DATA_PATH_DECODE_RF_n6359, DLX_INST_DATA_PATH_DECODE_RF_n6358, 
      DLX_INST_DATA_PATH_DECODE_RF_n6357, DLX_INST_DATA_PATH_DECODE_RF_n6356, 
      DLX_INST_DATA_PATH_DECODE_RF_n6355, DLX_INST_DATA_PATH_DECODE_RF_n6354, 
      DLX_INST_DATA_PATH_DECODE_RF_n6353, DLX_INST_DATA_PATH_DECODE_RF_n6352, 
      DLX_INST_DATA_PATH_DECODE_RF_n6351, DLX_INST_DATA_PATH_DECODE_RF_n6350, 
      DLX_INST_DATA_PATH_DECODE_RF_n6349, DLX_INST_DATA_PATH_DECODE_RF_n6348, 
      DLX_INST_DATA_PATH_DECODE_RF_n6347, DLX_INST_DATA_PATH_DECODE_RF_n6346, 
      DLX_INST_DATA_PATH_DECODE_RF_n6345, DLX_INST_DATA_PATH_DECODE_RF_n6344, 
      DLX_INST_DATA_PATH_DECODE_RF_n6343, DLX_INST_DATA_PATH_DECODE_RF_n6342, 
      DLX_INST_DATA_PATH_DECODE_RF_n6341, DLX_INST_DATA_PATH_DECODE_RF_n6340, 
      DLX_INST_DATA_PATH_DECODE_RF_n6339, DLX_INST_DATA_PATH_DECODE_RF_n6338, 
      DLX_INST_DATA_PATH_DECODE_RF_n6337, DLX_INST_DATA_PATH_DECODE_RF_n6336, 
      DLX_INST_DATA_PATH_DECODE_RF_n6335, DLX_INST_DATA_PATH_DECODE_RF_n6334, 
      DLX_INST_DATA_PATH_DECODE_RF_n6333, DLX_INST_DATA_PATH_DECODE_RF_n6332, 
      DLX_INST_DATA_PATH_DECODE_RF_n6331, DLX_INST_DATA_PATH_DECODE_RF_n6330, 
      DLX_INST_DATA_PATH_DECODE_RF_n6329, DLX_INST_DATA_PATH_DECODE_RF_n6328, 
      DLX_INST_DATA_PATH_DECODE_RF_n6327, DLX_INST_DATA_PATH_DECODE_RF_n6326, 
      DLX_INST_DATA_PATH_DECODE_RF_n6325, DLX_INST_DATA_PATH_DECODE_RF_n6324, 
      DLX_INST_DATA_PATH_DECODE_RF_n6323, DLX_INST_DATA_PATH_DECODE_RF_n6322, 
      DLX_INST_DATA_PATH_DECODE_RF_n6321, DLX_INST_DATA_PATH_DECODE_RF_n6320, 
      DLX_INST_DATA_PATH_DECODE_RF_n6319, DLX_INST_DATA_PATH_DECODE_RF_n6318, 
      DLX_INST_DATA_PATH_DECODE_RF_n6317, DLX_INST_DATA_PATH_DECODE_RF_n6316, 
      DLX_INST_DATA_PATH_DECODE_RF_n6315, DLX_INST_DATA_PATH_DECODE_RF_n6314, 
      DLX_INST_DATA_PATH_DECODE_RF_n6313, DLX_INST_DATA_PATH_DECODE_RF_n6312, 
      DLX_INST_DATA_PATH_DECODE_RF_n6311, DLX_INST_DATA_PATH_DECODE_RF_n6310, 
      DLX_INST_DATA_PATH_DECODE_RF_n6309, DLX_INST_DATA_PATH_DECODE_RF_n6308, 
      DLX_INST_DATA_PATH_DECODE_RF_n6307, DLX_INST_DATA_PATH_DECODE_RF_n6306, 
      DLX_INST_DATA_PATH_DECODE_RF_n6305, DLX_INST_DATA_PATH_DECODE_RF_n6304, 
      DLX_INST_DATA_PATH_DECODE_RF_n6303, DLX_INST_DATA_PATH_DECODE_RF_n6302, 
      DLX_INST_DATA_PATH_DECODE_RF_n6301, DLX_INST_DATA_PATH_DECODE_RF_n6300, 
      DLX_INST_DATA_PATH_DECODE_RF_n6299, DLX_INST_DATA_PATH_DECODE_RF_n6298, 
      DLX_INST_DATA_PATH_DECODE_RF_n6297, DLX_INST_DATA_PATH_DECODE_RF_n6296, 
      DLX_INST_DATA_PATH_DECODE_RF_n6295, DLX_INST_DATA_PATH_DECODE_RF_n6294, 
      DLX_INST_DATA_PATH_DECODE_RF_n6293, DLX_INST_DATA_PATH_DECODE_RF_n6292, 
      DLX_INST_DATA_PATH_DECODE_RF_n6291, DLX_INST_DATA_PATH_DECODE_RF_n6290, 
      DLX_INST_DATA_PATH_DECODE_RF_n6289, DLX_INST_DATA_PATH_DECODE_RF_n6288, 
      DLX_INST_DATA_PATH_DECODE_RF_n6287, DLX_INST_DATA_PATH_DECODE_RF_n6286, 
      DLX_INST_DATA_PATH_DECODE_RF_n6285, DLX_INST_DATA_PATH_DECODE_RF_n6284, 
      DLX_INST_DATA_PATH_DECODE_RF_n6283, DLX_INST_DATA_PATH_DECODE_RF_n6282, 
      DLX_INST_DATA_PATH_DECODE_RF_n6281, DLX_INST_DATA_PATH_DECODE_RF_n6280, 
      DLX_INST_DATA_PATH_DECODE_RF_n6279, DLX_INST_DATA_PATH_DECODE_RF_n6278, 
      DLX_INST_DATA_PATH_DECODE_RF_n6277, DLX_INST_DATA_PATH_DECODE_RF_n6276, 
      DLX_INST_DATA_PATH_DECODE_RF_n6275, DLX_INST_DATA_PATH_DECODE_RF_n6274, 
      DLX_INST_DATA_PATH_DECODE_RF_n6273, DLX_INST_DATA_PATH_DECODE_RF_n6272, 
      DLX_INST_DATA_PATH_DECODE_RF_n6271, DLX_INST_DATA_PATH_DECODE_RF_n6270, 
      DLX_INST_DATA_PATH_DECODE_RF_n6269, DLX_INST_DATA_PATH_DECODE_RF_n6268, 
      DLX_INST_DATA_PATH_DECODE_RF_n6267, DLX_INST_DATA_PATH_DECODE_RF_n6266, 
      DLX_INST_DATA_PATH_DECODE_RF_n6265, DLX_INST_DATA_PATH_DECODE_RF_n6264, 
      DLX_INST_DATA_PATH_DECODE_RF_n6263, DLX_INST_DATA_PATH_DECODE_RF_n6262, 
      DLX_INST_DATA_PATH_DECODE_RF_n6261, DLX_INST_DATA_PATH_DECODE_RF_n6260, 
      DLX_INST_DATA_PATH_DECODE_RF_n6259, DLX_INST_DATA_PATH_DECODE_RF_n6258, 
      DLX_INST_DATA_PATH_DECODE_RF_n6257, DLX_INST_DATA_PATH_DECODE_RF_n6256, 
      DLX_INST_DATA_PATH_DECODE_RF_n6255, DLX_INST_DATA_PATH_DECODE_RF_n6254, 
      DLX_INST_DATA_PATH_DECODE_RF_n6253, DLX_INST_DATA_PATH_DECODE_RF_n6252, 
      DLX_INST_DATA_PATH_DECODE_RF_n6251, DLX_INST_DATA_PATH_DECODE_RF_n6250, 
      DLX_INST_DATA_PATH_DECODE_RF_n6249, DLX_INST_DATA_PATH_DECODE_RF_n6248, 
      DLX_INST_DATA_PATH_DECODE_RF_n6247, DLX_INST_DATA_PATH_DECODE_RF_n6246, 
      DLX_INST_DATA_PATH_DECODE_RF_n6245, DLX_INST_DATA_PATH_DECODE_RF_n6244, 
      DLX_INST_DATA_PATH_DECODE_RF_n6243, DLX_INST_DATA_PATH_DECODE_RF_n6242, 
      DLX_INST_DATA_PATH_DECODE_RF_n6241, DLX_INST_DATA_PATH_DECODE_RF_n6240, 
      DLX_INST_DATA_PATH_DECODE_RF_n6239, DLX_INST_DATA_PATH_DECODE_RF_n6238, 
      DLX_INST_DATA_PATH_DECODE_RF_n6237, DLX_INST_DATA_PATH_DECODE_RF_n6236, 
      DLX_INST_DATA_PATH_DECODE_RF_n6235, DLX_INST_DATA_PATH_DECODE_RF_n6234, 
      DLX_INST_DATA_PATH_DECODE_RF_n6233, DLX_INST_DATA_PATH_DECODE_RF_n6232, 
      DLX_INST_DATA_PATH_DECODE_RF_n6231, DLX_INST_DATA_PATH_DECODE_RF_n6230, 
      DLX_INST_DATA_PATH_DECODE_RF_n6229, DLX_INST_DATA_PATH_DECODE_RF_n6228, 
      DLX_INST_DATA_PATH_DECODE_RF_n6227, DLX_INST_DATA_PATH_DECODE_RF_n6226, 
      DLX_INST_DATA_PATH_DECODE_RF_n6225, DLX_INST_DATA_PATH_DECODE_RF_n6224, 
      DLX_INST_DATA_PATH_DECODE_RF_n6223, DLX_INST_DATA_PATH_DECODE_RF_n6222, 
      DLX_INST_DATA_PATH_DECODE_RF_n6221, DLX_INST_DATA_PATH_DECODE_RF_n6220, 
      DLX_INST_DATA_PATH_DECODE_RF_n6219, DLX_INST_DATA_PATH_DECODE_RF_n6218, 
      DLX_INST_DATA_PATH_DECODE_RF_n6217, DLX_INST_DATA_PATH_DECODE_RF_n6216, 
      DLX_INST_DATA_PATH_DECODE_RF_n6215, DLX_INST_DATA_PATH_DECODE_RF_n6214, 
      DLX_INST_DATA_PATH_DECODE_RF_n6213, DLX_INST_DATA_PATH_DECODE_RF_n6212, 
      DLX_INST_DATA_PATH_DECODE_RF_n6211, DLX_INST_DATA_PATH_DECODE_RF_n6210, 
      DLX_INST_DATA_PATH_DECODE_RF_n6209, DLX_INST_DATA_PATH_DECODE_RF_n6208, 
      DLX_INST_DATA_PATH_DECODE_RF_n6207, DLX_INST_DATA_PATH_DECODE_RF_n6206, 
      DLX_INST_DATA_PATH_DECODE_RF_n6205, DLX_INST_DATA_PATH_DECODE_RF_n6204, 
      DLX_INST_DATA_PATH_DECODE_RF_n6203, DLX_INST_DATA_PATH_DECODE_RF_n6202, 
      DLX_INST_DATA_PATH_DECODE_RF_n6201, DLX_INST_DATA_PATH_DECODE_RF_n6200, 
      DLX_INST_DATA_PATH_DECODE_RF_n6199, DLX_INST_DATA_PATH_DECODE_RF_n6198, 
      DLX_INST_DATA_PATH_DECODE_RF_n6197, DLX_INST_DATA_PATH_DECODE_RF_n6196, 
      DLX_INST_DATA_PATH_DECODE_RF_n6195, DLX_INST_DATA_PATH_DECODE_RF_n6194, 
      DLX_INST_DATA_PATH_DECODE_RF_n6193, DLX_INST_DATA_PATH_DECODE_RF_n6192, 
      DLX_INST_DATA_PATH_DECODE_RF_n6191, DLX_INST_DATA_PATH_DECODE_RF_n6190, 
      DLX_INST_DATA_PATH_DECODE_RF_n6189, DLX_INST_DATA_PATH_DECODE_RF_n6188, 
      DLX_INST_DATA_PATH_DECODE_RF_n6187, DLX_INST_DATA_PATH_DECODE_RF_n6186, 
      DLX_INST_DATA_PATH_DECODE_RF_n6185, DLX_INST_DATA_PATH_DECODE_RF_n6184, 
      DLX_INST_DATA_PATH_DECODE_RF_n6183, DLX_INST_DATA_PATH_DECODE_RF_n6182, 
      DLX_INST_DATA_PATH_DECODE_RF_n6181, DLX_INST_DATA_PATH_DECODE_RF_n6180, 
      DLX_INST_DATA_PATH_DECODE_RF_n6179, DLX_INST_DATA_PATH_DECODE_RF_n6178, 
      DLX_INST_DATA_PATH_DECODE_RF_n6177, DLX_INST_DATA_PATH_DECODE_RF_n6176, 
      DLX_INST_DATA_PATH_DECODE_RF_n6175, DLX_INST_DATA_PATH_DECODE_RF_n6174, 
      DLX_INST_DATA_PATH_DECODE_RF_n6173, DLX_INST_DATA_PATH_DECODE_RF_n6172, 
      DLX_INST_DATA_PATH_DECODE_RF_n6171, DLX_INST_DATA_PATH_DECODE_RF_n6170, 
      DLX_INST_DATA_PATH_DECODE_RF_n6169, DLX_INST_DATA_PATH_DECODE_RF_n6168, 
      DLX_INST_DATA_PATH_DECODE_RF_n6167, DLX_INST_DATA_PATH_DECODE_RF_n6166, 
      DLX_INST_DATA_PATH_DECODE_RF_n6165, DLX_INST_DATA_PATH_DECODE_RF_n6164, 
      DLX_INST_DATA_PATH_DECODE_RF_n6163, DLX_INST_DATA_PATH_DECODE_RF_n6162, 
      DLX_INST_DATA_PATH_DECODE_RF_n6161, DLX_INST_DATA_PATH_DECODE_RF_n6160, 
      DLX_INST_DATA_PATH_DECODE_RF_n6159, DLX_INST_DATA_PATH_DECODE_RF_n6158, 
      DLX_INST_DATA_PATH_DECODE_RF_n6157, DLX_INST_DATA_PATH_DECODE_RF_n6156, 
      DLX_INST_DATA_PATH_DECODE_RF_n6155, DLX_INST_DATA_PATH_DECODE_RF_n6154, 
      DLX_INST_DATA_PATH_DECODE_RF_n6153, DLX_INST_DATA_PATH_DECODE_RF_n6152, 
      DLX_INST_DATA_PATH_DECODE_RF_n6151, DLX_INST_DATA_PATH_DECODE_RF_n6150, 
      DLX_INST_DATA_PATH_DECODE_RF_n6149, DLX_INST_DATA_PATH_DECODE_RF_n6148, 
      DLX_INST_DATA_PATH_DECODE_RF_n6147, DLX_INST_DATA_PATH_DECODE_RF_n6146, 
      DLX_INST_DATA_PATH_DECODE_RF_n6145, DLX_INST_DATA_PATH_DECODE_RF_n6144, 
      DLX_INST_DATA_PATH_DECODE_RF_n6143, DLX_INST_DATA_PATH_DECODE_RF_n6142, 
      DLX_INST_DATA_PATH_DECODE_RF_n6141, DLX_INST_DATA_PATH_DECODE_RF_n6140, 
      DLX_INST_DATA_PATH_DECODE_RF_n6139, DLX_INST_DATA_PATH_DECODE_RF_n6138, 
      DLX_INST_DATA_PATH_DECODE_RF_n6137, DLX_INST_DATA_PATH_DECODE_RF_n6136, 
      DLX_INST_DATA_PATH_DECODE_RF_n6135, DLX_INST_DATA_PATH_DECODE_RF_n6134, 
      DLX_INST_DATA_PATH_DECODE_RF_n6133, DLX_INST_DATA_PATH_DECODE_RF_n6132, 
      DLX_INST_DATA_PATH_DECODE_RF_n6131, DLX_INST_DATA_PATH_DECODE_RF_n6130, 
      DLX_INST_DATA_PATH_DECODE_RF_n6129, DLX_INST_DATA_PATH_DECODE_RF_n6128, 
      DLX_INST_DATA_PATH_DECODE_RF_n6127, DLX_INST_DATA_PATH_DECODE_RF_n6126, 
      DLX_INST_DATA_PATH_DECODE_RF_n6125, DLX_INST_DATA_PATH_DECODE_RF_n6124, 
      DLX_INST_DATA_PATH_DECODE_RF_n6123, DLX_INST_DATA_PATH_DECODE_RF_n6122, 
      DLX_INST_DATA_PATH_DECODE_RF_n6121, DLX_INST_DATA_PATH_DECODE_RF_n6120, 
      DLX_INST_DATA_PATH_DECODE_RF_n6119, DLX_INST_DATA_PATH_DECODE_RF_n6118, 
      DLX_INST_DATA_PATH_DECODE_RF_n6117, DLX_INST_DATA_PATH_DECODE_RF_n6116, 
      DLX_INST_DATA_PATH_DECODE_RF_n6115, DLX_INST_DATA_PATH_DECODE_RF_n6114, 
      DLX_INST_DATA_PATH_DECODE_RF_n6113, DLX_INST_DATA_PATH_DECODE_RF_n6112, 
      DLX_INST_DATA_PATH_DECODE_RF_n6111, DLX_INST_DATA_PATH_DECODE_RF_n6110, 
      DLX_INST_DATA_PATH_DECODE_RF_n6109, DLX_INST_DATA_PATH_DECODE_RF_n6108, 
      DLX_INST_DATA_PATH_DECODE_RF_n6107, DLX_INST_DATA_PATH_DECODE_RF_n6106, 
      DLX_INST_DATA_PATH_DECODE_RF_n6105, DLX_INST_DATA_PATH_DECODE_RF_n6104, 
      DLX_INST_DATA_PATH_DECODE_RF_n6103, DLX_INST_DATA_PATH_DECODE_RF_n6102, 
      DLX_INST_DATA_PATH_DECODE_RF_n6101, DLX_INST_DATA_PATH_DECODE_RF_n6100, 
      DLX_INST_DATA_PATH_DECODE_RF_n6099, DLX_INST_DATA_PATH_DECODE_RF_n6098, 
      DLX_INST_DATA_PATH_DECODE_RF_n6097, DLX_INST_DATA_PATH_DECODE_RF_n6096, 
      DLX_INST_DATA_PATH_DECODE_RF_n6095, DLX_INST_DATA_PATH_DECODE_RF_n6094, 
      DLX_INST_DATA_PATH_DECODE_RF_n6093, DLX_INST_DATA_PATH_DECODE_RF_n6092, 
      DLX_INST_DATA_PATH_DECODE_RF_n6091, DLX_INST_DATA_PATH_DECODE_RF_n6090, 
      DLX_INST_DATA_PATH_DECODE_RF_n6089, DLX_INST_DATA_PATH_DECODE_RF_n6088, 
      DLX_INST_DATA_PATH_DECODE_RF_n6087, DLX_INST_DATA_PATH_DECODE_RF_n6086, 
      DLX_INST_DATA_PATH_DECODE_RF_n6085, DLX_INST_DATA_PATH_DECODE_RF_n6084, 
      DLX_INST_DATA_PATH_DECODE_RF_n6083, DLX_INST_DATA_PATH_DECODE_RF_n6082, 
      DLX_INST_DATA_PATH_DECODE_RF_n6081, DLX_INST_DATA_PATH_DECODE_RF_n6080, 
      DLX_INST_DATA_PATH_DECODE_RF_n6079, DLX_INST_DATA_PATH_DECODE_RF_n6078, 
      DLX_INST_DATA_PATH_DECODE_RF_n6077, DLX_INST_DATA_PATH_DECODE_RF_n6076, 
      DLX_INST_DATA_PATH_DECODE_RF_n6075, DLX_INST_DATA_PATH_DECODE_RF_n6074, 
      DLX_INST_DATA_PATH_DECODE_RF_n6073, DLX_INST_DATA_PATH_DECODE_RF_n6072, 
      DLX_INST_DATA_PATH_DECODE_RF_n6071, DLX_INST_DATA_PATH_DECODE_RF_n6070, 
      DLX_INST_DATA_PATH_DECODE_RF_n6069, DLX_INST_DATA_PATH_DECODE_RF_n6068, 
      DLX_INST_DATA_PATH_DECODE_RF_n6067, DLX_INST_DATA_PATH_DECODE_RF_n6066, 
      DLX_INST_DATA_PATH_DECODE_RF_n6065, DLX_INST_DATA_PATH_DECODE_RF_n6064, 
      DLX_INST_DATA_PATH_DECODE_RF_n6063, DLX_INST_DATA_PATH_DECODE_RF_n6062, 
      DLX_INST_DATA_PATH_DECODE_RF_n6061, DLX_INST_DATA_PATH_DECODE_RF_n6060, 
      DLX_INST_DATA_PATH_DECODE_RF_n6059, DLX_INST_DATA_PATH_DECODE_RF_n6058, 
      DLX_INST_DATA_PATH_DECODE_RF_n6057, DLX_INST_DATA_PATH_DECODE_RF_n6056, 
      DLX_INST_DATA_PATH_DECODE_RF_n6055, DLX_INST_DATA_PATH_DECODE_RF_n6054, 
      DLX_INST_DATA_PATH_DECODE_RF_n6053, DLX_INST_DATA_PATH_DECODE_RF_n6052, 
      DLX_INST_DATA_PATH_DECODE_RF_n6051, DLX_INST_DATA_PATH_DECODE_RF_n6050, 
      DLX_INST_DATA_PATH_DECODE_RF_n6049, DLX_INST_DATA_PATH_DECODE_RF_n6048, 
      DLX_INST_DATA_PATH_DECODE_RF_n6047, DLX_INST_DATA_PATH_DECODE_RF_n6046, 
      DLX_INST_DATA_PATH_DECODE_RF_n6045, DLX_INST_DATA_PATH_DECODE_RF_n6044, 
      DLX_INST_DATA_PATH_DECODE_RF_n6043, DLX_INST_DATA_PATH_DECODE_RF_n6042, 
      DLX_INST_DATA_PATH_DECODE_RF_n6041, DLX_INST_DATA_PATH_DECODE_RF_n6040, 
      DLX_INST_DATA_PATH_DECODE_RF_n6039, DLX_INST_DATA_PATH_DECODE_RF_n6038, 
      DLX_INST_DATA_PATH_DECODE_RF_n6037, DLX_INST_DATA_PATH_DECODE_RF_n6036, 
      DLX_INST_DATA_PATH_DECODE_RF_n6035, DLX_INST_DATA_PATH_DECODE_RF_n6034, 
      DLX_INST_DATA_PATH_DECODE_RF_n6033, DLX_INST_DATA_PATH_DECODE_RF_n6032, 
      DLX_INST_DATA_PATH_DECODE_RF_n6031, DLX_INST_DATA_PATH_DECODE_RF_n6030, 
      DLX_INST_DATA_PATH_DECODE_RF_n6029, DLX_INST_DATA_PATH_DECODE_RF_n6028, 
      DLX_INST_DATA_PATH_DECODE_RF_n6027, DLX_INST_DATA_PATH_DECODE_RF_n6026, 
      DLX_INST_DATA_PATH_DECODE_RF_n6025, DLX_INST_DATA_PATH_DECODE_RF_n6024, 
      DLX_INST_DATA_PATH_DECODE_RF_n6023, DLX_INST_DATA_PATH_DECODE_RF_n6022, 
      DLX_INST_DATA_PATH_DECODE_RF_n6021, DLX_INST_DATA_PATH_DECODE_RF_n6020, 
      DLX_INST_DATA_PATH_DECODE_RF_n6019, DLX_INST_DATA_PATH_DECODE_RF_n6018, 
      DLX_INST_DATA_PATH_DECODE_RF_n6017, DLX_INST_DATA_PATH_DECODE_RF_n6016, 
      DLX_INST_DATA_PATH_DECODE_RF_n6015, DLX_INST_DATA_PATH_DECODE_RF_n6014, 
      DLX_INST_DATA_PATH_DECODE_RF_n6013, DLX_INST_DATA_PATH_DECODE_RF_n6012, 
      DLX_INST_DATA_PATH_DECODE_RF_n6011, DLX_INST_DATA_PATH_DECODE_RF_n6010, 
      DLX_INST_DATA_PATH_DECODE_RF_n6009, DLX_INST_DATA_PATH_DECODE_RF_n6008, 
      DLX_INST_DATA_PATH_DECODE_RF_n6007, DLX_INST_DATA_PATH_DECODE_RF_n6006, 
      DLX_INST_DATA_PATH_DECODE_RF_n6005, DLX_INST_DATA_PATH_DECODE_RF_n6004, 
      DLX_INST_DATA_PATH_DECODE_RF_n6003, DLX_INST_DATA_PATH_DECODE_RF_n6002, 
      DLX_INST_DATA_PATH_DECODE_RF_n6001, DLX_INST_DATA_PATH_DECODE_RF_n6000, 
      DLX_INST_DATA_PATH_DECODE_RF_n5999, DLX_INST_DATA_PATH_DECODE_RF_n5998, 
      DLX_INST_DATA_PATH_DECODE_RF_n5997, DLX_INST_DATA_PATH_DECODE_RF_n5996, 
      DLX_INST_DATA_PATH_DECODE_RF_n5995, DLX_INST_DATA_PATH_DECODE_RF_n5994, 
      DLX_INST_DATA_PATH_DECODE_RF_n5993, DLX_INST_DATA_PATH_DECODE_RF_n5992, 
      DLX_INST_DATA_PATH_DECODE_RF_n5991, DLX_INST_DATA_PATH_DECODE_RF_n5990, 
      DLX_INST_DATA_PATH_DECODE_RF_n5989, DLX_INST_DATA_PATH_DECODE_RF_n5988, 
      DLX_INST_DATA_PATH_DECODE_RF_n5987, DLX_INST_DATA_PATH_DECODE_RF_n5986, 
      DLX_INST_DATA_PATH_DECODE_RF_n5985, DLX_INST_DATA_PATH_DECODE_RF_n5984, 
      DLX_INST_DATA_PATH_DECODE_RF_n5983, DLX_INST_DATA_PATH_DECODE_RF_n5982, 
      DLX_INST_DATA_PATH_DECODE_RF_n5981, DLX_INST_DATA_PATH_DECODE_RF_n5980, 
      DLX_INST_DATA_PATH_DECODE_RF_n5979, DLX_INST_DATA_PATH_DECODE_RF_n5978, 
      DLX_INST_DATA_PATH_DECODE_RF_n5977, DLX_INST_DATA_PATH_DECODE_RF_n5976, 
      DLX_INST_DATA_PATH_DECODE_RF_n5975, DLX_INST_DATA_PATH_DECODE_RF_n5974, 
      DLX_INST_DATA_PATH_DECODE_RF_n5973, DLX_INST_DATA_PATH_DECODE_RF_n5972, 
      DLX_INST_DATA_PATH_DECODE_RF_n5971, DLX_INST_DATA_PATH_DECODE_RF_n5970, 
      DLX_INST_DATA_PATH_DECODE_RF_n5969, DLX_INST_DATA_PATH_DECODE_RF_n5968, 
      DLX_INST_DATA_PATH_DECODE_RF_n5967, DLX_INST_DATA_PATH_DECODE_RF_n5966, 
      DLX_INST_DATA_PATH_DECODE_RF_n5965, DLX_INST_DATA_PATH_DECODE_RF_n5964, 
      DLX_INST_DATA_PATH_DECODE_RF_n5963, DLX_INST_DATA_PATH_DECODE_RF_n5962, 
      DLX_INST_DATA_PATH_DECODE_RF_n5961, DLX_INST_DATA_PATH_DECODE_RF_n5960, 
      DLX_INST_DATA_PATH_DECODE_RF_n5959, DLX_INST_DATA_PATH_DECODE_RF_n5958, 
      DLX_INST_DATA_PATH_DECODE_RF_n5957, DLX_INST_DATA_PATH_DECODE_RF_n5956, 
      DLX_INST_DATA_PATH_DECODE_RF_n5955, DLX_INST_DATA_PATH_DECODE_RF_n5954, 
      DLX_INST_DATA_PATH_DECODE_RF_n5953, DLX_INST_DATA_PATH_DECODE_RF_n5952, 
      DLX_INST_DATA_PATH_DECODE_RF_n5951, DLX_INST_DATA_PATH_DECODE_RF_n5950, 
      DLX_INST_DATA_PATH_DECODE_RF_n5949, DLX_INST_DATA_PATH_DECODE_RF_n5948, 
      DLX_INST_DATA_PATH_DECODE_RF_n5947, DLX_INST_DATA_PATH_DECODE_RF_n5946, 
      DLX_INST_DATA_PATH_DECODE_RF_n5945, DLX_INST_DATA_PATH_DECODE_RF_n5944, 
      DLX_INST_DATA_PATH_DECODE_RF_n5943, DLX_INST_DATA_PATH_DECODE_RF_n5942, 
      DLX_INST_DATA_PATH_DECODE_RF_n5941, DLX_INST_DATA_PATH_DECODE_RF_n5940, 
      DLX_INST_DATA_PATH_DECODE_RF_n5939, DLX_INST_DATA_PATH_DECODE_RF_n5938, 
      DLX_INST_DATA_PATH_DECODE_RF_n5937, DLX_INST_DATA_PATH_DECODE_RF_n5936, 
      DLX_INST_DATA_PATH_DECODE_RF_n5935, DLX_INST_DATA_PATH_DECODE_RF_n5934, 
      DLX_INST_DATA_PATH_DECODE_RF_n5933, DLX_INST_DATA_PATH_DECODE_RF_n5932, 
      DLX_INST_DATA_PATH_DECODE_RF_n5931, DLX_INST_DATA_PATH_DECODE_RF_n5930, 
      DLX_INST_DATA_PATH_DECODE_RF_n5929, DLX_INST_DATA_PATH_DECODE_RF_n5928, 
      DLX_INST_DATA_PATH_DECODE_RF_n5927, DLX_INST_DATA_PATH_DECODE_RF_n5926, 
      DLX_INST_DATA_PATH_DECODE_RF_n5925, DLX_INST_DATA_PATH_DECODE_RF_n5924, 
      DLX_INST_DATA_PATH_DECODE_RF_n5923, DLX_INST_DATA_PATH_DECODE_RF_n5922, 
      DLX_INST_DATA_PATH_DECODE_RF_n5921, DLX_INST_DATA_PATH_DECODE_RF_n5920, 
      DLX_INST_DATA_PATH_DECODE_RF_n5919, DLX_INST_DATA_PATH_DECODE_RF_n5918, 
      DLX_INST_DATA_PATH_DECODE_RF_n5917, DLX_INST_DATA_PATH_DECODE_RF_n5916, 
      DLX_INST_DATA_PATH_DECODE_RF_n5915, DLX_INST_DATA_PATH_DECODE_RF_n5914, 
      DLX_INST_DATA_PATH_DECODE_RF_n5913, DLX_INST_DATA_PATH_DECODE_RF_n5912, 
      DLX_INST_DATA_PATH_DECODE_RF_n5911, DLX_INST_DATA_PATH_DECODE_RF_n5910, 
      DLX_INST_DATA_PATH_DECODE_RF_n5909, DLX_INST_DATA_PATH_DECODE_RF_n5908, 
      DLX_INST_DATA_PATH_DECODE_RF_n5907, DLX_INST_DATA_PATH_DECODE_RF_n5906, 
      DLX_INST_DATA_PATH_DECODE_RF_n5905, DLX_INST_DATA_PATH_DECODE_RF_n5904, 
      DLX_INST_DATA_PATH_DECODE_RF_n5903, DLX_INST_DATA_PATH_DECODE_RF_n5902, 
      DLX_INST_DATA_PATH_DECODE_RF_n5901, DLX_INST_DATA_PATH_DECODE_RF_n5900, 
      DLX_INST_DATA_PATH_DECODE_RF_n5899, DLX_INST_DATA_PATH_DECODE_RF_n5898, 
      DLX_INST_DATA_PATH_DECODE_RF_n5897, DLX_INST_DATA_PATH_DECODE_RF_n5896, 
      DLX_INST_DATA_PATH_DECODE_RF_n5895, DLX_INST_DATA_PATH_DECODE_RF_n5894, 
      DLX_INST_DATA_PATH_DECODE_RF_n5893, DLX_INST_DATA_PATH_DECODE_RF_n5892, 
      DLX_INST_DATA_PATH_DECODE_RF_n5891, DLX_INST_DATA_PATH_DECODE_RF_n5890, 
      DLX_INST_DATA_PATH_DECODE_RF_n5889, DLX_INST_DATA_PATH_DECODE_RF_n5888, 
      DLX_INST_DATA_PATH_DECODE_RF_n5887, DLX_INST_DATA_PATH_DECODE_RF_n5886, 
      DLX_INST_DATA_PATH_DECODE_RF_n5885, DLX_INST_DATA_PATH_DECODE_RF_n5884, 
      DLX_INST_DATA_PATH_DECODE_RF_n5883, DLX_INST_DATA_PATH_DECODE_RF_n5882, 
      DLX_INST_DATA_PATH_DECODE_RF_n5881, DLX_INST_DATA_PATH_DECODE_RF_n5880, 
      DLX_INST_DATA_PATH_DECODE_RF_n5879, DLX_INST_DATA_PATH_DECODE_RF_n5878, 
      DLX_INST_DATA_PATH_DECODE_RF_n5877, DLX_INST_DATA_PATH_DECODE_RF_n5876, 
      DLX_INST_DATA_PATH_DECODE_RF_n5875, DLX_INST_DATA_PATH_DECODE_RF_n5874, 
      DLX_INST_DATA_PATH_DECODE_RF_n5873, DLX_INST_DATA_PATH_DECODE_RF_n5872, 
      DLX_INST_DATA_PATH_DECODE_RF_n5871, DLX_INST_DATA_PATH_DECODE_RF_n5870, 
      DLX_INST_DATA_PATH_DECODE_RF_n5869, DLX_INST_DATA_PATH_DECODE_RF_n5868, 
      DLX_INST_DATA_PATH_DECODE_RF_n5867, DLX_INST_DATA_PATH_DECODE_RF_n5866, 
      DLX_INST_DATA_PATH_DECODE_RF_n5865, DLX_INST_DATA_PATH_DECODE_RF_n5864, 
      DLX_INST_DATA_PATH_DECODE_RF_n5863, DLX_INST_DATA_PATH_DECODE_RF_n5862, 
      DLX_INST_DATA_PATH_DECODE_RF_n5861, DLX_INST_DATA_PATH_DECODE_RF_n5860, 
      DLX_INST_DATA_PATH_DECODE_RF_n5859, DLX_INST_DATA_PATH_DECODE_RF_n5858, 
      DLX_INST_DATA_PATH_DECODE_RF_n5857, DLX_INST_DATA_PATH_DECODE_RF_n5856, 
      DLX_INST_DATA_PATH_DECODE_RF_n5855, DLX_INST_DATA_PATH_DECODE_RF_n5854, 
      DLX_INST_DATA_PATH_DECODE_RF_n5853, DLX_INST_DATA_PATH_DECODE_RF_n5852, 
      DLX_INST_DATA_PATH_DECODE_RF_n5851, DLX_INST_DATA_PATH_DECODE_RF_n5850, 
      DLX_INST_DATA_PATH_DECODE_RF_n5849, DLX_INST_DATA_PATH_DECODE_RF_n5848, 
      DLX_INST_DATA_PATH_DECODE_RF_n5847, DLX_INST_DATA_PATH_DECODE_RF_n5846, 
      DLX_INST_DATA_PATH_DECODE_RF_n5845, DLX_INST_DATA_PATH_DECODE_RF_n5844, 
      DLX_INST_DATA_PATH_DECODE_RF_n5843, DLX_INST_DATA_PATH_DECODE_RF_n5842, 
      DLX_INST_DATA_PATH_DECODE_RF_n5841, DLX_INST_DATA_PATH_DECODE_RF_n5840, 
      DLX_INST_DATA_PATH_DECODE_RF_n5839, DLX_INST_DATA_PATH_DECODE_RF_n5838, 
      DLX_INST_DATA_PATH_DECODE_RF_n5837, DLX_INST_DATA_PATH_DECODE_RF_n5836, 
      DLX_INST_DATA_PATH_DECODE_RF_n5835, DLX_INST_DATA_PATH_DECODE_RF_n5834, 
      DLX_INST_DATA_PATH_DECODE_RF_n5833, DLX_INST_DATA_PATH_DECODE_RF_n5832, 
      DLX_INST_DATA_PATH_DECODE_RF_n5831, DLX_INST_DATA_PATH_DECODE_RF_n5830, 
      DLX_INST_DATA_PATH_DECODE_RF_n5829, DLX_INST_DATA_PATH_DECODE_RF_n5828, 
      DLX_INST_DATA_PATH_DECODE_RF_n5827, DLX_INST_DATA_PATH_DECODE_RF_n5826, 
      DLX_INST_DATA_PATH_DECODE_RF_n5825, DLX_INST_DATA_PATH_DECODE_RF_n5824, 
      DLX_INST_DATA_PATH_DECODE_RF_n5823, DLX_INST_DATA_PATH_DECODE_RF_n5822, 
      DLX_INST_DATA_PATH_DECODE_RF_n5821, DLX_INST_DATA_PATH_DECODE_RF_n5820, 
      DLX_INST_DATA_PATH_DECODE_RF_n5819, DLX_INST_DATA_PATH_DECODE_RF_n5818, 
      DLX_INST_DATA_PATH_DECODE_RF_n5817, DLX_INST_DATA_PATH_DECODE_RF_n5816, 
      DLX_INST_DATA_PATH_DECODE_RF_n5815, DLX_INST_DATA_PATH_DECODE_RF_n5814, 
      DLX_INST_DATA_PATH_DECODE_RF_n5813, DLX_INST_DATA_PATH_DECODE_RF_n5812, 
      DLX_INST_DATA_PATH_DECODE_RF_n5811, DLX_INST_DATA_PATH_DECODE_RF_n5810, 
      DLX_INST_DATA_PATH_DECODE_RF_n5809, DLX_INST_DATA_PATH_DECODE_RF_n5808, 
      DLX_INST_DATA_PATH_DECODE_RF_n5807, DLX_INST_DATA_PATH_DECODE_RF_n5806, 
      DLX_INST_DATA_PATH_DECODE_RF_n5805, DLX_INST_DATA_PATH_DECODE_RF_n5804, 
      DLX_INST_DATA_PATH_DECODE_RF_n5803, DLX_INST_DATA_PATH_DECODE_RF_n5802, 
      DLX_INST_DATA_PATH_DECODE_RF_n5801, DLX_INST_DATA_PATH_DECODE_RF_n5800, 
      DLX_INST_DATA_PATH_DECODE_RF_n5799, DLX_INST_DATA_PATH_DECODE_RF_n5798, 
      DLX_INST_DATA_PATH_DECODE_RF_n5797, DLX_INST_DATA_PATH_DECODE_RF_n5796, 
      DLX_INST_DATA_PATH_DECODE_RF_n5795, DLX_INST_DATA_PATH_DECODE_RF_n5794, 
      DLX_INST_DATA_PATH_DECODE_RF_n5793, DLX_INST_DATA_PATH_DECODE_RF_n5792, 
      DLX_INST_DATA_PATH_DECODE_RF_n5791, DLX_INST_DATA_PATH_DECODE_RF_n5790, 
      DLX_INST_DATA_PATH_DECODE_RF_n5789, DLX_INST_DATA_PATH_DECODE_RF_n5788, 
      DLX_INST_DATA_PATH_DECODE_RF_n5787, DLX_INST_DATA_PATH_DECODE_RF_n5786, 
      DLX_INST_DATA_PATH_DECODE_RF_n5785, DLX_INST_DATA_PATH_DECODE_RF_n5784, 
      DLX_INST_DATA_PATH_DECODE_RF_n5783, DLX_INST_DATA_PATH_DECODE_RF_n5782, 
      DLX_INST_DATA_PATH_DECODE_RF_n5781, DLX_INST_DATA_PATH_DECODE_RF_n5780, 
      DLX_INST_DATA_PATH_DECODE_RF_n5779, DLX_INST_DATA_PATH_DECODE_RF_n5778, 
      DLX_INST_DATA_PATH_DECODE_RF_n5777, DLX_INST_DATA_PATH_DECODE_RF_n5776, 
      DLX_INST_DATA_PATH_DECODE_RF_n5775, DLX_INST_DATA_PATH_DECODE_RF_n5774, 
      DLX_INST_DATA_PATH_DECODE_RF_n5773, DLX_INST_DATA_PATH_DECODE_RF_n5772, 
      DLX_INST_DATA_PATH_DECODE_RF_n5771, DLX_INST_DATA_PATH_DECODE_RF_n5770, 
      DLX_INST_DATA_PATH_DECODE_RF_n5769, DLX_INST_DATA_PATH_DECODE_RF_n5768, 
      DLX_INST_DATA_PATH_DECODE_RF_n5767, DLX_INST_DATA_PATH_DECODE_RF_n5766, 
      DLX_INST_DATA_PATH_DECODE_RF_n5765, DLX_INST_DATA_PATH_DECODE_RF_n5764, 
      DLX_INST_DATA_PATH_DECODE_RF_n5763, DLX_INST_DATA_PATH_DECODE_RF_n5762, 
      DLX_INST_DATA_PATH_DECODE_RF_n5761, DLX_INST_DATA_PATH_DECODE_RF_n5760, 
      DLX_INST_DATA_PATH_DECODE_RF_n5759, DLX_INST_DATA_PATH_DECODE_RF_n5758, 
      DLX_INST_DATA_PATH_DECODE_RF_n5757, DLX_INST_DATA_PATH_DECODE_RF_n5756, 
      DLX_INST_DATA_PATH_DECODE_RF_n5755, DLX_INST_DATA_PATH_DECODE_RF_n5754, 
      DLX_INST_DATA_PATH_DECODE_RF_n5753, DLX_INST_DATA_PATH_DECODE_RF_n5752, 
      DLX_INST_DATA_PATH_DECODE_RF_n5751, DLX_INST_DATA_PATH_DECODE_RF_n5750, 
      DLX_INST_DATA_PATH_DECODE_RF_n5749, DLX_INST_DATA_PATH_DECODE_RF_n5748, 
      DLX_INST_DATA_PATH_DECODE_RF_n5747, DLX_INST_DATA_PATH_DECODE_RF_n5746, 
      DLX_INST_DATA_PATH_DECODE_RF_n5745, DLX_INST_DATA_PATH_DECODE_RF_n5744, 
      DLX_INST_DATA_PATH_DECODE_RF_n5743, DLX_INST_DATA_PATH_DECODE_RF_n5742, 
      DLX_INST_DATA_PATH_DECODE_RF_n5741, DLX_INST_DATA_PATH_DECODE_RF_n5740, 
      DLX_INST_DATA_PATH_DECODE_RF_n5739, DLX_INST_DATA_PATH_DECODE_RF_n5738, 
      DLX_INST_DATA_PATH_DECODE_RF_n5737, DLX_INST_DATA_PATH_DECODE_RF_n5736, 
      DLX_INST_DATA_PATH_DECODE_RF_n5735, DLX_INST_DATA_PATH_DECODE_RF_n5734, 
      DLX_INST_DATA_PATH_DECODE_RF_n5733, DLX_INST_DATA_PATH_DECODE_RF_n5732, 
      DLX_INST_DATA_PATH_DECODE_RF_n5731, DLX_INST_DATA_PATH_DECODE_RF_n5730, 
      DLX_INST_DATA_PATH_DECODE_RF_n5729, DLX_INST_DATA_PATH_DECODE_RF_n5728, 
      DLX_INST_DATA_PATH_DECODE_RF_n5727, DLX_INST_DATA_PATH_DECODE_RF_n5726, 
      DLX_INST_DATA_PATH_DECODE_RF_n5725, DLX_INST_DATA_PATH_DECODE_RF_n5724, 
      DLX_INST_DATA_PATH_DECODE_RF_n5723, DLX_INST_DATA_PATH_DECODE_RF_n5722, 
      DLX_INST_DATA_PATH_DECODE_RF_n5721, DLX_INST_DATA_PATH_DECODE_RF_n5720, 
      DLX_INST_DATA_PATH_DECODE_RF_n5719, DLX_INST_DATA_PATH_DECODE_RF_n5718, 
      DLX_INST_DATA_PATH_DECODE_RF_n5717, DLX_INST_DATA_PATH_DECODE_RF_n5716, 
      DLX_INST_DATA_PATH_DECODE_RF_n5715, DLX_INST_DATA_PATH_DECODE_RF_n5714, 
      DLX_INST_DATA_PATH_DECODE_RF_n5713, DLX_INST_DATA_PATH_DECODE_RF_n5712, 
      DLX_INST_DATA_PATH_DECODE_RF_n5711, DLX_INST_DATA_PATH_DECODE_RF_n5710, 
      DLX_INST_DATA_PATH_DECODE_RF_n5709, DLX_INST_DATA_PATH_DECODE_RF_n5708, 
      DLX_INST_DATA_PATH_DECODE_RF_n5707, DLX_INST_DATA_PATH_DECODE_RF_n5706, 
      DLX_INST_DATA_PATH_DECODE_RF_n5705, DLX_INST_DATA_PATH_DECODE_RF_n5704, 
      DLX_INST_DATA_PATH_DECODE_RF_n5703, DLX_INST_DATA_PATH_DECODE_RF_n5702, 
      DLX_INST_DATA_PATH_DECODE_RF_n5701, DLX_INST_DATA_PATH_DECODE_RF_n5700, 
      DLX_INST_DATA_PATH_DECODE_RF_n5699, DLX_INST_DATA_PATH_DECODE_RF_n5698, 
      DLX_INST_DATA_PATH_DECODE_RF_n5697, DLX_INST_DATA_PATH_DECODE_RF_n5696, 
      DLX_INST_DATA_PATH_DECODE_RF_n5695, DLX_INST_DATA_PATH_DECODE_RF_n5694, 
      DLX_INST_DATA_PATH_DECODE_RF_n5693, DLX_INST_DATA_PATH_DECODE_RF_n5692, 
      DLX_INST_DATA_PATH_DECODE_RF_n5691, DLX_INST_DATA_PATH_DECODE_RF_n5690, 
      DLX_INST_DATA_PATH_DECODE_RF_n5689, DLX_INST_DATA_PATH_DECODE_RF_n5688, 
      DLX_INST_DATA_PATH_DECODE_RF_n5687, DLX_INST_DATA_PATH_DECODE_RF_n5686, 
      DLX_INST_DATA_PATH_DECODE_RF_n5685, DLX_INST_DATA_PATH_DECODE_RF_n5684, 
      DLX_INST_DATA_PATH_DECODE_RF_n5683, DLX_INST_DATA_PATH_DECODE_RF_n5682, 
      DLX_INST_DATA_PATH_DECODE_RF_n5681, DLX_INST_DATA_PATH_DECODE_RF_n5680, 
      DLX_INST_DATA_PATH_DECODE_RF_n5679, DLX_INST_DATA_PATH_DECODE_RF_n5678, 
      DLX_INST_DATA_PATH_DECODE_RF_n5677, DLX_INST_DATA_PATH_DECODE_RF_n5676, 
      DLX_INST_DATA_PATH_DECODE_RF_n5675, DLX_INST_DATA_PATH_DECODE_RF_n5674, 
      DLX_INST_DATA_PATH_DECODE_RF_n5673, DLX_INST_DATA_PATH_DECODE_RF_n5672, 
      DLX_INST_DATA_PATH_DECODE_RF_n5671, DLX_INST_DATA_PATH_DECODE_RF_n5670, 
      DLX_INST_DATA_PATH_DECODE_RF_n5669, DLX_INST_DATA_PATH_DECODE_RF_n5668, 
      DLX_INST_DATA_PATH_DECODE_RF_n5667, DLX_INST_DATA_PATH_DECODE_RF_n5666, 
      DLX_INST_DATA_PATH_DECODE_RF_n5665, DLX_INST_DATA_PATH_DECODE_RF_n5664, 
      DLX_INST_DATA_PATH_DECODE_RF_n5663, DLX_INST_DATA_PATH_DECODE_RF_n5662, 
      DLX_INST_DATA_PATH_DECODE_RF_n5661, DLX_INST_DATA_PATH_DECODE_RF_n5660, 
      DLX_INST_DATA_PATH_DECODE_RF_n5659, DLX_INST_DATA_PATH_DECODE_RF_n5658, 
      DLX_INST_DATA_PATH_DECODE_RF_n5657, DLX_INST_DATA_PATH_DECODE_RF_n5656, 
      DLX_INST_DATA_PATH_DECODE_RF_n5655, DLX_INST_DATA_PATH_DECODE_RF_n5654, 
      DLX_INST_DATA_PATH_DECODE_RF_n5653, DLX_INST_DATA_PATH_DECODE_RF_n5652, 
      DLX_INST_DATA_PATH_DECODE_RF_n5651, DLX_INST_DATA_PATH_DECODE_RF_n5650, 
      DLX_INST_DATA_PATH_DECODE_RF_n5649, DLX_INST_DATA_PATH_DECODE_RF_n5648, 
      DLX_INST_DATA_PATH_DECODE_RF_n5647, DLX_INST_DATA_PATH_DECODE_RF_n5646, 
      DLX_INST_DATA_PATH_DECODE_RF_n5645, DLX_INST_DATA_PATH_DECODE_RF_n5644, 
      DLX_INST_DATA_PATH_DECODE_RF_n5643, DLX_INST_DATA_PATH_DECODE_RF_n5642, 
      DLX_INST_DATA_PATH_DECODE_RF_n5641, DLX_INST_DATA_PATH_DECODE_RF_n5640, 
      DLX_INST_DATA_PATH_DECODE_RF_n5639, DLX_INST_DATA_PATH_DECODE_RF_n5638, 
      DLX_INST_DATA_PATH_DECODE_RF_n5637, DLX_INST_DATA_PATH_DECODE_RF_n5636, 
      DLX_INST_DATA_PATH_DECODE_RF_n5635, DLX_INST_DATA_PATH_DECODE_RF_n5634, 
      DLX_INST_DATA_PATH_DECODE_RF_n5633, DLX_INST_DATA_PATH_DECODE_RF_n5632, 
      DLX_INST_DATA_PATH_DECODE_RF_n5631, DLX_INST_DATA_PATH_DECODE_RF_n5630, 
      DLX_INST_DATA_PATH_DECODE_RF_n5629, DLX_INST_DATA_PATH_DECODE_RF_n5628, 
      DLX_INST_DATA_PATH_DECODE_RF_n5627, DLX_INST_DATA_PATH_DECODE_RF_n5626, 
      DLX_INST_DATA_PATH_DECODE_RF_n5625, DLX_INST_DATA_PATH_DECODE_RF_n5624, 
      DLX_INST_DATA_PATH_DECODE_RF_n5623, DLX_INST_DATA_PATH_DECODE_RF_n5622, 
      DLX_INST_DATA_PATH_DECODE_RF_n5621, DLX_INST_DATA_PATH_DECODE_RF_n5620, 
      DLX_INST_DATA_PATH_DECODE_RF_n5619, DLX_INST_DATA_PATH_DECODE_RF_n5618, 
      DLX_INST_DATA_PATH_DECODE_RF_n5617, DLX_INST_DATA_PATH_DECODE_RF_n5616, 
      DLX_INST_DATA_PATH_DECODE_RF_n5615, DLX_INST_DATA_PATH_DECODE_RF_n5614, 
      DLX_INST_DATA_PATH_DECODE_RF_n5613, DLX_INST_DATA_PATH_DECODE_RF_n5612, 
      DLX_INST_DATA_PATH_DECODE_RF_n5611, DLX_INST_DATA_PATH_DECODE_RF_n5610, 
      DLX_INST_DATA_PATH_DECODE_RF_n5609, DLX_INST_DATA_PATH_DECODE_RF_n5608, 
      DLX_INST_DATA_PATH_DECODE_RF_n5607, DLX_INST_DATA_PATH_DECODE_RF_n5606, 
      DLX_INST_DATA_PATH_DECODE_RF_n5605, DLX_INST_DATA_PATH_DECODE_RF_n5604, 
      DLX_INST_DATA_PATH_DECODE_RF_n5603, DLX_INST_DATA_PATH_DECODE_RF_n5602, 
      DLX_INST_DATA_PATH_DECODE_RF_n5601, DLX_INST_DATA_PATH_DECODE_RF_n5600, 
      DLX_INST_DATA_PATH_DECODE_RF_n5599, DLX_INST_DATA_PATH_DECODE_RF_n5598, 
      DLX_INST_DATA_PATH_DECODE_RF_n5597, DLX_INST_DATA_PATH_DECODE_RF_n5596, 
      DLX_INST_DATA_PATH_DECODE_RF_n5595, DLX_INST_DATA_PATH_DECODE_RF_n5594, 
      DLX_INST_DATA_PATH_DECODE_RF_n5593, DLX_INST_DATA_PATH_DECODE_RF_n5592, 
      DLX_INST_DATA_PATH_DECODE_RF_n5591, DLX_INST_DATA_PATH_DECODE_RF_n5590, 
      DLX_INST_DATA_PATH_DECODE_RF_n5589, DLX_INST_DATA_PATH_DECODE_RF_n5588, 
      DLX_INST_DATA_PATH_DECODE_RF_n5587, DLX_INST_DATA_PATH_DECODE_RF_n5586, 
      DLX_INST_DATA_PATH_DECODE_RF_n5585, DLX_INST_DATA_PATH_DECODE_RF_n5584, 
      DLX_INST_DATA_PATH_DECODE_RF_n5583, DLX_INST_DATA_PATH_DECODE_RF_n5582, 
      DLX_INST_DATA_PATH_DECODE_RF_n5581, DLX_INST_DATA_PATH_DECODE_RF_n5580, 
      DLX_INST_DATA_PATH_DECODE_RF_n5579, DLX_INST_DATA_PATH_DECODE_RF_n5578, 
      DLX_INST_DATA_PATH_DECODE_RF_n5577, DLX_INST_DATA_PATH_DECODE_RF_n5576, 
      DLX_INST_DATA_PATH_DECODE_RF_n5575, DLX_INST_DATA_PATH_DECODE_RF_n5574, 
      DLX_INST_DATA_PATH_DECODE_RF_n5573, DLX_INST_DATA_PATH_DECODE_RF_n5572, 
      DLX_INST_DATA_PATH_DECODE_RF_n5571, DLX_INST_DATA_PATH_DECODE_RF_n5570, 
      DLX_INST_DATA_PATH_DECODE_RF_n5569, DLX_INST_DATA_PATH_DECODE_RF_n5568, 
      DLX_INST_DATA_PATH_DECODE_RF_n5567, DLX_INST_DATA_PATH_DECODE_RF_n5566, 
      DLX_INST_DATA_PATH_DECODE_RF_n5565, DLX_INST_DATA_PATH_DECODE_RF_n5564, 
      DLX_INST_DATA_PATH_DECODE_RF_n5563, DLX_INST_DATA_PATH_DECODE_RF_n5562, 
      DLX_INST_DATA_PATH_DECODE_RF_n5561, DLX_INST_DATA_PATH_DECODE_RF_n5560, 
      DLX_INST_DATA_PATH_DECODE_RF_n5559, DLX_INST_DATA_PATH_DECODE_RF_n5558, 
      DLX_INST_DATA_PATH_DECODE_RF_n5557, DLX_INST_DATA_PATH_DECODE_RF_n5556, 
      DLX_INST_DATA_PATH_DECODE_RF_n5555, DLX_INST_DATA_PATH_DECODE_RF_n5554, 
      DLX_INST_DATA_PATH_DECODE_RF_n5553, DLX_INST_DATA_PATH_DECODE_RF_n5552, 
      DLX_INST_DATA_PATH_DECODE_RF_n5551, DLX_INST_DATA_PATH_DECODE_RF_n5550, 
      DLX_INST_DATA_PATH_DECODE_RF_n5549, DLX_INST_DATA_PATH_DECODE_RF_n5548, 
      DLX_INST_DATA_PATH_DECODE_RF_n5547, DLX_INST_DATA_PATH_DECODE_RF_n5546, 
      DLX_INST_DATA_PATH_DECODE_RF_n5545, DLX_INST_DATA_PATH_DECODE_RF_n5544, 
      DLX_INST_DATA_PATH_DECODE_RF_n5543, DLX_INST_DATA_PATH_DECODE_RF_n5542, 
      DLX_INST_DATA_PATH_DECODE_RF_n5541, DLX_INST_DATA_PATH_DECODE_RF_n5540, 
      DLX_INST_DATA_PATH_DECODE_RF_n5539, DLX_INST_DATA_PATH_DECODE_RF_n5538, 
      DLX_INST_DATA_PATH_DECODE_RF_n5537, DLX_INST_DATA_PATH_DECODE_RF_n5536, 
      DLX_INST_DATA_PATH_DECODE_RF_n5535, DLX_INST_DATA_PATH_DECODE_RF_n5534, 
      DLX_INST_DATA_PATH_DECODE_RF_n5533, DLX_INST_DATA_PATH_DECODE_RF_n5532, 
      DLX_INST_DATA_PATH_DECODE_RF_n5531, DLX_INST_DATA_PATH_DECODE_RF_n5530, 
      DLX_INST_DATA_PATH_DECODE_RF_n5529, DLX_INST_DATA_PATH_DECODE_RF_n5528, 
      DLX_INST_DATA_PATH_DECODE_RF_n5527, DLX_INST_DATA_PATH_DECODE_RF_n5526, 
      DLX_INST_DATA_PATH_DECODE_RF_n5525, DLX_INST_DATA_PATH_DECODE_RF_n5524, 
      DLX_INST_DATA_PATH_DECODE_RF_n5523, DLX_INST_DATA_PATH_DECODE_RF_n5522, 
      DLX_INST_DATA_PATH_DECODE_RF_n5521, DLX_INST_DATA_PATH_DECODE_RF_n5520, 
      DLX_INST_DATA_PATH_DECODE_RF_n5519, DLX_INST_DATA_PATH_DECODE_RF_n5518, 
      DLX_INST_DATA_PATH_DECODE_RF_n5517, DLX_INST_DATA_PATH_DECODE_RF_n5516, 
      DLX_INST_DATA_PATH_DECODE_RF_n5515, DLX_INST_DATA_PATH_DECODE_RF_n5514, 
      DLX_INST_DATA_PATH_DECODE_RF_n5513, DLX_INST_DATA_PATH_DECODE_RF_n5512, 
      DLX_INST_DATA_PATH_DECODE_RF_n5511, DLX_INST_DATA_PATH_DECODE_RF_n5510, 
      DLX_INST_DATA_PATH_DECODE_RF_n5509, DLX_INST_DATA_PATH_DECODE_RF_n5508, 
      DLX_INST_DATA_PATH_DECODE_RF_n5507, DLX_INST_DATA_PATH_DECODE_RF_n5506, 
      DLX_INST_DATA_PATH_DECODE_RF_n5505, DLX_INST_DATA_PATH_DECODE_RF_n5504, 
      DLX_INST_DATA_PATH_DECODE_RF_n5503, DLX_INST_DATA_PATH_DECODE_RF_n5502, 
      DLX_INST_DATA_PATH_DECODE_RF_n5501, DLX_INST_DATA_PATH_DECODE_RF_n5500, 
      DLX_INST_DATA_PATH_DECODE_RF_n5499, DLX_INST_DATA_PATH_DECODE_RF_n5498, 
      DLX_INST_DATA_PATH_DECODE_RF_n5497, DLX_INST_DATA_PATH_DECODE_RF_n5496, 
      DLX_INST_DATA_PATH_DECODE_RF_n5495, DLX_INST_DATA_PATH_DECODE_RF_n5494, 
      DLX_INST_DATA_PATH_DECODE_RF_n5493, DLX_INST_DATA_PATH_DECODE_RF_n5492, 
      DLX_INST_DATA_PATH_DECODE_RF_n5491, DLX_INST_DATA_PATH_DECODE_RF_n5490, 
      DLX_INST_DATA_PATH_DECODE_RF_n5489, DLX_INST_DATA_PATH_DECODE_RF_n5488, 
      DLX_INST_DATA_PATH_DECODE_RF_n5487, DLX_INST_DATA_PATH_DECODE_RF_n5486, 
      DLX_INST_DATA_PATH_DECODE_RF_n5485, DLX_INST_DATA_PATH_DECODE_RF_n5484, 
      DLX_INST_DATA_PATH_DECODE_RF_n5483, DLX_INST_DATA_PATH_DECODE_RF_n5482, 
      DLX_INST_DATA_PATH_DECODE_RF_n5481, DLX_INST_DATA_PATH_DECODE_RF_n5480, 
      DLX_INST_DATA_PATH_DECODE_RF_n5479, DLX_INST_DATA_PATH_DECODE_RF_n5478, 
      DLX_INST_DATA_PATH_DECODE_RF_n5477, DLX_INST_DATA_PATH_DECODE_RF_n5476, 
      DLX_INST_DATA_PATH_DECODE_RF_n5475, DLX_INST_DATA_PATH_DECODE_RF_n5474, 
      DLX_INST_DATA_PATH_DECODE_RF_n5473, DLX_INST_DATA_PATH_DECODE_RF_n5472, 
      DLX_INST_DATA_PATH_DECODE_RF_n5471, DLX_INST_DATA_PATH_DECODE_RF_n5470, 
      DLX_INST_DATA_PATH_DECODE_RF_n5469, DLX_INST_DATA_PATH_DECODE_RF_n5468, 
      DLX_INST_DATA_PATH_DECODE_RF_n5467, DLX_INST_DATA_PATH_DECODE_RF_n5466, 
      DLX_INST_DATA_PATH_DECODE_RF_n5465, DLX_INST_DATA_PATH_DECODE_RF_n5464, 
      DLX_INST_DATA_PATH_DECODE_RF_n5463, DLX_INST_DATA_PATH_DECODE_RF_n5462, 
      DLX_INST_DATA_PATH_DECODE_RF_n5461, DLX_INST_DATA_PATH_DECODE_RF_n5460, 
      DLX_INST_DATA_PATH_DECODE_RF_n5459, DLX_INST_DATA_PATH_DECODE_RF_n5458, 
      DLX_INST_DATA_PATH_DECODE_RF_n5457, DLX_INST_DATA_PATH_DECODE_RF_n5456, 
      DLX_INST_DATA_PATH_DECODE_RF_n5455, DLX_INST_DATA_PATH_DECODE_RF_n5454, 
      DLX_INST_DATA_PATH_DECODE_RF_n5453, DLX_INST_DATA_PATH_DECODE_RF_n5452, 
      DLX_INST_DATA_PATH_DECODE_RF_n5451, DLX_INST_DATA_PATH_DECODE_RF_n5450, 
      DLX_INST_DATA_PATH_DECODE_RF_n5449, DLX_INST_DATA_PATH_DECODE_RF_n5448, 
      DLX_INST_DATA_PATH_DECODE_RF_n5447, DLX_INST_DATA_PATH_DECODE_RF_n5446, 
      DLX_INST_DATA_PATH_DECODE_RF_n5445, DLX_INST_DATA_PATH_DECODE_RF_n5444, 
      DLX_INST_DATA_PATH_DECODE_RF_n5443, DLX_INST_DATA_PATH_DECODE_RF_n5442, 
      DLX_INST_DATA_PATH_DECODE_RF_n5441, DLX_INST_DATA_PATH_DECODE_RF_n5440, 
      DLX_INST_DATA_PATH_DECODE_RF_n5439, DLX_INST_DATA_PATH_DECODE_RF_n5438, 
      DLX_INST_DATA_PATH_DECODE_RF_n5437, DLX_INST_DATA_PATH_DECODE_RF_n5436, 
      DLX_INST_DATA_PATH_DECODE_RF_n5435, DLX_INST_DATA_PATH_DECODE_RF_n5434, 
      DLX_INST_DATA_PATH_DECODE_RF_n5433, DLX_INST_DATA_PATH_DECODE_RF_n5432, 
      DLX_INST_DATA_PATH_DECODE_RF_n5431, DLX_INST_DATA_PATH_DECODE_RF_n5430, 
      DLX_INST_DATA_PATH_DECODE_RF_n5429, DLX_INST_DATA_PATH_DECODE_RF_n5428, 
      DLX_INST_DATA_PATH_DECODE_RF_n5427, DLX_INST_DATA_PATH_DECODE_RF_n5426, 
      DLX_INST_DATA_PATH_DECODE_RF_n5425, DLX_INST_DATA_PATH_DECODE_RF_n5424, 
      DLX_INST_DATA_PATH_DECODE_RF_n5423, DLX_INST_DATA_PATH_DECODE_RF_n5422, 
      DLX_INST_DATA_PATH_DECODE_RF_n5421, DLX_INST_DATA_PATH_DECODE_RF_n5420, 
      DLX_INST_DATA_PATH_DECODE_RF_n5419, DLX_INST_DATA_PATH_DECODE_RF_n5418, 
      DLX_INST_DATA_PATH_DECODE_RF_n5417, DLX_INST_DATA_PATH_DECODE_RF_n5416, 
      DLX_INST_DATA_PATH_DECODE_RF_n5415, DLX_INST_DATA_PATH_DECODE_RF_n5414, 
      DLX_INST_DATA_PATH_DECODE_RF_n5413, DLX_INST_DATA_PATH_DECODE_RF_n5412, 
      DLX_INST_DATA_PATH_DECODE_RF_n5411, DLX_INST_DATA_PATH_DECODE_RF_n5410, 
      DLX_INST_DATA_PATH_DECODE_RF_n5409, DLX_INST_DATA_PATH_DECODE_RF_n5408, 
      DLX_INST_DATA_PATH_DECODE_RF_n5407, DLX_INST_DATA_PATH_DECODE_RF_n5406, 
      DLX_INST_DATA_PATH_DECODE_RF_n5405, DLX_INST_DATA_PATH_DECODE_RF_n5404, 
      DLX_INST_DATA_PATH_DECODE_RF_n5403, DLX_INST_DATA_PATH_DECODE_RF_n5402, 
      DLX_INST_DATA_PATH_DECODE_RF_n5401, DLX_INST_DATA_PATH_DECODE_RF_n5400, 
      DLX_INST_DATA_PATH_DECODE_RF_n5399, DLX_INST_DATA_PATH_DECODE_RF_n5398, 
      DLX_INST_DATA_PATH_DECODE_RF_n5397, DLX_INST_DATA_PATH_DECODE_RF_n5396, 
      DLX_INST_DATA_PATH_DECODE_RF_n5395, DLX_INST_DATA_PATH_DECODE_RF_n5394, 
      DLX_INST_DATA_PATH_DECODE_RF_n5393, DLX_INST_DATA_PATH_DECODE_RF_n5392, 
      DLX_INST_DATA_PATH_DECODE_RF_n5391, DLX_INST_DATA_PATH_DECODE_RF_n5390, 
      DLX_INST_DATA_PATH_DECODE_RF_n5389, DLX_INST_DATA_PATH_DECODE_RF_n5388, 
      DLX_INST_DATA_PATH_DECODE_RF_n5387, DLX_INST_DATA_PATH_DECODE_RF_n5386, 
      DLX_INST_DATA_PATH_DECODE_RF_n5385, DLX_INST_DATA_PATH_DECODE_RF_n5384, 
      DLX_INST_DATA_PATH_DECODE_RF_n5383, DLX_INST_DATA_PATH_DECODE_RF_n5382, 
      DLX_INST_DATA_PATH_DECODE_RF_n5381, DLX_INST_DATA_PATH_DECODE_RF_n5380, 
      DLX_INST_DATA_PATH_DECODE_RF_n5379, DLX_INST_DATA_PATH_DECODE_RF_n5378, 
      DLX_INST_DATA_PATH_DECODE_RF_n5377, DLX_INST_DATA_PATH_DECODE_RF_n5376, 
      DLX_INST_DATA_PATH_DECODE_RF_n5375, DLX_INST_DATA_PATH_DECODE_RF_n5374, 
      DLX_INST_DATA_PATH_DECODE_RF_n5373, DLX_INST_DATA_PATH_DECODE_RF_n5372, 
      DLX_INST_DATA_PATH_DECODE_RF_n5371, DLX_INST_DATA_PATH_DECODE_RF_n5370, 
      DLX_INST_DATA_PATH_DECODE_RF_n5369, DLX_INST_DATA_PATH_DECODE_RF_n5368, 
      DLX_INST_DATA_PATH_DECODE_RF_n5367, DLX_INST_DATA_PATH_DECODE_RF_n5366, 
      DLX_INST_DATA_PATH_DECODE_RF_n5365, DLX_INST_DATA_PATH_DECODE_RF_n5364, 
      DLX_INST_DATA_PATH_DECODE_RF_n5363, DLX_INST_DATA_PATH_DECODE_RF_n5362, 
      DLX_INST_DATA_PATH_DECODE_RF_n5361, DLX_INST_DATA_PATH_DECODE_RF_n5360, 
      DLX_INST_DATA_PATH_DECODE_RF_n5359, DLX_INST_DATA_PATH_DECODE_RF_n5358, 
      DLX_INST_DATA_PATH_DECODE_RF_n5357, DLX_INST_DATA_PATH_DECODE_RF_n5356, 
      DLX_INST_DATA_PATH_DECODE_RF_n5355, DLX_INST_DATA_PATH_DECODE_RF_n5354, 
      DLX_INST_DATA_PATH_DECODE_RF_n5353, DLX_INST_DATA_PATH_DECODE_RF_n5352, 
      DLX_INST_DATA_PATH_DECODE_RF_n5351, DLX_INST_DATA_PATH_DECODE_RF_n5350, 
      DLX_INST_DATA_PATH_DECODE_RF_n5349, DLX_INST_DATA_PATH_DECODE_RF_n5348, 
      DLX_INST_DATA_PATH_DECODE_RF_n5347, DLX_INST_DATA_PATH_DECODE_RF_n5346, 
      DLX_INST_DATA_PATH_DECODE_RF_n5345, DLX_INST_DATA_PATH_DECODE_RF_n5344, 
      DLX_INST_DATA_PATH_DECODE_RF_n5343, DLX_INST_DATA_PATH_DECODE_RF_n5342, 
      DLX_INST_DATA_PATH_DECODE_RF_n5341, DLX_INST_DATA_PATH_DECODE_RF_n5340, 
      DLX_INST_DATA_PATH_DECODE_RF_n5339, DLX_INST_DATA_PATH_DECODE_RF_n5338, 
      DLX_INST_DATA_PATH_DECODE_RF_n5337, DLX_INST_DATA_PATH_DECODE_RF_n5336, 
      DLX_INST_DATA_PATH_DECODE_RF_n5335, DLX_INST_DATA_PATH_DECODE_RF_n5334, 
      DLX_INST_DATA_PATH_DECODE_RF_n5333, DLX_INST_DATA_PATH_DECODE_RF_n5332, 
      DLX_INST_DATA_PATH_DECODE_RF_n5331, DLX_INST_DATA_PATH_DECODE_RF_n5330, 
      DLX_INST_DATA_PATH_DECODE_RF_n5329, DLX_INST_DATA_PATH_DECODE_RF_n5328, 
      DLX_INST_DATA_PATH_DECODE_RF_n5327, DLX_INST_DATA_PATH_DECODE_RF_n5326, 
      DLX_INST_DATA_PATH_DECODE_RF_n5325, DLX_INST_DATA_PATH_DECODE_RF_n5324, 
      DLX_INST_DATA_PATH_DECODE_RF_n5323, DLX_INST_DATA_PATH_DECODE_RF_n5322, 
      DLX_INST_DATA_PATH_DECODE_RF_n5321, DLX_INST_DATA_PATH_DECODE_RF_n5320, 
      DLX_INST_DATA_PATH_DECODE_RF_n5319, DLX_INST_DATA_PATH_DECODE_RF_n5318, 
      DLX_INST_DATA_PATH_DECODE_RF_n5317, DLX_INST_DATA_PATH_DECODE_RF_n5316, 
      DLX_INST_DATA_PATH_DECODE_RF_n5315, DLX_INST_DATA_PATH_DECODE_RF_n5314, 
      DLX_INST_DATA_PATH_DECODE_RF_n5313, DLX_INST_DATA_PATH_DECODE_RF_n5312, 
      DLX_INST_DATA_PATH_DECODE_RF_n5311, DLX_INST_DATA_PATH_DECODE_RF_n5310, 
      DLX_INST_DATA_PATH_DECODE_RF_n5309, DLX_INST_DATA_PATH_DECODE_RF_n5308, 
      DLX_INST_DATA_PATH_DECODE_RF_n5307, DLX_INST_DATA_PATH_DECODE_RF_n5306, 
      DLX_INST_DATA_PATH_DECODE_RF_n5305, DLX_INST_DATA_PATH_DECODE_RF_n5304, 
      DLX_INST_DATA_PATH_DECODE_RF_n5303, DLX_INST_DATA_PATH_DECODE_RF_n5302, 
      DLX_INST_DATA_PATH_DECODE_RF_n5301, DLX_INST_DATA_PATH_DECODE_RF_n5300, 
      DLX_INST_DATA_PATH_DECODE_RF_n5299, DLX_INST_DATA_PATH_DECODE_RF_n5298, 
      DLX_INST_DATA_PATH_DECODE_RF_n5297, DLX_INST_DATA_PATH_DECODE_RF_n5296, 
      DLX_INST_DATA_PATH_DECODE_RF_n5295, DLX_INST_DATA_PATH_DECODE_RF_n5294, 
      DLX_INST_DATA_PATH_DECODE_RF_n5293, DLX_INST_DATA_PATH_DECODE_RF_n5292, 
      DLX_INST_DATA_PATH_DECODE_RF_n5291, DLX_INST_DATA_PATH_DECODE_RF_n5290, 
      DLX_INST_DATA_PATH_DECODE_RF_n5289, DLX_INST_DATA_PATH_DECODE_RF_n5288, 
      DLX_INST_DATA_PATH_DECODE_RF_n5287, DLX_INST_DATA_PATH_DECODE_RF_n5286, 
      DLX_INST_DATA_PATH_DECODE_RF_n5285, DLX_INST_DATA_PATH_DECODE_RF_n5284, 
      DLX_INST_DATA_PATH_DECODE_RF_n5283, DLX_INST_DATA_PATH_DECODE_RF_n5282, 
      DLX_INST_DATA_PATH_DECODE_RF_n5281, DLX_INST_DATA_PATH_DECODE_RF_n5280, 
      DLX_INST_DATA_PATH_DECODE_RF_n5279, DLX_INST_DATA_PATH_DECODE_RF_n5278, 
      DLX_INST_DATA_PATH_DECODE_RF_n5277, DLX_INST_DATA_PATH_DECODE_RF_n5276, 
      DLX_INST_DATA_PATH_DECODE_RF_n5275, DLX_INST_DATA_PATH_DECODE_RF_n5274, 
      DLX_INST_DATA_PATH_DECODE_RF_n5273, DLX_INST_DATA_PATH_DECODE_RF_n5272, 
      DLX_INST_DATA_PATH_DECODE_RF_n5271, DLX_INST_DATA_PATH_DECODE_RF_n5270, 
      DLX_INST_DATA_PATH_DECODE_RF_n5269, DLX_INST_DATA_PATH_DECODE_RF_n5268, 
      DLX_INST_DATA_PATH_DECODE_RF_n5267, DLX_INST_DATA_PATH_DECODE_RF_n5266, 
      DLX_INST_DATA_PATH_DECODE_RF_n5265, DLX_INST_DATA_PATH_DECODE_RF_n5264, 
      DLX_INST_DATA_PATH_DECODE_RF_n5263, DLX_INST_DATA_PATH_DECODE_RF_n5262, 
      DLX_INST_DATA_PATH_DECODE_RF_n5261, DLX_INST_DATA_PATH_DECODE_RF_n5260, 
      DLX_INST_DATA_PATH_DECODE_RF_n5259, DLX_INST_DATA_PATH_DECODE_RF_n5258, 
      DLX_INST_DATA_PATH_DECODE_RF_n5257, DLX_INST_DATA_PATH_DECODE_RF_n5256, 
      DLX_INST_DATA_PATH_DECODE_RF_n5255, DLX_INST_DATA_PATH_DECODE_RF_n5254, 
      DLX_INST_DATA_PATH_DECODE_RF_n5253, DLX_INST_DATA_PATH_DECODE_RF_n5252, 
      DLX_INST_DATA_PATH_DECODE_RF_n5251, DLX_INST_DATA_PATH_DECODE_RF_n5250, 
      DLX_INST_DATA_PATH_DECODE_RF_n5249, DLX_INST_DATA_PATH_DECODE_RF_n5248, 
      DLX_INST_DATA_PATH_DECODE_RF_n5247, DLX_INST_DATA_PATH_DECODE_RF_n5246, 
      DLX_INST_DATA_PATH_DECODE_RF_n5245, DLX_INST_DATA_PATH_DECODE_RF_n5244, 
      DLX_INST_DATA_PATH_DECODE_RF_n5243, DLX_INST_DATA_PATH_DECODE_RF_n5242, 
      DLX_INST_DATA_PATH_DECODE_RF_n5241, DLX_INST_DATA_PATH_DECODE_RF_n5240, 
      DLX_INST_DATA_PATH_DECODE_RF_n5239, DLX_INST_DATA_PATH_DECODE_RF_n5238, 
      DLX_INST_DATA_PATH_DECODE_RF_n5237, DLX_INST_DATA_PATH_DECODE_RF_n5236, 
      DLX_INST_DATA_PATH_DECODE_RF_n5235, DLX_INST_DATA_PATH_DECODE_RF_n5234, 
      DLX_INST_DATA_PATH_DECODE_RF_n5233, DLX_INST_DATA_PATH_DECODE_RF_n5232, 
      DLX_INST_DATA_PATH_DECODE_RF_n5231, DLX_INST_DATA_PATH_DECODE_RF_n5230, 
      DLX_INST_DATA_PATH_DECODE_RF_n5229, DLX_INST_DATA_PATH_DECODE_RF_n5228, 
      DLX_INST_DATA_PATH_DECODE_RF_n5227, DLX_INST_DATA_PATH_DECODE_RF_n5226, 
      DLX_INST_DATA_PATH_DECODE_RF_n5225, DLX_INST_DATA_PATH_DECODE_RF_n5224, 
      DLX_INST_DATA_PATH_DECODE_RF_n5223, DLX_INST_DATA_PATH_DECODE_RF_n5222, 
      DLX_INST_DATA_PATH_DECODE_RF_n5221, DLX_INST_DATA_PATH_DECODE_RF_n5220, 
      DLX_INST_DATA_PATH_DECODE_RF_n5219, DLX_INST_DATA_PATH_DECODE_RF_n5218, 
      DLX_INST_DATA_PATH_DECODE_RF_n5217, DLX_INST_DATA_PATH_DECODE_RF_n5216, 
      DLX_INST_DATA_PATH_DECODE_RF_n5215, DLX_INST_DATA_PATH_DECODE_RF_n5214, 
      DLX_INST_DATA_PATH_DECODE_RF_n5213, DLX_INST_DATA_PATH_DECODE_RF_n5212, 
      DLX_INST_DATA_PATH_DECODE_RF_n5211, DLX_INST_DATA_PATH_DECODE_RF_n5210, 
      DLX_INST_DATA_PATH_DECODE_RF_n5209, DLX_INST_DATA_PATH_DECODE_RF_n5208, 
      DLX_INST_DATA_PATH_DECODE_RF_n5207, DLX_INST_DATA_PATH_DECODE_RF_n5206, 
      DLX_INST_DATA_PATH_DECODE_RF_n5205, DLX_INST_DATA_PATH_DECODE_RF_n5204, 
      DLX_INST_DATA_PATH_DECODE_RF_n5203, DLX_INST_DATA_PATH_DECODE_RF_n5202, 
      DLX_INST_DATA_PATH_DECODE_RF_n5201, DLX_INST_DATA_PATH_DECODE_RF_n5200, 
      DLX_INST_DATA_PATH_DECODE_RF_n5199, DLX_INST_DATA_PATH_DECODE_RF_n5198, 
      DLX_INST_DATA_PATH_DECODE_RF_n5197, DLX_INST_DATA_PATH_DECODE_RF_n5196, 
      DLX_INST_DATA_PATH_DECODE_RF_n5195, DLX_INST_DATA_PATH_DECODE_RF_n5194, 
      DLX_INST_DATA_PATH_DECODE_RF_n5193, DLX_INST_DATA_PATH_DECODE_RF_n5192, 
      DLX_INST_DATA_PATH_DECODE_RF_n5191, DLX_INST_DATA_PATH_DECODE_RF_n5190, 
      DLX_INST_DATA_PATH_DECODE_RF_n5189, DLX_INST_DATA_PATH_DECODE_RF_n5188, 
      DLX_INST_DATA_PATH_DECODE_RF_n5187, DLX_INST_DATA_PATH_DECODE_RF_n5186, 
      DLX_INST_DATA_PATH_DECODE_RF_n5185, DLX_INST_DATA_PATH_DECODE_RF_n5184, 
      DLX_INST_DATA_PATH_DECODE_RF_n5183, DLX_INST_DATA_PATH_DECODE_RF_n5182, 
      DLX_INST_DATA_PATH_DECODE_RF_n5181, DLX_INST_DATA_PATH_DECODE_RF_n5180, 
      DLX_INST_DATA_PATH_DECODE_RF_n5179, DLX_INST_DATA_PATH_DECODE_RF_n5178, 
      DLX_INST_DATA_PATH_DECODE_RF_n5177, DLX_INST_DATA_PATH_DECODE_RF_n5176, 
      DLX_INST_DATA_PATH_DECODE_RF_n5175, DLX_INST_DATA_PATH_DECODE_RF_n5174, 
      DLX_INST_DATA_PATH_DECODE_RF_n5173, DLX_INST_DATA_PATH_DECODE_RF_n5172, 
      DLX_INST_DATA_PATH_DECODE_RF_n5171, DLX_INST_DATA_PATH_DECODE_RF_n5170, 
      DLX_INST_DATA_PATH_DECODE_RF_n5169, DLX_INST_DATA_PATH_DECODE_RF_n5168, 
      DLX_INST_DATA_PATH_DECODE_RF_n5167, DLX_INST_DATA_PATH_DECODE_RF_n5166, 
      DLX_INST_DATA_PATH_DECODE_RF_n5165, DLX_INST_DATA_PATH_DECODE_RF_n5164, 
      DLX_INST_DATA_PATH_DECODE_RF_n5163, DLX_INST_DATA_PATH_DECODE_RF_n5162, 
      DLX_INST_DATA_PATH_DECODE_RF_n5161, DLX_INST_DATA_PATH_DECODE_RF_n5160, 
      DLX_INST_DATA_PATH_DECODE_RF_n5159, DLX_INST_DATA_PATH_DECODE_RF_n5158, 
      DLX_INST_DATA_PATH_DECODE_RF_n5157, DLX_INST_DATA_PATH_DECODE_RF_n5156, 
      DLX_INST_DATA_PATH_DECODE_RF_n5155, DLX_INST_DATA_PATH_DECODE_RF_n5154, 
      DLX_INST_DATA_PATH_DECODE_RF_n5153, DLX_INST_DATA_PATH_DECODE_RF_n5152, 
      DLX_INST_DATA_PATH_DECODE_RF_n5151, DLX_INST_DATA_PATH_DECODE_RF_n5150, 
      DLX_INST_DATA_PATH_DECODE_RF_n5149, DLX_INST_DATA_PATH_DECODE_RF_n5148, 
      DLX_INST_DATA_PATH_DECODE_RF_n5147, DLX_INST_DATA_PATH_DECODE_RF_n5146, 
      DLX_INST_DATA_PATH_DECODE_RF_n5145, DLX_INST_DATA_PATH_DECODE_RF_n5144, 
      DLX_INST_DATA_PATH_DECODE_RF_n5143, DLX_INST_DATA_PATH_DECODE_RF_n5142, 
      DLX_INST_DATA_PATH_DECODE_RF_n5141, DLX_INST_DATA_PATH_DECODE_RF_n5140, 
      DLX_INST_DATA_PATH_DECODE_RF_n5139, DLX_INST_DATA_PATH_DECODE_RF_n5138, 
      DLX_INST_DATA_PATH_DECODE_RF_n5137, DLX_INST_DATA_PATH_DECODE_RF_n5136, 
      DLX_INST_DATA_PATH_DECODE_RF_n5135, DLX_INST_DATA_PATH_DECODE_RF_n5134, 
      DLX_INST_DATA_PATH_DECODE_RF_n5133, DLX_INST_DATA_PATH_DECODE_RF_n5132, 
      DLX_INST_DATA_PATH_DECODE_RF_n5131, DLX_INST_DATA_PATH_DECODE_RF_n5130, 
      DLX_INST_DATA_PATH_DECODE_RF_n5129, DLX_INST_DATA_PATH_DECODE_RF_n5128, 
      DLX_INST_DATA_PATH_DECODE_RF_n5127, DLX_INST_DATA_PATH_DECODE_RF_n5126, 
      DLX_INST_DATA_PATH_DECODE_RF_n5125, DLX_INST_DATA_PATH_DECODE_RF_n5124, 
      DLX_INST_DATA_PATH_DECODE_RF_n5123, DLX_INST_DATA_PATH_DECODE_RF_n5122, 
      DLX_INST_DATA_PATH_DECODE_RF_n5121, DLX_INST_DATA_PATH_DECODE_RF_n5120, 
      DLX_INST_DATA_PATH_DECODE_RF_n5119, DLX_INST_DATA_PATH_DECODE_RF_n5118, 
      DLX_INST_DATA_PATH_DECODE_RF_n5117, DLX_INST_DATA_PATH_DECODE_RF_n5116, 
      DLX_INST_DATA_PATH_DECODE_RF_n5115, DLX_INST_DATA_PATH_DECODE_RF_n5114, 
      DLX_INST_DATA_PATH_DECODE_RF_n5113, DLX_INST_DATA_PATH_DECODE_RF_n5112, 
      DLX_INST_DATA_PATH_DECODE_RF_n5111, DLX_INST_DATA_PATH_DECODE_RF_n5110, 
      DLX_INST_DATA_PATH_DECODE_RF_n5109, DLX_INST_DATA_PATH_DECODE_RF_n5108, 
      DLX_INST_DATA_PATH_DECODE_RF_n5107, DLX_INST_DATA_PATH_DECODE_RF_n5106, 
      DLX_INST_DATA_PATH_DECODE_RF_n5105, DLX_INST_DATA_PATH_DECODE_RF_n5104, 
      DLX_INST_DATA_PATH_DECODE_RF_n5103, DLX_INST_DATA_PATH_DECODE_RF_n5102, 
      DLX_INST_DATA_PATH_DECODE_RF_n5101, DLX_INST_DATA_PATH_DECODE_RF_n5100, 
      DLX_INST_DATA_PATH_DECODE_RF_n5099, DLX_INST_DATA_PATH_DECODE_RF_n5098, 
      DLX_INST_DATA_PATH_DECODE_RF_n5097, DLX_INST_DATA_PATH_DECODE_RF_n5096, 
      DLX_INST_DATA_PATH_DECODE_RF_n5095, DLX_INST_DATA_PATH_DECODE_RF_n5094, 
      DLX_INST_DATA_PATH_DECODE_RF_n5093, DLX_INST_DATA_PATH_DECODE_RF_n5092, 
      DLX_INST_DATA_PATH_DECODE_RF_n5091, DLX_INST_DATA_PATH_DECODE_RF_n5090, 
      DLX_INST_DATA_PATH_DECODE_RF_n5089, DLX_INST_DATA_PATH_DECODE_RF_n5088, 
      DLX_INST_DATA_PATH_DECODE_RF_n5087, DLX_INST_DATA_PATH_DECODE_RF_n5086, 
      DLX_INST_DATA_PATH_DECODE_RF_n5085, DLX_INST_DATA_PATH_DECODE_RF_n5084, 
      DLX_INST_DATA_PATH_DECODE_RF_n5083, DLX_INST_DATA_PATH_DECODE_RF_n5082, 
      DLX_INST_DATA_PATH_DECODE_RF_n5081, DLX_INST_DATA_PATH_DECODE_RF_n5080, 
      DLX_INST_DATA_PATH_DECODE_RF_n5079, DLX_INST_DATA_PATH_DECODE_RF_n5078, 
      DLX_INST_DATA_PATH_DECODE_RF_n5077, DLX_INST_DATA_PATH_DECODE_RF_n5076, 
      DLX_INST_DATA_PATH_DECODE_RF_n5075, DLX_INST_DATA_PATH_DECODE_RF_n5074, 
      DLX_INST_DATA_PATH_DECODE_RF_n5073, DLX_INST_DATA_PATH_DECODE_RF_n5072, 
      DLX_INST_DATA_PATH_DECODE_RF_n5071, DLX_INST_DATA_PATH_DECODE_RF_n5070, 
      DLX_INST_DATA_PATH_DECODE_RF_n5069, DLX_INST_DATA_PATH_DECODE_RF_n5068, 
      DLX_INST_DATA_PATH_DECODE_RF_n5067, DLX_INST_DATA_PATH_DECODE_RF_n5066, 
      DLX_INST_DATA_PATH_DECODE_RF_n5065, DLX_INST_DATA_PATH_DECODE_RF_n5064, 
      DLX_INST_DATA_PATH_DECODE_RF_n5063, DLX_INST_DATA_PATH_DECODE_RF_n5062, 
      DLX_INST_DATA_PATH_DECODE_RF_n5061, DLX_INST_DATA_PATH_DECODE_RF_n5060, 
      DLX_INST_DATA_PATH_DECODE_RF_n5059, DLX_INST_DATA_PATH_DECODE_RF_n5058, 
      DLX_INST_DATA_PATH_DECODE_RF_n5057, DLX_INST_DATA_PATH_DECODE_RF_n5056, 
      DLX_INST_DATA_PATH_DECODE_RF_n5055, DLX_INST_DATA_PATH_DECODE_RF_n5054, 
      DLX_INST_DATA_PATH_DECODE_RF_n5053, DLX_INST_DATA_PATH_DECODE_RF_n5052, 
      DLX_INST_DATA_PATH_DECODE_RF_n5051, DLX_INST_DATA_PATH_DECODE_RF_n5050, 
      DLX_INST_DATA_PATH_DECODE_RF_n5049, DLX_INST_DATA_PATH_DECODE_RF_n5048, 
      DLX_INST_DATA_PATH_DECODE_RF_n5047, DLX_INST_DATA_PATH_DECODE_RF_n5046, 
      DLX_INST_DATA_PATH_DECODE_RF_n5045, DLX_INST_DATA_PATH_DECODE_RF_n5044, 
      DLX_INST_DATA_PATH_DECODE_RF_n5043, DLX_INST_DATA_PATH_DECODE_RF_n5042, 
      DLX_INST_DATA_PATH_DECODE_RF_n5041, DLX_INST_DATA_PATH_DECODE_RF_n5040, 
      DLX_INST_DATA_PATH_DECODE_RF_n5039, DLX_INST_DATA_PATH_DECODE_RF_n5038, 
      DLX_INST_DATA_PATH_DECODE_RF_n5037, DLX_INST_DATA_PATH_DECODE_RF_n5036, 
      DLX_INST_DATA_PATH_DECODE_RF_n5035, DLX_INST_DATA_PATH_DECODE_RF_n5034, 
      DLX_INST_DATA_PATH_DECODE_RF_n5033, DLX_INST_DATA_PATH_DECODE_RF_n5032, 
      DLX_INST_DATA_PATH_DECODE_RF_n5031, DLX_INST_DATA_PATH_DECODE_RF_n5030, 
      DLX_INST_DATA_PATH_DECODE_RF_n5029, DLX_INST_DATA_PATH_DECODE_RF_n5028, 
      DLX_INST_DATA_PATH_DECODE_RF_n5027, DLX_INST_DATA_PATH_DECODE_RF_n5026, 
      DLX_INST_DATA_PATH_DECODE_RF_n5025, DLX_INST_DATA_PATH_DECODE_RF_n5024, 
      DLX_INST_DATA_PATH_DECODE_RF_n5023, DLX_INST_DATA_PATH_DECODE_RF_n5022, 
      DLX_INST_DATA_PATH_DECODE_RF_n5021, DLX_INST_DATA_PATH_DECODE_RF_n5020, 
      DLX_INST_DATA_PATH_DECODE_RF_n5019, DLX_INST_DATA_PATH_DECODE_RF_n5018, 
      DLX_INST_DATA_PATH_DECODE_RF_n5017, DLX_INST_DATA_PATH_DECODE_RF_n5016, 
      DLX_INST_DATA_PATH_DECODE_RF_n5015, DLX_INST_DATA_PATH_DECODE_RF_n5014, 
      DLX_INST_DATA_PATH_DECODE_RF_n5013, DLX_INST_DATA_PATH_DECODE_RF_n5012, 
      DLX_INST_DATA_PATH_DECODE_RF_n5011, DLX_INST_DATA_PATH_DECODE_RF_n5010, 
      DLX_INST_DATA_PATH_DECODE_RF_n5009, DLX_INST_DATA_PATH_DECODE_RF_n5008, 
      DLX_INST_DATA_PATH_DECODE_RF_n5007, DLX_INST_DATA_PATH_DECODE_RF_n5006, 
      DLX_INST_DATA_PATH_DECODE_RF_n5005, DLX_INST_DATA_PATH_DECODE_RF_n5004, 
      DLX_INST_DATA_PATH_DECODE_RF_n5003, DLX_INST_DATA_PATH_DECODE_RF_n5002, 
      DLX_INST_DATA_PATH_DECODE_RF_n5001, DLX_INST_DATA_PATH_DECODE_RF_n5000, 
      DLX_INST_DATA_PATH_DECODE_RF_n4999, DLX_INST_DATA_PATH_DECODE_RF_n4998, 
      DLX_INST_DATA_PATH_DECODE_RF_n4997, DLX_INST_DATA_PATH_DECODE_RF_n4996, 
      DLX_INST_DATA_PATH_DECODE_RF_n4995, DLX_INST_DATA_PATH_DECODE_RF_n4994, 
      DLX_INST_DATA_PATH_DECODE_RF_n4993, DLX_INST_DATA_PATH_DECODE_RF_n4992, 
      DLX_INST_DATA_PATH_DECODE_RF_n4991, DLX_INST_DATA_PATH_DECODE_RF_n4990, 
      DLX_INST_DATA_PATH_DECODE_RF_n4989, DLX_INST_DATA_PATH_DECODE_RF_n4988, 
      DLX_INST_DATA_PATH_DECODE_RF_n4987, DLX_INST_DATA_PATH_DECODE_RF_n4986, 
      DLX_INST_DATA_PATH_DECODE_RF_n4985, DLX_INST_DATA_PATH_DECODE_RF_n4984, 
      DLX_INST_DATA_PATH_DECODE_RF_n4983, DLX_INST_DATA_PATH_DECODE_RF_n4982, 
      DLX_INST_DATA_PATH_DECODE_RF_n4981, DLX_INST_DATA_PATH_DECODE_RF_n4980, 
      DLX_INST_DATA_PATH_DECODE_RF_n4979, DLX_INST_DATA_PATH_DECODE_RF_n4978, 
      DLX_INST_DATA_PATH_DECODE_RF_n4977, DLX_INST_DATA_PATH_DECODE_RF_n4976, 
      DLX_INST_DATA_PATH_DECODE_RF_n4975, DLX_INST_DATA_PATH_DECODE_RF_n4974, 
      DLX_INST_DATA_PATH_DECODE_RF_n4973, DLX_INST_DATA_PATH_DECODE_RF_n4972, 
      DLX_INST_DATA_PATH_DECODE_RF_n4971, DLX_INST_DATA_PATH_DECODE_RF_n4970, 
      DLX_INST_DATA_PATH_DECODE_RF_n4969, DLX_INST_DATA_PATH_DECODE_RF_n4968, 
      DLX_INST_DATA_PATH_DECODE_RF_n4967, DLX_INST_DATA_PATH_DECODE_RF_n4966, 
      DLX_INST_DATA_PATH_DECODE_RF_n4965, DLX_INST_DATA_PATH_DECODE_RF_n4964, 
      DLX_INST_DATA_PATH_DECODE_RF_n4963, DLX_INST_DATA_PATH_DECODE_RF_n4962, 
      DLX_INST_DATA_PATH_DECODE_RF_n4961, DLX_INST_DATA_PATH_DECODE_RF_n4960, 
      DLX_INST_DATA_PATH_DECODE_RF_n4959, DLX_INST_DATA_PATH_DECODE_RF_n4958, 
      DLX_INST_DATA_PATH_DECODE_RF_n4957, DLX_INST_DATA_PATH_DECODE_RF_n4956, 
      DLX_INST_DATA_PATH_DECODE_RF_n4955, DLX_INST_DATA_PATH_DECODE_RF_n4954, 
      DLX_INST_DATA_PATH_DECODE_RF_n4953, DLX_INST_DATA_PATH_DECODE_RF_n4952, 
      DLX_INST_DATA_PATH_DECODE_RF_n4951, DLX_INST_DATA_PATH_DECODE_RF_n4950, 
      DLX_INST_DATA_PATH_DECODE_RF_n4949, DLX_INST_DATA_PATH_DECODE_RF_n4948, 
      DLX_INST_DATA_PATH_DECODE_RF_n4947, DLX_INST_DATA_PATH_DECODE_RF_n4946, 
      DLX_INST_DATA_PATH_DECODE_RF_n4945, DLX_INST_DATA_PATH_DECODE_RF_n4944, 
      DLX_INST_DATA_PATH_DECODE_RF_n4943, DLX_INST_DATA_PATH_DECODE_RF_n4942, 
      DLX_INST_DATA_PATH_DECODE_RF_n4941, DLX_INST_DATA_PATH_DECODE_RF_n4940, 
      DLX_INST_DATA_PATH_DECODE_RF_n4939, DLX_INST_DATA_PATH_DECODE_RF_n4938, 
      DLX_INST_DATA_PATH_DECODE_RF_n4937, DLX_INST_DATA_PATH_DECODE_RF_n4936, 
      DLX_INST_DATA_PATH_DECODE_RF_n4935, DLX_INST_DATA_PATH_DECODE_RF_n4934, 
      DLX_INST_DATA_PATH_DECODE_RF_n4933, DLX_INST_DATA_PATH_DECODE_RF_n4932, 
      DLX_INST_DATA_PATH_DECODE_RF_n4931, DLX_INST_DATA_PATH_DECODE_RF_n4930, 
      DLX_INST_DATA_PATH_DECODE_RF_n4929, DLX_INST_DATA_PATH_DECODE_RF_n4928, 
      DLX_INST_DATA_PATH_DECODE_RF_n4927, DLX_INST_DATA_PATH_DECODE_RF_n4926, 
      DLX_INST_DATA_PATH_DECODE_RF_n4925, DLX_INST_DATA_PATH_DECODE_RF_n4924, 
      DLX_INST_DATA_PATH_DECODE_RF_n4923, DLX_INST_DATA_PATH_DECODE_RF_n4922, 
      DLX_INST_DATA_PATH_DECODE_RF_n4921, DLX_INST_DATA_PATH_DECODE_RF_n4920, 
      DLX_INST_DATA_PATH_DECODE_RF_n4919, DLX_INST_DATA_PATH_DECODE_RF_n4918, 
      DLX_INST_DATA_PATH_DECODE_RF_n4917, DLX_INST_DATA_PATH_DECODE_RF_n4916, 
      DLX_INST_DATA_PATH_DECODE_RF_n4915, DLX_INST_DATA_PATH_DECODE_RF_n4914, 
      DLX_INST_DATA_PATH_DECODE_RF_n4913, DLX_INST_DATA_PATH_DECODE_RF_n4912, 
      DLX_INST_DATA_PATH_DECODE_RF_n4911, DLX_INST_DATA_PATH_DECODE_RF_n4910, 
      DLX_INST_DATA_PATH_DECODE_RF_n4909, DLX_INST_DATA_PATH_DECODE_RF_n4908, 
      DLX_INST_DATA_PATH_DECODE_RF_n4907, DLX_INST_DATA_PATH_DECODE_RF_n4906, 
      DLX_INST_DATA_PATH_DECODE_RF_n4905, DLX_INST_DATA_PATH_DECODE_RF_n4904, 
      DLX_INST_DATA_PATH_DECODE_RF_n4903, DLX_INST_DATA_PATH_DECODE_RF_n4902, 
      DLX_INST_DATA_PATH_DECODE_RF_n4901, DLX_INST_DATA_PATH_DECODE_RF_n4900, 
      DLX_INST_DATA_PATH_DECODE_RF_n4899, DLX_INST_DATA_PATH_DECODE_RF_n4898, 
      DLX_INST_DATA_PATH_DECODE_RF_n4897, DLX_INST_DATA_PATH_DECODE_RF_n4896, 
      DLX_INST_DATA_PATH_DECODE_RF_n4895, DLX_INST_DATA_PATH_DECODE_RF_n4894, 
      DLX_INST_DATA_PATH_DECODE_RF_n4893, DLX_INST_DATA_PATH_DECODE_RF_n4892, 
      DLX_INST_DATA_PATH_DECODE_RF_n4891, DLX_INST_DATA_PATH_DECODE_RF_n4890, 
      DLX_INST_DATA_PATH_DECODE_RF_n4889, DLX_INST_DATA_PATH_DECODE_RF_n4888, 
      DLX_INST_DATA_PATH_DECODE_RF_n4887, DLX_INST_DATA_PATH_DECODE_RF_n4886, 
      DLX_INST_DATA_PATH_DECODE_RF_n4885, DLX_INST_DATA_PATH_DECODE_RF_n4884, 
      DLX_INST_DATA_PATH_DECODE_RF_n4883, DLX_INST_DATA_PATH_DECODE_RF_n4882, 
      DLX_INST_DATA_PATH_DECODE_RF_n4881, DLX_INST_DATA_PATH_DECODE_RF_n4880, 
      DLX_INST_DATA_PATH_DECODE_RF_n4879, DLX_INST_DATA_PATH_DECODE_RF_n4878, 
      DLX_INST_DATA_PATH_DECODE_RF_n4877, DLX_INST_DATA_PATH_DECODE_RF_n4876, 
      DLX_INST_DATA_PATH_DECODE_RF_n4875, DLX_INST_DATA_PATH_DECODE_RF_n4874, 
      DLX_INST_DATA_PATH_DECODE_RF_n4873, DLX_INST_DATA_PATH_DECODE_RF_n4872, 
      DLX_INST_DATA_PATH_DECODE_RF_n4871, DLX_INST_DATA_PATH_DECODE_RF_n4870, 
      DLX_INST_DATA_PATH_DECODE_RF_n4869, DLX_INST_DATA_PATH_DECODE_RF_n4868, 
      DLX_INST_DATA_PATH_DECODE_RF_n4867, DLX_INST_DATA_PATH_DECODE_RF_n4866, 
      DLX_INST_DATA_PATH_DECODE_RF_n4865, DLX_INST_DATA_PATH_DECODE_RF_n4864, 
      DLX_INST_DATA_PATH_DECODE_RF_n4863, DLX_INST_DATA_PATH_DECODE_RF_n4862, 
      DLX_INST_DATA_PATH_DECODE_RF_n4861, DLX_INST_DATA_PATH_DECODE_RF_n4860, 
      DLX_INST_DATA_PATH_DECODE_RF_n4859, DLX_INST_DATA_PATH_DECODE_RF_n4858, 
      DLX_INST_DATA_PATH_DECODE_RF_n4857, DLX_INST_DATA_PATH_DECODE_RF_n4856, 
      DLX_INST_DATA_PATH_DECODE_RF_n4855, DLX_INST_DATA_PATH_DECODE_RF_n4854, 
      DLX_INST_DATA_PATH_DECODE_RF_n4853, DLX_INST_DATA_PATH_DECODE_RF_n4852, 
      DLX_INST_DATA_PATH_DECODE_RF_n4851, DLX_INST_DATA_PATH_DECODE_RF_n4850, 
      DLX_INST_DATA_PATH_DECODE_RF_n4849, DLX_INST_DATA_PATH_DECODE_RF_n4848, 
      DLX_INST_DATA_PATH_DECODE_RF_n4847, DLX_INST_DATA_PATH_DECODE_RF_n4846, 
      DLX_INST_DATA_PATH_DECODE_RF_n4845, DLX_INST_DATA_PATH_DECODE_RF_n4844, 
      DLX_INST_DATA_PATH_DECODE_RF_n4843, DLX_INST_DATA_PATH_DECODE_RF_n4842, 
      DLX_INST_DATA_PATH_DECODE_RF_n4841, DLX_INST_DATA_PATH_DECODE_RF_n4840, 
      DLX_INST_DATA_PATH_DECODE_RF_n4839, DLX_INST_DATA_PATH_DECODE_RF_n4838, 
      DLX_INST_DATA_PATH_DECODE_RF_n4837, DLX_INST_DATA_PATH_DECODE_RF_n4836, 
      DLX_INST_DATA_PATH_DECODE_RF_n4835, DLX_INST_DATA_PATH_DECODE_RF_n4834, 
      DLX_INST_DATA_PATH_DECODE_RF_n4833, DLX_INST_DATA_PATH_DECODE_RF_n4832, 
      DLX_INST_DATA_PATH_DECODE_RF_n4831, DLX_INST_DATA_PATH_DECODE_RF_n4830, 
      DLX_INST_DATA_PATH_DECODE_RF_n4829, DLX_INST_DATA_PATH_DECODE_RF_n4828, 
      DLX_INST_DATA_PATH_DECODE_RF_n4827, DLX_INST_DATA_PATH_DECODE_RF_n4826, 
      DLX_INST_DATA_PATH_DECODE_RF_n4825, DLX_INST_DATA_PATH_DECODE_RF_n4824, 
      DLX_INST_DATA_PATH_DECODE_RF_n4823, DLX_INST_DATA_PATH_DECODE_RF_n4822, 
      DLX_INST_DATA_PATH_DECODE_RF_n4821, DLX_INST_DATA_PATH_DECODE_RF_n4820, 
      DLX_INST_DATA_PATH_DECODE_RF_n4819, DLX_INST_DATA_PATH_DECODE_RF_n4818, 
      DLX_INST_DATA_PATH_DECODE_RF_n4817, DLX_INST_DATA_PATH_DECODE_RF_n4816, 
      DLX_INST_DATA_PATH_DECODE_RF_n4815, DLX_INST_DATA_PATH_DECODE_RF_n4814, 
      DLX_INST_DATA_PATH_DECODE_RF_n4813, DLX_INST_DATA_PATH_DECODE_RF_n4812, 
      DLX_INST_DATA_PATH_DECODE_RF_n4811, DLX_INST_DATA_PATH_DECODE_RF_n4810, 
      DLX_INST_DATA_PATH_DECODE_RF_n4809, DLX_INST_DATA_PATH_DECODE_RF_n4808, 
      DLX_INST_DATA_PATH_DECODE_RF_n4807, DLX_INST_DATA_PATH_DECODE_RF_n4806, 
      DLX_INST_DATA_PATH_DECODE_RF_n4805, DLX_INST_DATA_PATH_DECODE_RF_n4804, 
      DLX_INST_DATA_PATH_DECODE_RF_n4803, DLX_INST_DATA_PATH_DECODE_RF_n4802, 
      DLX_INST_DATA_PATH_DECODE_RF_n4801, DLX_INST_DATA_PATH_DECODE_RF_n4800, 
      DLX_INST_DATA_PATH_DECODE_RF_n4799, DLX_INST_DATA_PATH_DECODE_RF_n4798, 
      DLX_INST_DATA_PATH_DECODE_RF_n4797, DLX_INST_DATA_PATH_DECODE_RF_n4796, 
      DLX_INST_DATA_PATH_DECODE_RF_n4795, DLX_INST_DATA_PATH_DECODE_RF_n4794, 
      DLX_INST_DATA_PATH_DECODE_RF_n4793, DLX_INST_DATA_PATH_DECODE_RF_n4792, 
      DLX_INST_DATA_PATH_DECODE_RF_n4791, DLX_INST_DATA_PATH_DECODE_RF_n4790, 
      DLX_INST_DATA_PATH_DECODE_RF_n4789, DLX_INST_DATA_PATH_DECODE_RF_n4788, 
      DLX_INST_DATA_PATH_DECODE_RF_n4787, DLX_INST_DATA_PATH_DECODE_RF_n4786, 
      DLX_INST_DATA_PATH_DECODE_RF_n4785, DLX_INST_DATA_PATH_DECODE_RF_n4784, 
      DLX_INST_DATA_PATH_DECODE_RF_n4783, DLX_INST_DATA_PATH_DECODE_RF_n4782, 
      DLX_INST_DATA_PATH_DECODE_RF_n4781, DLX_INST_DATA_PATH_DECODE_RF_n4780, 
      DLX_INST_DATA_PATH_DECODE_RF_n4779, DLX_INST_DATA_PATH_DECODE_RF_n4778, 
      DLX_INST_DATA_PATH_DECODE_RF_n4777, DLX_INST_DATA_PATH_DECODE_RF_n4776, 
      DLX_INST_DATA_PATH_DECODE_RF_n4775, DLX_INST_DATA_PATH_DECODE_RF_n4774, 
      DLX_INST_DATA_PATH_DECODE_RF_n4773, DLX_INST_DATA_PATH_DECODE_RF_n4772, 
      DLX_INST_DATA_PATH_DECODE_RF_n4771, DLX_INST_DATA_PATH_DECODE_RF_n4770, 
      DLX_INST_DATA_PATH_DECODE_RF_n4769, DLX_INST_DATA_PATH_DECODE_RF_n4768, 
      DLX_INST_DATA_PATH_DECODE_RF_n4767, DLX_INST_DATA_PATH_DECODE_RF_n4766, 
      DLX_INST_DATA_PATH_DECODE_RF_n4765, DLX_INST_DATA_PATH_DECODE_RF_n4764, 
      DLX_INST_DATA_PATH_DECODE_RF_n4763, DLX_INST_DATA_PATH_DECODE_RF_n4762, 
      DLX_INST_DATA_PATH_DECODE_RF_n4761, DLX_INST_DATA_PATH_DECODE_RF_n4760, 
      DLX_INST_DATA_PATH_DECODE_RF_n4759, DLX_INST_DATA_PATH_DECODE_RF_n4758, 
      DLX_INST_DATA_PATH_DECODE_RF_n4757, DLX_INST_DATA_PATH_DECODE_RF_n4756, 
      DLX_INST_DATA_PATH_DECODE_RF_n4755, DLX_INST_DATA_PATH_DECODE_RF_n4754, 
      DLX_INST_DATA_PATH_DECODE_RF_n4753, DLX_INST_DATA_PATH_DECODE_RF_n4752, 
      DLX_INST_DATA_PATH_DECODE_RF_n4751, DLX_INST_DATA_PATH_DECODE_RF_n4750, 
      DLX_INST_DATA_PATH_DECODE_RF_n4749, DLX_INST_DATA_PATH_DECODE_RF_n4748, 
      DLX_INST_DATA_PATH_DECODE_RF_n4747, DLX_INST_DATA_PATH_DECODE_RF_n4746, 
      DLX_INST_DATA_PATH_DECODE_RF_n4745, DLX_INST_DATA_PATH_DECODE_RF_n4744, 
      DLX_INST_DATA_PATH_DECODE_RF_n4743, DLX_INST_DATA_PATH_DECODE_RF_n4742, 
      DLX_INST_DATA_PATH_DECODE_RF_n4741, DLX_INST_DATA_PATH_DECODE_RF_n4740, 
      DLX_INST_DATA_PATH_DECODE_RF_n4739, DLX_INST_DATA_PATH_DECODE_RF_n4738, 
      DLX_INST_DATA_PATH_DECODE_RF_n4737, DLX_INST_DATA_PATH_DECODE_RF_n4736, 
      DLX_INST_DATA_PATH_DECODE_RF_n4735, DLX_INST_DATA_PATH_DECODE_RF_n4734, 
      DLX_INST_DATA_PATH_DECODE_RF_n4733, DLX_INST_DATA_PATH_DECODE_RF_n4732, 
      DLX_INST_DATA_PATH_DECODE_RF_n4731, DLX_INST_DATA_PATH_DECODE_RF_n4730, 
      DLX_INST_DATA_PATH_DECODE_RF_n4729, DLX_INST_DATA_PATH_DECODE_RF_n4728, 
      DLX_INST_DATA_PATH_DECODE_RF_n4727, DLX_INST_DATA_PATH_DECODE_RF_n4726, 
      DLX_INST_DATA_PATH_DECODE_RF_n4725, DLX_INST_DATA_PATH_DECODE_RF_n4724, 
      DLX_INST_DATA_PATH_DECODE_RF_n4723, DLX_INST_DATA_PATH_DECODE_RF_n4722, 
      DLX_INST_DATA_PATH_DECODE_RF_n4721, DLX_INST_DATA_PATH_DECODE_RF_n4720, 
      DLX_INST_DATA_PATH_DECODE_RF_n4719, DLX_INST_DATA_PATH_DECODE_RF_n4718, 
      DLX_INST_DATA_PATH_DECODE_RF_n4717, DLX_INST_DATA_PATH_DECODE_RF_n4716, 
      DLX_INST_DATA_PATH_DECODE_RF_n4715, DLX_INST_DATA_PATH_DECODE_RF_n4714, 
      DLX_INST_DATA_PATH_DECODE_RF_n4713, DLX_INST_DATA_PATH_DECODE_RF_n4712, 
      DLX_INST_DATA_PATH_DECODE_RF_n4711, DLX_INST_DATA_PATH_DECODE_RF_n4710, 
      DLX_INST_DATA_PATH_DECODE_RF_n4709, DLX_INST_DATA_PATH_DECODE_RF_n4708, 
      DLX_INST_DATA_PATH_DECODE_RF_n4707, DLX_INST_DATA_PATH_DECODE_RF_n4706, 
      DLX_INST_DATA_PATH_DECODE_RF_n4705, DLX_INST_DATA_PATH_DECODE_RF_n4704, 
      DLX_INST_DATA_PATH_DECODE_RF_n4703, DLX_INST_DATA_PATH_DECODE_RF_n4702, 
      DLX_INST_DATA_PATH_DECODE_RF_n4701, DLX_INST_DATA_PATH_DECODE_RF_n4700, 
      DLX_INST_DATA_PATH_DECODE_RF_n4699, DLX_INST_DATA_PATH_DECODE_RF_n4698, 
      DLX_INST_DATA_PATH_DECODE_RF_n4697, DLX_INST_DATA_PATH_DECODE_RF_n4696, 
      DLX_INST_DATA_PATH_DECODE_RF_n4695, DLX_INST_DATA_PATH_DECODE_RF_n4694, 
      DLX_INST_DATA_PATH_DECODE_RF_n4693, DLX_INST_DATA_PATH_DECODE_RF_n4692, 
      DLX_INST_DATA_PATH_DECODE_RF_n4691, DLX_INST_DATA_PATH_DECODE_RF_n4690, 
      DLX_INST_DATA_PATH_DECODE_RF_n4689, DLX_INST_DATA_PATH_DECODE_RF_n4688, 
      DLX_INST_DATA_PATH_DECODE_RF_n4687, DLX_INST_DATA_PATH_DECODE_RF_n4686, 
      DLX_INST_DATA_PATH_DECODE_RF_n4685, DLX_INST_DATA_PATH_DECODE_RF_n4684, 
      DLX_INST_DATA_PATH_DECODE_RF_n4683, DLX_INST_DATA_PATH_DECODE_RF_n4682, 
      DLX_INST_DATA_PATH_DECODE_RF_n4681, DLX_INST_DATA_PATH_DECODE_RF_n4680, 
      DLX_INST_DATA_PATH_DECODE_RF_n4679, DLX_INST_DATA_PATH_DECODE_RF_n4678, 
      DLX_INST_DATA_PATH_DECODE_RF_n4677, DLX_INST_DATA_PATH_DECODE_RF_n4676, 
      DLX_INST_DATA_PATH_DECODE_RF_n4675, DLX_INST_DATA_PATH_DECODE_RF_n4674, 
      DLX_INST_DATA_PATH_DECODE_RF_n4673, DLX_INST_DATA_PATH_DECODE_RF_n4672, 
      DLX_INST_DATA_PATH_DECODE_RF_n4671, DLX_INST_DATA_PATH_DECODE_RF_n4670, 
      DLX_INST_DATA_PATH_DECODE_RF_n4669, DLX_INST_DATA_PATH_DECODE_RF_n4668, 
      DLX_INST_DATA_PATH_DECODE_RF_n4667, DLX_INST_DATA_PATH_DECODE_RF_n4666, 
      DLX_INST_DATA_PATH_DECODE_RF_n4665, DLX_INST_DATA_PATH_DECODE_RF_n4664, 
      DLX_INST_DATA_PATH_DECODE_RF_n4663, DLX_INST_DATA_PATH_DECODE_RF_n4662, 
      DLX_INST_DATA_PATH_DECODE_RF_n4661, DLX_INST_DATA_PATH_DECODE_RF_n4660, 
      DLX_INST_DATA_PATH_DECODE_RF_n4659, DLX_INST_DATA_PATH_DECODE_RF_n4658, 
      DLX_INST_DATA_PATH_DECODE_RF_n4657, DLX_INST_DATA_PATH_DECODE_RF_n4656, 
      DLX_INST_DATA_PATH_DECODE_RF_n4655, DLX_INST_DATA_PATH_DECODE_RF_n4654, 
      DLX_INST_DATA_PATH_DECODE_RF_n4653, DLX_INST_DATA_PATH_DECODE_RF_n4652, 
      DLX_INST_DATA_PATH_DECODE_RF_n4651, DLX_INST_DATA_PATH_DECODE_RF_n4650, 
      DLX_INST_DATA_PATH_DECODE_RF_n4649, DLX_INST_DATA_PATH_DECODE_RF_n4648, 
      DLX_INST_DATA_PATH_DECODE_RF_n4647, DLX_INST_DATA_PATH_DECODE_RF_n4646, 
      DLX_INST_DATA_PATH_DECODE_RF_n4645, DLX_INST_DATA_PATH_DECODE_RF_n4644, 
      DLX_INST_DATA_PATH_DECODE_RF_n4643, DLX_INST_DATA_PATH_DECODE_RF_n4642, 
      DLX_INST_DATA_PATH_DECODE_RF_n4641, DLX_INST_DATA_PATH_DECODE_RF_n4640, 
      DLX_INST_DATA_PATH_DECODE_RF_n4639, DLX_INST_DATA_PATH_DECODE_RF_n4638, 
      DLX_INST_DATA_PATH_DECODE_RF_n4637, DLX_INST_DATA_PATH_DECODE_RF_n4636, 
      DLX_INST_DATA_PATH_DECODE_RF_n4635, DLX_INST_DATA_PATH_DECODE_RF_n4634, 
      DLX_INST_DATA_PATH_DECODE_RF_n4633, DLX_INST_DATA_PATH_DECODE_RF_n4632, 
      DLX_INST_DATA_PATH_DECODE_RF_n4631, DLX_INST_DATA_PATH_DECODE_RF_n4630, 
      DLX_INST_DATA_PATH_DECODE_RF_n4629, DLX_INST_DATA_PATH_DECODE_RF_n4628, 
      DLX_INST_DATA_PATH_DECODE_RF_n4627, DLX_INST_DATA_PATH_DECODE_RF_n4626, 
      DLX_INST_DATA_PATH_DECODE_RF_n4625, DLX_INST_DATA_PATH_DECODE_RF_n4624, 
      DLX_INST_DATA_PATH_DECODE_RF_n4623, DLX_INST_DATA_PATH_DECODE_RF_n4622, 
      DLX_INST_DATA_PATH_DECODE_RF_n4621, DLX_INST_DATA_PATH_DECODE_RF_n4620, 
      DLX_INST_DATA_PATH_DECODE_RF_n4619, DLX_INST_DATA_PATH_DECODE_RF_n4618, 
      DLX_INST_DATA_PATH_DECODE_RF_n4617, DLX_INST_DATA_PATH_DECODE_RF_n4616, 
      DLX_INST_DATA_PATH_DECODE_RF_n4615, DLX_INST_DATA_PATH_DECODE_RF_n4614, 
      DLX_INST_DATA_PATH_DECODE_RF_n4613, DLX_INST_DATA_PATH_DECODE_RF_n4612, 
      DLX_INST_DATA_PATH_DECODE_RF_n4611, DLX_INST_DATA_PATH_DECODE_RF_n4610, 
      DLX_INST_DATA_PATH_DECODE_RF_n4609, DLX_INST_DATA_PATH_DECODE_RF_n4608, 
      DLX_INST_DATA_PATH_DECODE_RF_n4607, DLX_INST_DATA_PATH_DECODE_RF_n4606, 
      DLX_INST_DATA_PATH_DECODE_RF_n4605, DLX_INST_DATA_PATH_DECODE_RF_n4604, 
      DLX_INST_DATA_PATH_DECODE_RF_n4603, DLX_INST_DATA_PATH_DECODE_RF_n4602, 
      DLX_INST_DATA_PATH_DECODE_RF_n4601, DLX_INST_DATA_PATH_DECODE_RF_n4600, 
      DLX_INST_DATA_PATH_DECODE_RF_n4599, DLX_INST_DATA_PATH_DECODE_RF_n4598, 
      DLX_INST_DATA_PATH_DECODE_RF_n4597, DLX_INST_DATA_PATH_DECODE_RF_n4596, 
      DLX_INST_DATA_PATH_DECODE_RF_n4595, DLX_INST_DATA_PATH_DECODE_RF_n4594, 
      DLX_INST_DATA_PATH_DECODE_RF_n4593, DLX_INST_DATA_PATH_DECODE_RF_n4592, 
      DLX_INST_DATA_PATH_DECODE_RF_n4591, DLX_INST_DATA_PATH_DECODE_RF_n4590, 
      DLX_INST_DATA_PATH_DECODE_RF_n4589, DLX_INST_DATA_PATH_DECODE_RF_n4588, 
      DLX_INST_DATA_PATH_DECODE_RF_n4587, DLX_INST_DATA_PATH_DECODE_RF_n4586, 
      DLX_INST_DATA_PATH_DECODE_RF_n4585, DLX_INST_DATA_PATH_DECODE_RF_n4584, 
      DLX_INST_DATA_PATH_DECODE_RF_n4583, DLX_INST_DATA_PATH_DECODE_RF_n4582, 
      DLX_INST_DATA_PATH_DECODE_RF_n4581, DLX_INST_DATA_PATH_DECODE_RF_n4580, 
      DLX_INST_DATA_PATH_DECODE_RF_n4579, DLX_INST_DATA_PATH_DECODE_RF_n4578, 
      DLX_INST_DATA_PATH_DECODE_RF_n4577, DLX_INST_DATA_PATH_DECODE_RF_n4576, 
      DLX_INST_DATA_PATH_DECODE_RF_n4575, DLX_INST_DATA_PATH_DECODE_RF_n4574, 
      DLX_INST_DATA_PATH_DECODE_RF_n4573, DLX_INST_DATA_PATH_DECODE_RF_n4572, 
      DLX_INST_DATA_PATH_DECODE_RF_n4571, DLX_INST_DATA_PATH_DECODE_RF_n4570, 
      DLX_INST_DATA_PATH_DECODE_RF_n4569, DLX_INST_DATA_PATH_DECODE_RF_n4568, 
      DLX_INST_DATA_PATH_DECODE_RF_n4567, DLX_INST_DATA_PATH_DECODE_RF_n4566, 
      DLX_INST_DATA_PATH_DECODE_RF_n4565, DLX_INST_DATA_PATH_DECODE_RF_n4564, 
      DLX_INST_DATA_PATH_DECODE_RF_n4563, DLX_INST_DATA_PATH_DECODE_RF_n4562, 
      DLX_INST_DATA_PATH_DECODE_RF_n4561, DLX_INST_DATA_PATH_DECODE_RF_n4560, 
      DLX_INST_DATA_PATH_DECODE_RF_n4559, DLX_INST_DATA_PATH_DECODE_RF_n4558, 
      DLX_INST_DATA_PATH_DECODE_RF_n4557, DLX_INST_DATA_PATH_DECODE_RF_n4556, 
      DLX_INST_DATA_PATH_DECODE_RF_n4555, DLX_INST_DATA_PATH_DECODE_RF_n4554, 
      DLX_INST_DATA_PATH_DECODE_RF_n4553, DLX_INST_DATA_PATH_DECODE_RF_n4552, 
      DLX_INST_DATA_PATH_DECODE_RF_n4551, DLX_INST_DATA_PATH_DECODE_RF_n4550, 
      DLX_INST_DATA_PATH_DECODE_RF_n4549, DLX_INST_DATA_PATH_DECODE_RF_n4548, 
      DLX_INST_DATA_PATH_DECODE_RF_n4547, DLX_INST_DATA_PATH_DECODE_RF_n4546, 
      DLX_INST_DATA_PATH_DECODE_RF_n4545, DLX_INST_DATA_PATH_DECODE_RF_n4544, 
      DLX_INST_DATA_PATH_DECODE_RF_n4543, DLX_INST_DATA_PATH_DECODE_RF_n4542, 
      DLX_INST_DATA_PATH_DECODE_RF_n4541, DLX_INST_DATA_PATH_DECODE_RF_n4540, 
      DLX_INST_DATA_PATH_DECODE_RF_n4539, DLX_INST_DATA_PATH_DECODE_RF_n4538, 
      DLX_INST_DATA_PATH_DECODE_RF_n4537, DLX_INST_DATA_PATH_DECODE_RF_n4536, 
      DLX_INST_DATA_PATH_DECODE_RF_n4535, DLX_INST_DATA_PATH_DECODE_RF_n4534, 
      DLX_INST_DATA_PATH_DECODE_RF_n4533, DLX_INST_DATA_PATH_DECODE_RF_n4532, 
      DLX_INST_DATA_PATH_DECODE_RF_n4531, DLX_INST_DATA_PATH_DECODE_RF_n4530, 
      DLX_INST_DATA_PATH_DECODE_RF_n4529, DLX_INST_DATA_PATH_DECODE_RF_n4528, 
      DLX_INST_DATA_PATH_DECODE_RF_n4527, DLX_INST_DATA_PATH_DECODE_RF_n4526, 
      DLX_INST_DATA_PATH_DECODE_RF_n4525, DLX_INST_DATA_PATH_DECODE_RF_n4524, 
      DLX_INST_DATA_PATH_DECODE_RF_n4523, DLX_INST_DATA_PATH_DECODE_RF_n4522, 
      DLX_INST_DATA_PATH_DECODE_RF_n4521, DLX_INST_DATA_PATH_DECODE_RF_n4520, 
      DLX_INST_DATA_PATH_DECODE_RF_n4519, DLX_INST_DATA_PATH_DECODE_RF_n4518, 
      DLX_INST_DATA_PATH_DECODE_RF_n4517, DLX_INST_DATA_PATH_DECODE_RF_n4516, 
      DLX_INST_DATA_PATH_DECODE_RF_n4515, DLX_INST_DATA_PATH_DECODE_RF_n4514, 
      DLX_INST_DATA_PATH_DECODE_RF_n4513, DLX_INST_DATA_PATH_DECODE_RF_n4512, 
      DLX_INST_DATA_PATH_DECODE_RF_n4511, DLX_INST_DATA_PATH_DECODE_RF_n4510, 
      DLX_INST_DATA_PATH_DECODE_RF_n4509, DLX_INST_DATA_PATH_DECODE_RF_n4508, 
      DLX_INST_DATA_PATH_DECODE_RF_n4507, DLX_INST_DATA_PATH_DECODE_RF_n4506, 
      DLX_INST_DATA_PATH_DECODE_RF_n4505, DLX_INST_DATA_PATH_DECODE_RF_n4504, 
      DLX_INST_DATA_PATH_DECODE_RF_n4503, DLX_INST_DATA_PATH_DECODE_RF_n4502, 
      DLX_INST_DATA_PATH_DECODE_RF_n4501, DLX_INST_DATA_PATH_DECODE_RF_n4500, 
      DLX_INST_DATA_PATH_DECODE_RF_n4499, DLX_INST_DATA_PATH_DECODE_RF_n4498, 
      DLX_INST_DATA_PATH_DECODE_RF_n4497, DLX_INST_DATA_PATH_DECODE_RF_n4496, 
      DLX_INST_DATA_PATH_DECODE_RF_n4495, DLX_INST_DATA_PATH_DECODE_RF_n4494, 
      DLX_INST_DATA_PATH_DECODE_RF_n4493, DLX_INST_DATA_PATH_DECODE_RF_n4492, 
      DLX_INST_DATA_PATH_DECODE_RF_n4491, DLX_INST_DATA_PATH_DECODE_RF_n4490, 
      DLX_INST_DATA_PATH_DECODE_RF_n4489, DLX_INST_DATA_PATH_DECODE_RF_n4488, 
      DLX_INST_DATA_PATH_DECODE_RF_n4487, DLX_INST_DATA_PATH_DECODE_RF_n4486, 
      DLX_INST_DATA_PATH_DECODE_RF_n4485, DLX_INST_DATA_PATH_DECODE_RF_n4484, 
      DLX_INST_DATA_PATH_DECODE_RF_n4483, DLX_INST_DATA_PATH_DECODE_RF_n4482, 
      DLX_INST_DATA_PATH_DECODE_RF_n4481, DLX_INST_DATA_PATH_DECODE_RF_n4480, 
      DLX_INST_DATA_PATH_DECODE_RF_n4479, DLX_INST_DATA_PATH_DECODE_RF_n4478, 
      DLX_INST_DATA_PATH_DECODE_RF_n4477, DLX_INST_DATA_PATH_DECODE_RF_n4476, 
      DLX_INST_DATA_PATH_DECODE_RF_n4475, DLX_INST_DATA_PATH_DECODE_RF_n4474, 
      DLX_INST_DATA_PATH_DECODE_RF_n4473, DLX_INST_DATA_PATH_DECODE_RF_n4472, 
      DLX_INST_DATA_PATH_DECODE_RF_n4471, DLX_INST_DATA_PATH_DECODE_RF_n4470, 
      DLX_INST_DATA_PATH_DECODE_RF_n4469, DLX_INST_DATA_PATH_DECODE_RF_n4468, 
      DLX_INST_DATA_PATH_DECODE_RF_n4467, DLX_INST_DATA_PATH_DECODE_RF_n4466, 
      DLX_INST_DATA_PATH_DECODE_RF_n4465, DLX_INST_DATA_PATH_DECODE_RF_n4464, 
      DLX_INST_DATA_PATH_DECODE_RF_n4463, DLX_INST_DATA_PATH_DECODE_RF_n4462, 
      DLX_INST_DATA_PATH_DECODE_RF_n4461, DLX_INST_DATA_PATH_DECODE_RF_n4460, 
      DLX_INST_DATA_PATH_DECODE_RF_n4459, DLX_INST_DATA_PATH_DECODE_RF_n4458, 
      DLX_INST_DATA_PATH_DECODE_RF_n4457, DLX_INST_DATA_PATH_DECODE_RF_n4456, 
      DLX_INST_DATA_PATH_DECODE_RF_n4455, DLX_INST_DATA_PATH_DECODE_RF_n4454, 
      DLX_INST_DATA_PATH_DECODE_RF_n4453, DLX_INST_DATA_PATH_DECODE_RF_n4452, 
      DLX_INST_DATA_PATH_DECODE_RF_n4451, DLX_INST_DATA_PATH_DECODE_RF_n4450, 
      DLX_INST_DATA_PATH_DECODE_RF_n4449, DLX_INST_DATA_PATH_DECODE_RF_n4448, 
      DLX_INST_DATA_PATH_DECODE_RF_n4447, DLX_INST_DATA_PATH_DECODE_RF_n4446, 
      DLX_INST_DATA_PATH_DECODE_RF_n4445, DLX_INST_DATA_PATH_DECODE_RF_n4444, 
      DLX_INST_DATA_PATH_DECODE_RF_n4443, DLX_INST_DATA_PATH_DECODE_RF_n4442, 
      DLX_INST_DATA_PATH_DECODE_RF_n4441, DLX_INST_DATA_PATH_DECODE_RF_n4440, 
      DLX_INST_DATA_PATH_DECODE_RF_n4439, DLX_INST_DATA_PATH_DECODE_RF_n4438, 
      DLX_INST_DATA_PATH_DECODE_RF_n4437, DLX_INST_DATA_PATH_DECODE_RF_n4436, 
      DLX_INST_DATA_PATH_DECODE_RF_n4435, DLX_INST_DATA_PATH_DECODE_RF_n4434, 
      DLX_INST_DATA_PATH_DECODE_RF_n4433, DLX_INST_DATA_PATH_DECODE_RF_n4432, 
      DLX_INST_DATA_PATH_DECODE_RF_n4431, DLX_INST_DATA_PATH_DECODE_RF_n4430, 
      DLX_INST_DATA_PATH_DECODE_RF_n4429, DLX_INST_DATA_PATH_DECODE_RF_n4428, 
      DLX_INST_DATA_PATH_DECODE_RF_n4427, DLX_INST_DATA_PATH_DECODE_RF_n4426, 
      DLX_INST_DATA_PATH_DECODE_RF_n4425, DLX_INST_DATA_PATH_DECODE_RF_n4424, 
      DLX_INST_DATA_PATH_DECODE_RF_n4423, DLX_INST_DATA_PATH_DECODE_RF_n4422, 
      DLX_INST_DATA_PATH_DECODE_RF_n4421, DLX_INST_DATA_PATH_DECODE_RF_n4420, 
      DLX_INST_DATA_PATH_DECODE_RF_n4419, DLX_INST_DATA_PATH_DECODE_RF_n4418, 
      DLX_INST_DATA_PATH_DECODE_RF_n4417, DLX_INST_DATA_PATH_DECODE_RF_n4416, 
      DLX_INST_DATA_PATH_DECODE_RF_n4415, DLX_INST_DATA_PATH_DECODE_RF_n4414, 
      DLX_INST_DATA_PATH_DECODE_RF_n4413, DLX_INST_DATA_PATH_DECODE_RF_n4412, 
      DLX_INST_DATA_PATH_DECODE_RF_n4411, DLX_INST_DATA_PATH_DECODE_RF_n4410, 
      DLX_INST_DATA_PATH_DECODE_RF_n4409, DLX_INST_DATA_PATH_DECODE_RF_n4408, 
      DLX_INST_DATA_PATH_DECODE_RF_n4407, DLX_INST_DATA_PATH_DECODE_RF_n4406, 
      DLX_INST_DATA_PATH_DECODE_RF_n4405, DLX_INST_DATA_PATH_DECODE_RF_n4404, 
      DLX_INST_DATA_PATH_DECODE_RF_n4403, DLX_INST_DATA_PATH_DECODE_RF_n4402, 
      DLX_INST_DATA_PATH_DECODE_RF_n4401, DLX_INST_DATA_PATH_DECODE_RF_n4400, 
      DLX_INST_DATA_PATH_DECODE_RF_n4399, DLX_INST_DATA_PATH_DECODE_RF_n4398, 
      DLX_INST_DATA_PATH_DECODE_RF_n4397, DLX_INST_DATA_PATH_DECODE_RF_n4396, 
      DLX_INST_DATA_PATH_DECODE_RF_n4395, DLX_INST_DATA_PATH_DECODE_RF_n4394, 
      DLX_INST_DATA_PATH_DECODE_RF_n4393, DLX_INST_DATA_PATH_DECODE_RF_n4392, 
      DLX_INST_DATA_PATH_DECODE_RF_n4391, DLX_INST_DATA_PATH_DECODE_RF_n4390, 
      DLX_INST_DATA_PATH_DECODE_RF_n4389, DLX_INST_DATA_PATH_DECODE_RF_n4388, 
      DLX_INST_DATA_PATH_DECODE_RF_n4387, DLX_INST_DATA_PATH_DECODE_RF_n4386, 
      DLX_INST_DATA_PATH_DECODE_RF_n4385, DLX_INST_DATA_PATH_DECODE_RF_n4384, 
      DLX_INST_DATA_PATH_DECODE_RF_n4383, DLX_INST_DATA_PATH_DECODE_RF_n4382, 
      DLX_INST_DATA_PATH_DECODE_RF_n4381, DLX_INST_DATA_PATH_DECODE_RF_n4380, 
      DLX_INST_DATA_PATH_DECODE_RF_n4379, DLX_INST_DATA_PATH_DECODE_RF_n4378, 
      DLX_INST_DATA_PATH_DECODE_RF_n4377, DLX_INST_DATA_PATH_DECODE_RF_n4376, 
      DLX_INST_DATA_PATH_DECODE_RF_n4375, DLX_INST_DATA_PATH_DECODE_RF_n4374, 
      DLX_INST_DATA_PATH_DECODE_RF_n4373, DLX_INST_DATA_PATH_DECODE_RF_n4372, 
      DLX_INST_DATA_PATH_DECODE_RF_n4371, DLX_INST_DATA_PATH_DECODE_RF_n4370, 
      DLX_INST_DATA_PATH_DECODE_RF_n4369, DLX_INST_DATA_PATH_DECODE_RF_n4368, 
      DLX_INST_DATA_PATH_DECODE_RF_n4367, DLX_INST_DATA_PATH_DECODE_RF_n4366, 
      DLX_INST_DATA_PATH_DECODE_RF_n4365, DLX_INST_DATA_PATH_DECODE_RF_n4364, 
      DLX_INST_DATA_PATH_DECODE_RF_n4363, DLX_INST_DATA_PATH_DECODE_RF_n4362, 
      DLX_INST_DATA_PATH_DECODE_RF_n4361, DLX_INST_DATA_PATH_DECODE_RF_n4360, 
      DLX_INST_DATA_PATH_DECODE_RF_n4359, DLX_INST_DATA_PATH_DECODE_RF_n4358, 
      DLX_INST_DATA_PATH_DECODE_RF_n4357, DLX_INST_DATA_PATH_DECODE_RF_n4356, 
      DLX_INST_DATA_PATH_DECODE_RF_n4355, DLX_INST_DATA_PATH_DECODE_RF_n4354, 
      DLX_INST_DATA_PATH_DECODE_RF_n4353, DLX_INST_DATA_PATH_DECODE_RF_n4352, 
      DLX_INST_DATA_PATH_DECODE_RF_n4351, DLX_INST_DATA_PATH_DECODE_RF_n4350, 
      DLX_INST_DATA_PATH_DECODE_RF_n4349, DLX_INST_DATA_PATH_DECODE_RF_n4348, 
      DLX_INST_DATA_PATH_DECODE_RF_n4347, DLX_INST_DATA_PATH_DECODE_RF_n4346, 
      DLX_INST_DATA_PATH_DECODE_RF_n4345, DLX_INST_DATA_PATH_DECODE_RF_n4344, 
      DLX_INST_DATA_PATH_DECODE_RF_n4343, DLX_INST_DATA_PATH_DECODE_RF_n4342, 
      DLX_INST_DATA_PATH_DECODE_RF_n4341, DLX_INST_DATA_PATH_DECODE_RF_n4340, 
      DLX_INST_DATA_PATH_DECODE_RF_n4339, DLX_INST_DATA_PATH_DECODE_RF_n4338, 
      DLX_INST_DATA_PATH_DECODE_RF_n4337, DLX_INST_DATA_PATH_DECODE_RF_n4336, 
      DLX_INST_DATA_PATH_DECODE_RF_n4335, DLX_INST_DATA_PATH_DECODE_RF_n4334, 
      DLX_INST_DATA_PATH_DECODE_RF_n4333, DLX_INST_DATA_PATH_DECODE_RF_n4332, 
      DLX_INST_DATA_PATH_DECODE_RF_n4331, DLX_INST_DATA_PATH_DECODE_RF_n4330, 
      DLX_INST_DATA_PATH_DECODE_RF_n4329, DLX_INST_DATA_PATH_DECODE_RF_n4328, 
      DLX_INST_DATA_PATH_DECODE_RF_n4327, DLX_INST_DATA_PATH_DECODE_RF_n4326, 
      DLX_INST_DATA_PATH_DECODE_RF_n4325, DLX_INST_DATA_PATH_DECODE_RF_n4324, 
      DLX_INST_DATA_PATH_DECODE_RF_n4323, DLX_INST_DATA_PATH_DECODE_RF_n4322, 
      DLX_INST_DATA_PATH_DECODE_RF_n4321, DLX_INST_DATA_PATH_DECODE_RF_n4320, 
      DLX_INST_DATA_PATH_DECODE_RF_n4319, DLX_INST_DATA_PATH_DECODE_RF_n4318, 
      DLX_INST_DATA_PATH_DECODE_RF_n4317, DLX_INST_DATA_PATH_DECODE_RF_n4316, 
      DLX_INST_DATA_PATH_DECODE_RF_n4315, DLX_INST_DATA_PATH_DECODE_RF_n4314, 
      DLX_INST_DATA_PATH_DECODE_RF_n4313, DLX_INST_DATA_PATH_DECODE_RF_n4312, 
      DLX_INST_DATA_PATH_DECODE_RF_n4311, DLX_INST_DATA_PATH_DECODE_RF_n4310, 
      DLX_INST_DATA_PATH_DECODE_RF_n4309, DLX_INST_DATA_PATH_DECODE_RF_n4308, 
      DLX_INST_DATA_PATH_DECODE_RF_n4307, DLX_INST_DATA_PATH_DECODE_RF_n4306, 
      DLX_INST_DATA_PATH_DECODE_RF_n4305, DLX_INST_DATA_PATH_DECODE_RF_n4304, 
      DLX_INST_DATA_PATH_DECODE_RF_n4303, DLX_INST_DATA_PATH_DECODE_RF_n4302, 
      DLX_INST_DATA_PATH_DECODE_RF_n4301, DLX_INST_DATA_PATH_DECODE_RF_n4300, 
      DLX_INST_DATA_PATH_DECODE_RF_n4299, DLX_INST_DATA_PATH_DECODE_RF_n4298, 
      DLX_INST_DATA_PATH_DECODE_RF_n4297, DLX_INST_DATA_PATH_DECODE_RF_n4296, 
      DLX_INST_DATA_PATH_DECODE_RF_n4295, DLX_INST_DATA_PATH_DECODE_RF_n4294, 
      DLX_INST_DATA_PATH_DECODE_RF_n4293, DLX_INST_DATA_PATH_DECODE_RF_n4292, 
      DLX_INST_DATA_PATH_DECODE_RF_n4291, DLX_INST_DATA_PATH_DECODE_RF_n4290, 
      DLX_INST_DATA_PATH_DECODE_RF_n4289, DLX_INST_DATA_PATH_DECODE_RF_n4288, 
      DLX_INST_DATA_PATH_DECODE_RF_n4287, DLX_INST_DATA_PATH_DECODE_RF_n4286, 
      DLX_INST_DATA_PATH_DECODE_RF_n4285, DLX_INST_DATA_PATH_DECODE_RF_n4284, 
      DLX_INST_DATA_PATH_DECODE_RF_n4283, DLX_INST_DATA_PATH_DECODE_RF_n4282, 
      DLX_INST_DATA_PATH_DECODE_RF_n4281, DLX_INST_DATA_PATH_DECODE_RF_n4280, 
      DLX_INST_DATA_PATH_DECODE_RF_n4279, DLX_INST_DATA_PATH_DECODE_RF_n4278, 
      DLX_INST_DATA_PATH_DECODE_RF_n4277, DLX_INST_DATA_PATH_DECODE_RF_n4276, 
      DLX_INST_DATA_PATH_DECODE_RF_n4275, DLX_INST_DATA_PATH_DECODE_RF_n4274, 
      DLX_INST_DATA_PATH_DECODE_RF_n4273, DLX_INST_DATA_PATH_DECODE_RF_n4272, 
      DLX_INST_DATA_PATH_DECODE_RF_n4271, DLX_INST_DATA_PATH_DECODE_RF_n4270, 
      DLX_INST_DATA_PATH_DECODE_RF_n4269, DLX_INST_DATA_PATH_DECODE_RF_n4268, 
      DLX_INST_DATA_PATH_DECODE_RF_n4267, DLX_INST_DATA_PATH_DECODE_RF_n4266, 
      DLX_INST_DATA_PATH_DECODE_RF_n4265, DLX_INST_DATA_PATH_DECODE_RF_n4264, 
      DLX_INST_DATA_PATH_DECODE_RF_n4263, DLX_INST_DATA_PATH_DECODE_RF_n4262, 
      DLX_INST_DATA_PATH_DECODE_RF_n4261, DLX_INST_DATA_PATH_DECODE_RF_n4260, 
      DLX_INST_DATA_PATH_DECODE_RF_n4259, DLX_INST_DATA_PATH_DECODE_RF_n4258, 
      DLX_INST_DATA_PATH_DECODE_RF_n4257, DLX_INST_DATA_PATH_DECODE_RF_n4256, 
      DLX_INST_DATA_PATH_DECODE_RF_n4255, DLX_INST_DATA_PATH_DECODE_RF_n4254, 
      DLX_INST_DATA_PATH_DECODE_RF_n4253, DLX_INST_DATA_PATH_DECODE_RF_n4252, 
      DLX_INST_DATA_PATH_DECODE_RF_n4251, DLX_INST_DATA_PATH_DECODE_RF_n4250, 
      DLX_INST_DATA_PATH_DECODE_RF_n4249, DLX_INST_DATA_PATH_DECODE_RF_n4248, 
      DLX_INST_DATA_PATH_DECODE_RF_n4247, DLX_INST_DATA_PATH_DECODE_RF_n4246, 
      DLX_INST_DATA_PATH_DECODE_RF_n4245, DLX_INST_DATA_PATH_DECODE_RF_n4244, 
      DLX_INST_DATA_PATH_DECODE_RF_n4243, DLX_INST_DATA_PATH_DECODE_RF_n4242, 
      DLX_INST_DATA_PATH_DECODE_RF_n4241, DLX_INST_DATA_PATH_DECODE_RF_n4240, 
      DLX_INST_DATA_PATH_DECODE_RF_n4239, DLX_INST_DATA_PATH_DECODE_RF_n4238, 
      DLX_INST_DATA_PATH_DECODE_RF_n4237, DLX_INST_DATA_PATH_DECODE_RF_n4236, 
      DLX_INST_DATA_PATH_DECODE_RF_n4235, DLX_INST_DATA_PATH_DECODE_RF_n4234, 
      DLX_INST_DATA_PATH_DECODE_RF_n4233, DLX_INST_DATA_PATH_DECODE_RF_n4232, 
      DLX_INST_DATA_PATH_DECODE_RF_n4231, DLX_INST_DATA_PATH_DECODE_RF_n4230, 
      DLX_INST_DATA_PATH_DECODE_RF_n4229, DLX_INST_DATA_PATH_DECODE_RF_n4228, 
      DLX_INST_DATA_PATH_DECODE_RF_n4227, DLX_INST_DATA_PATH_DECODE_RF_n4226, 
      DLX_INST_DATA_PATH_DECODE_RF_n4225, DLX_INST_DATA_PATH_DECODE_RF_n4224, 
      DLX_INST_DATA_PATH_DECODE_RF_n4223, DLX_INST_DATA_PATH_DECODE_RF_n4222, 
      DLX_INST_DATA_PATH_DECODE_RF_n4221, DLX_INST_DATA_PATH_DECODE_RF_n4220, 
      DLX_INST_DATA_PATH_DECODE_RF_n4219, DLX_INST_DATA_PATH_DECODE_RF_n4218, 
      DLX_INST_DATA_PATH_DECODE_RF_n4217, DLX_INST_DATA_PATH_DECODE_RF_n4216, 
      DLX_INST_DATA_PATH_DECODE_RF_n4215, DLX_INST_DATA_PATH_DECODE_RF_n4214, 
      DLX_INST_DATA_PATH_DECODE_RF_n4213, DLX_INST_DATA_PATH_DECODE_RF_n4212, 
      DLX_INST_DATA_PATH_DECODE_RF_n4211, DLX_INST_DATA_PATH_DECODE_RF_n4210, 
      DLX_INST_DATA_PATH_DECODE_RF_n4209, DLX_INST_DATA_PATH_DECODE_RF_n4208, 
      DLX_INST_DATA_PATH_DECODE_RF_n4207, DLX_INST_DATA_PATH_DECODE_RF_n4206, 
      DLX_INST_DATA_PATH_DECODE_RF_n4205, DLX_INST_DATA_PATH_DECODE_RF_n4204, 
      DLX_INST_DATA_PATH_DECODE_RF_n4203, DLX_INST_DATA_PATH_DECODE_RF_n4202, 
      DLX_INST_DATA_PATH_DECODE_RF_n4201, DLX_INST_DATA_PATH_DECODE_RF_n4200, 
      DLX_INST_DATA_PATH_DECODE_RF_n4199, DLX_INST_DATA_PATH_DECODE_RF_n4198, 
      DLX_INST_DATA_PATH_DECODE_RF_n4197, DLX_INST_DATA_PATH_DECODE_RF_n4196, 
      DLX_INST_DATA_PATH_DECODE_RF_n4195, DLX_INST_DATA_PATH_DECODE_RF_n4194, 
      DLX_INST_DATA_PATH_DECODE_RF_n4193, DLX_INST_DATA_PATH_DECODE_RF_n4192, 
      DLX_INST_DATA_PATH_DECODE_RF_n4191, DLX_INST_DATA_PATH_DECODE_RF_n4190, 
      DLX_INST_DATA_PATH_DECODE_RF_n4189, DLX_INST_DATA_PATH_DECODE_RF_n4188, 
      DLX_INST_DATA_PATH_DECODE_RF_n4187, DLX_INST_DATA_PATH_DECODE_RF_n4186, 
      DLX_INST_DATA_PATH_DECODE_RF_n4185, DLX_INST_DATA_PATH_DECODE_RF_n4184, 
      DLX_INST_DATA_PATH_DECODE_RF_n4183, DLX_INST_DATA_PATH_DECODE_RF_n4182, 
      DLX_INST_DATA_PATH_DECODE_RF_n4181, DLX_INST_DATA_PATH_DECODE_RF_n4180, 
      DLX_INST_DATA_PATH_DECODE_RF_n4179, DLX_INST_DATA_PATH_DECODE_RF_n4178, 
      DLX_INST_DATA_PATH_DECODE_RF_n4177, DLX_INST_DATA_PATH_DECODE_RF_n4176, 
      DLX_INST_DATA_PATH_DECODE_RF_n4175, DLX_INST_DATA_PATH_DECODE_RF_n4174, 
      DLX_INST_DATA_PATH_DECODE_RF_n4173, DLX_INST_DATA_PATH_DECODE_RF_n4172, 
      DLX_INST_DATA_PATH_DECODE_RF_n4171, DLX_INST_DATA_PATH_DECODE_RF_n4170, 
      DLX_INST_DATA_PATH_DECODE_RF_n4169, DLX_INST_DATA_PATH_DECODE_RF_n4168, 
      DLX_INST_DATA_PATH_DECODE_RF_n4167, DLX_INST_DATA_PATH_DECODE_RF_n4166, 
      DLX_INST_DATA_PATH_DECODE_RF_n4165, DLX_INST_DATA_PATH_DECODE_RF_n4164, 
      DLX_INST_DATA_PATH_DECODE_RF_n4163, DLX_INST_DATA_PATH_DECODE_RF_n4162, 
      DLX_INST_DATA_PATH_DECODE_RF_n4161, DLX_INST_DATA_PATH_DECODE_RF_n4160, 
      DLX_INST_DATA_PATH_DECODE_RF_n4159, DLX_INST_DATA_PATH_DECODE_RF_n4158, 
      DLX_INST_DATA_PATH_DECODE_RF_n4157, DLX_INST_DATA_PATH_DECODE_RF_n4156, 
      DLX_INST_DATA_PATH_DECODE_RF_n4155, DLX_INST_DATA_PATH_DECODE_RF_n4154, 
      DLX_INST_DATA_PATH_DECODE_RF_n4153, DLX_INST_DATA_PATH_DECODE_RF_n4152, 
      DLX_INST_DATA_PATH_DECODE_RF_n4151, DLX_INST_DATA_PATH_DECODE_RF_n4150, 
      DLX_INST_DATA_PATH_DECODE_RF_n4149, DLX_INST_DATA_PATH_DECODE_RF_n4148, 
      DLX_INST_DATA_PATH_DECODE_RF_n4147, DLX_INST_DATA_PATH_DECODE_RF_n4146, 
      DLX_INST_DATA_PATH_DECODE_RF_n4145, DLX_INST_DATA_PATH_DECODE_RF_n4144, 
      DLX_INST_DATA_PATH_DECODE_RF_n4143, DLX_INST_DATA_PATH_DECODE_RF_n4142, 
      DLX_INST_DATA_PATH_DECODE_RF_n4141, DLX_INST_DATA_PATH_DECODE_RF_n4140, 
      DLX_INST_DATA_PATH_DECODE_RF_n4139, DLX_INST_DATA_PATH_DECODE_RF_n4138, 
      DLX_INST_DATA_PATH_DECODE_RF_n4137, DLX_INST_DATA_PATH_DECODE_RF_n4136, 
      DLX_INST_DATA_PATH_DECODE_RF_n4135, DLX_INST_DATA_PATH_DECODE_RF_n4134, 
      DLX_INST_DATA_PATH_DECODE_RF_n4133, DLX_INST_DATA_PATH_DECODE_RF_n4132, 
      DLX_INST_DATA_PATH_DECODE_RF_n4131, DLX_INST_DATA_PATH_DECODE_RF_n4130, 
      DLX_INST_DATA_PATH_DECODE_RF_n4129, DLX_INST_DATA_PATH_DECODE_RF_n4128, 
      DLX_INST_DATA_PATH_DECODE_RF_n4127, DLX_INST_DATA_PATH_DECODE_RF_n4126, 
      DLX_INST_DATA_PATH_DECODE_RF_n4125, DLX_INST_DATA_PATH_DECODE_RF_n4124, 
      DLX_INST_DATA_PATH_DECODE_RF_n4123, DLX_INST_DATA_PATH_DECODE_RF_n4122, 
      DLX_INST_DATA_PATH_DECODE_RF_n4121, DLX_INST_DATA_PATH_DECODE_RF_n4120, 
      DLX_INST_DATA_PATH_DECODE_RF_n4119, DLX_INST_DATA_PATH_DECODE_RF_n4118, 
      DLX_INST_DATA_PATH_DECODE_RF_n4117, DLX_INST_DATA_PATH_DECODE_RF_n4116, 
      DLX_INST_DATA_PATH_DECODE_RF_n4115, DLX_INST_DATA_PATH_DECODE_RF_n4114, 
      DLX_INST_DATA_PATH_DECODE_RF_n4113, DLX_INST_DATA_PATH_DECODE_RF_n4112, 
      DLX_INST_DATA_PATH_DECODE_RF_n4111, DLX_INST_DATA_PATH_DECODE_RF_n4110, 
      DLX_INST_DATA_PATH_DECODE_RF_n4109, DLX_INST_DATA_PATH_DECODE_RF_n4108, 
      DLX_INST_DATA_PATH_DECODE_RF_n4107, DLX_INST_DATA_PATH_DECODE_RF_n4106, 
      DLX_INST_DATA_PATH_DECODE_RF_n4105, DLX_INST_DATA_PATH_DECODE_RF_n4104, 
      DLX_INST_DATA_PATH_DECODE_RF_n4103, DLX_INST_DATA_PATH_DECODE_RF_n4102, 
      DLX_INST_DATA_PATH_DECODE_RF_n4101, DLX_INST_DATA_PATH_DECODE_RF_n4100, 
      DLX_INST_DATA_PATH_DECODE_RF_n4099, DLX_INST_DATA_PATH_DECODE_RF_n2326, 
      DLX_INST_DATA_PATH_DECODE_RF_n2325, DLX_INST_DATA_PATH_DECODE_RF_n2324, 
      DLX_INST_DATA_PATH_DECODE_RF_n2323, DLX_INST_DATA_PATH_DECODE_RF_n2322, 
      DLX_INST_DATA_PATH_DECODE_RF_n2321, DLX_INST_DATA_PATH_DECODE_RF_n2320, 
      DLX_INST_DATA_PATH_DECODE_RF_n2319, DLX_INST_DATA_PATH_DECODE_RF_n2318, 
      DLX_INST_DATA_PATH_DECODE_RF_n2317, DLX_INST_DATA_PATH_DECODE_RF_n2316, 
      DLX_INST_DATA_PATH_DECODE_RF_n2315, DLX_INST_DATA_PATH_DECODE_RF_n2314, 
      DLX_INST_DATA_PATH_DECODE_RF_n2313, DLX_INST_DATA_PATH_DECODE_RF_n2312, 
      DLX_INST_DATA_PATH_DECODE_RF_n2311, DLX_INST_DATA_PATH_DECODE_RF_n2310, 
      DLX_INST_DATA_PATH_DECODE_RF_n2309, DLX_INST_DATA_PATH_DECODE_RF_n2308, 
      DLX_INST_DATA_PATH_DECODE_RF_n2307, DLX_INST_DATA_PATH_DECODE_RF_n2306, 
      DLX_INST_DATA_PATH_DECODE_RF_n2305, DLX_INST_DATA_PATH_DECODE_RF_n2304, 
      DLX_INST_DATA_PATH_DECODE_RF_n2303, DLX_INST_DATA_PATH_DECODE_RF_n2302, 
      DLX_INST_DATA_PATH_DECODE_RF_n2301, DLX_INST_DATA_PATH_DECODE_RF_n2300, 
      DLX_INST_DATA_PATH_DECODE_RF_n2299, DLX_INST_DATA_PATH_DECODE_RF_n2298, 
      DLX_INST_DATA_PATH_DECODE_RF_n2297, DLX_INST_DATA_PATH_DECODE_RF_n2296, 
      DLX_INST_DATA_PATH_DECODE_RF_n2295, DLX_INST_DATA_PATH_DECODE_RF_n2294, 
      DLX_INST_DATA_PATH_DECODE_RF_n2293, DLX_INST_DATA_PATH_DECODE_RF_n2292, 
      DLX_INST_DATA_PATH_DECODE_RF_n2291, DLX_INST_DATA_PATH_DECODE_RF_n2290, 
      DLX_INST_DATA_PATH_DECODE_RF_n2289, DLX_INST_DATA_PATH_DECODE_RF_n2288, 
      DLX_INST_DATA_PATH_DECODE_RF_n2287, DLX_INST_DATA_PATH_DECODE_RF_n2286, 
      DLX_INST_DATA_PATH_DECODE_RF_n2285, DLX_INST_DATA_PATH_DECODE_RF_n2284, 
      DLX_INST_DATA_PATH_DECODE_RF_n2283, DLX_INST_DATA_PATH_DECODE_RF_n2282, 
      DLX_INST_DATA_PATH_DECODE_RF_n2281, DLX_INST_DATA_PATH_DECODE_RF_n2280, 
      DLX_INST_DATA_PATH_DECODE_RF_n2279, DLX_INST_DATA_PATH_DECODE_RF_n2278, 
      DLX_INST_DATA_PATH_DECODE_RF_n2277, DLX_INST_DATA_PATH_DECODE_RF_n2276, 
      DLX_INST_DATA_PATH_DECODE_RF_n2275, DLX_INST_DATA_PATH_DECODE_RF_n2274, 
      DLX_INST_DATA_PATH_DECODE_RF_n2273, DLX_INST_DATA_PATH_DECODE_RF_n2272, 
      DLX_INST_DATA_PATH_DECODE_RF_n2271, DLX_INST_DATA_PATH_DECODE_RF_n2270, 
      DLX_INST_DATA_PATH_DECODE_RF_n2269, DLX_INST_DATA_PATH_DECODE_RF_n2268, 
      DLX_INST_DATA_PATH_DECODE_RF_n2267, DLX_INST_DATA_PATH_DECODE_RF_n2266, 
      DLX_INST_DATA_PATH_DECODE_RF_n2265, DLX_INST_DATA_PATH_DECODE_RF_n2264, 
      DLX_INST_DATA_PATH_DECODE_RF_n2263, DLX_INST_DATA_PATH_DECODE_RF_n2262, 
      DLX_INST_DATA_PATH_DECODE_RF_n2261, DLX_INST_DATA_PATH_DECODE_RF_n2260, 
      DLX_INST_DATA_PATH_DECODE_RF_n2259, DLX_INST_DATA_PATH_DECODE_RF_n2258, 
      DLX_INST_DATA_PATH_DECODE_RF_n2257, DLX_INST_DATA_PATH_DECODE_RF_n2256, 
      DLX_INST_DATA_PATH_DECODE_RF_n2255, DLX_INST_DATA_PATH_DECODE_RF_n2254, 
      DLX_INST_DATA_PATH_DECODE_RF_n2253, DLX_INST_DATA_PATH_DECODE_RF_n2252, 
      DLX_INST_DATA_PATH_DECODE_RF_n2251, DLX_INST_DATA_PATH_DECODE_RF_n2250, 
      DLX_INST_DATA_PATH_DECODE_RF_n2249, DLX_INST_DATA_PATH_DECODE_RF_n2248, 
      DLX_INST_DATA_PATH_DECODE_RF_n2247, DLX_INST_DATA_PATH_DECODE_RF_n2246, 
      DLX_INST_DATA_PATH_DECODE_RF_n2245, DLX_INST_DATA_PATH_DECODE_RF_n2244, 
      DLX_INST_DATA_PATH_DECODE_RF_n2243, DLX_INST_DATA_PATH_DECODE_RF_n2242, 
      DLX_INST_DATA_PATH_DECODE_RF_n2241, DLX_INST_DATA_PATH_DECODE_RF_n2240, 
      DLX_INST_DATA_PATH_DECODE_RF_n2239, DLX_INST_DATA_PATH_DECODE_RF_n2238, 
      DLX_INST_DATA_PATH_DECODE_RF_n2237, DLX_INST_DATA_PATH_DECODE_RF_n2236, 
      DLX_INST_DATA_PATH_DECODE_RF_n2235, DLX_INST_DATA_PATH_DECODE_RF_n2234, 
      DLX_INST_DATA_PATH_DECODE_RF_n2233, DLX_INST_DATA_PATH_DECODE_RF_n2232, 
      DLX_INST_DATA_PATH_DECODE_RF_n2231, DLX_INST_DATA_PATH_DECODE_RF_n2230, 
      DLX_INST_DATA_PATH_DECODE_RF_n2229, DLX_INST_DATA_PATH_DECODE_RF_n2228, 
      DLX_INST_DATA_PATH_DECODE_RF_n2227, DLX_INST_DATA_PATH_DECODE_RF_n2226, 
      DLX_INST_DATA_PATH_DECODE_RF_n2225, DLX_INST_DATA_PATH_DECODE_RF_n2224, 
      DLX_INST_DATA_PATH_DECODE_RF_n2223, DLX_INST_DATA_PATH_DECODE_RF_n2222, 
      DLX_INST_DATA_PATH_DECODE_RF_n2221, DLX_INST_DATA_PATH_DECODE_RF_n2220, 
      DLX_INST_DATA_PATH_DECODE_RF_n2219, DLX_INST_DATA_PATH_DECODE_RF_n2218, 
      DLX_INST_DATA_PATH_DECODE_RF_n2217, DLX_INST_DATA_PATH_DECODE_RF_n2216, 
      DLX_INST_DATA_PATH_DECODE_RF_n2215, DLX_INST_DATA_PATH_DECODE_RF_n2214, 
      DLX_INST_DATA_PATH_DECODE_RF_n2213, DLX_INST_DATA_PATH_DECODE_RF_n2212, 
      DLX_INST_DATA_PATH_DECODE_RF_n2211, DLX_INST_DATA_PATH_DECODE_RF_n2210, 
      DLX_INST_DATA_PATH_DECODE_RF_n2209, DLX_INST_DATA_PATH_DECODE_RF_n2208, 
      DLX_INST_DATA_PATH_DECODE_RF_n2207, DLX_INST_DATA_PATH_DECODE_RF_n2206, 
      DLX_INST_DATA_PATH_DECODE_RF_n2205, DLX_INST_DATA_PATH_DECODE_RF_n2204, 
      DLX_INST_DATA_PATH_DECODE_RF_n2203, DLX_INST_DATA_PATH_DECODE_RF_n2202, 
      DLX_INST_DATA_PATH_DECODE_RF_n2201, DLX_INST_DATA_PATH_DECODE_RF_n2200, 
      DLX_INST_DATA_PATH_DECODE_RF_n2199, DLX_INST_DATA_PATH_DECODE_RF_n2198, 
      DLX_INST_DATA_PATH_DECODE_RF_n2197, DLX_INST_DATA_PATH_DECODE_RF_n2196, 
      DLX_INST_DATA_PATH_DECODE_RF_n2195, DLX_INST_DATA_PATH_DECODE_RF_n2194, 
      DLX_INST_DATA_PATH_DECODE_RF_n2193, DLX_INST_DATA_PATH_DECODE_RF_n2192, 
      DLX_INST_DATA_PATH_DECODE_RF_n2191, DLX_INST_DATA_PATH_DECODE_RF_n2190, 
      DLX_INST_DATA_PATH_DECODE_RF_n2189, DLX_INST_DATA_PATH_DECODE_RF_n2188, 
      DLX_INST_DATA_PATH_DECODE_RF_n2187, DLX_INST_DATA_PATH_DECODE_RF_n2186, 
      DLX_INST_DATA_PATH_DECODE_RF_n2185, DLX_INST_DATA_PATH_DECODE_RF_n2184, 
      DLX_INST_DATA_PATH_DECODE_RF_n2183, DLX_INST_DATA_PATH_DECODE_RF_n2182, 
      DLX_INST_DATA_PATH_DECODE_RF_n2181, DLX_INST_DATA_PATH_DECODE_RF_n2180, 
      DLX_INST_DATA_PATH_DECODE_RF_n2179, DLX_INST_DATA_PATH_DECODE_RF_n2178, 
      DLX_INST_DATA_PATH_DECODE_RF_n2177, DLX_INST_DATA_PATH_DECODE_RF_n2176, 
      DLX_INST_DATA_PATH_DECODE_RF_n2175, DLX_INST_DATA_PATH_DECODE_RF_n2174, 
      DLX_INST_DATA_PATH_DECODE_RF_n2173, DLX_INST_DATA_PATH_DECODE_RF_n2172, 
      DLX_INST_DATA_PATH_DECODE_RF_n2171, DLX_INST_DATA_PATH_DECODE_RF_n2170, 
      DLX_INST_DATA_PATH_DECODE_RF_n2169, DLX_INST_DATA_PATH_DECODE_RF_n2168, 
      DLX_INST_DATA_PATH_DECODE_RF_n2167, DLX_INST_DATA_PATH_DECODE_RF_n2166, 
      DLX_INST_DATA_PATH_DECODE_RF_n2165, DLX_INST_DATA_PATH_DECODE_RF_n2164, 
      DLX_INST_DATA_PATH_DECODE_RF_n2163, DLX_INST_DATA_PATH_DECODE_RF_n2162, 
      DLX_INST_DATA_PATH_DECODE_RF_n2161, DLX_INST_DATA_PATH_DECODE_RF_n2160, 
      DLX_INST_DATA_PATH_DECODE_RF_n2159, DLX_INST_DATA_PATH_DECODE_RF_n2158, 
      DLX_INST_DATA_PATH_DECODE_RF_n2157, DLX_INST_DATA_PATH_DECODE_RF_n2156, 
      DLX_INST_DATA_PATH_DECODE_RF_n2155, DLX_INST_DATA_PATH_DECODE_RF_n2154, 
      DLX_INST_DATA_PATH_DECODE_RF_n2153, DLX_INST_DATA_PATH_DECODE_RF_n2152, 
      DLX_INST_DATA_PATH_DECODE_RF_n2151, DLX_INST_DATA_PATH_DECODE_RF_n2150, 
      DLX_INST_DATA_PATH_DECODE_RF_n2149, DLX_INST_DATA_PATH_DECODE_RF_n2148, 
      DLX_INST_DATA_PATH_DECODE_RF_n2147, DLX_INST_DATA_PATH_DECODE_RF_n2146, 
      DLX_INST_DATA_PATH_DECODE_RF_n2145, DLX_INST_DATA_PATH_DECODE_RF_n2144, 
      DLX_INST_DATA_PATH_DECODE_RF_n2143, DLX_INST_DATA_PATH_DECODE_RF_n2142, 
      DLX_INST_DATA_PATH_DECODE_RF_n2141, DLX_INST_DATA_PATH_DECODE_RF_n2140, 
      DLX_INST_DATA_PATH_DECODE_RF_n2139, DLX_INST_DATA_PATH_DECODE_RF_n2138, 
      DLX_INST_DATA_PATH_DECODE_RF_n2137, DLX_INST_DATA_PATH_DECODE_RF_n2136, 
      DLX_INST_DATA_PATH_DECODE_RF_n2135, DLX_INST_DATA_PATH_DECODE_RF_n2134, 
      DLX_INST_DATA_PATH_DECODE_RF_n2133, DLX_INST_DATA_PATH_DECODE_RF_n2132, 
      DLX_INST_DATA_PATH_DECODE_RF_n2131, DLX_INST_DATA_PATH_DECODE_RF_n2130, 
      DLX_INST_DATA_PATH_DECODE_RF_n2129, DLX_INST_DATA_PATH_DECODE_RF_n2128, 
      DLX_INST_DATA_PATH_DECODE_RF_n2127, DLX_INST_DATA_PATH_DECODE_RF_n2126, 
      DLX_INST_DATA_PATH_DECODE_RF_n2125, DLX_INST_DATA_PATH_DECODE_RF_n2124, 
      DLX_INST_DATA_PATH_DECODE_RF_n2123, DLX_INST_DATA_PATH_DECODE_RF_n2122, 
      DLX_INST_DATA_PATH_DECODE_RF_n2121, DLX_INST_DATA_PATH_DECODE_RF_n2120, 
      DLX_INST_DATA_PATH_DECODE_RF_n2119, DLX_INST_DATA_PATH_DECODE_RF_n2118, 
      DLX_INST_DATA_PATH_DECODE_RF_n2117, DLX_INST_DATA_PATH_DECODE_RF_n2116, 
      DLX_INST_DATA_PATH_DECODE_RF_n2115, DLX_INST_DATA_PATH_DECODE_RF_n2114, 
      DLX_INST_DATA_PATH_DECODE_RF_n2113, DLX_INST_DATA_PATH_DECODE_RF_n2112, 
      DLX_INST_DATA_PATH_DECODE_RF_n2111, DLX_INST_DATA_PATH_DECODE_RF_n2110, 
      DLX_INST_DATA_PATH_DECODE_RF_n2109, DLX_INST_DATA_PATH_DECODE_RF_n2108, 
      DLX_INST_DATA_PATH_DECODE_RF_n2107, DLX_INST_DATA_PATH_DECODE_RF_n2106, 
      DLX_INST_DATA_PATH_DECODE_RF_n2105, DLX_INST_DATA_PATH_DECODE_RF_n2104, 
      DLX_INST_DATA_PATH_DECODE_RF_n2103, DLX_INST_DATA_PATH_DECODE_RF_n2102, 
      DLX_INST_DATA_PATH_DECODE_RF_n2101, DLX_INST_DATA_PATH_DECODE_RF_n2100, 
      DLX_INST_DATA_PATH_DECODE_RF_n2099, DLX_INST_DATA_PATH_DECODE_RF_n2098, 
      DLX_INST_DATA_PATH_DECODE_RF_n2097, DLX_INST_DATA_PATH_DECODE_RF_n2096, 
      DLX_INST_DATA_PATH_DECODE_RF_n2095, DLX_INST_DATA_PATH_DECODE_RF_n2094, 
      DLX_INST_DATA_PATH_DECODE_RF_n2093, DLX_INST_DATA_PATH_DECODE_RF_n2092, 
      DLX_INST_DATA_PATH_DECODE_RF_n2091, DLX_INST_DATA_PATH_DECODE_RF_n2090, 
      DLX_INST_DATA_PATH_DECODE_RF_n2089, DLX_INST_DATA_PATH_DECODE_RF_n2088, 
      DLX_INST_DATA_PATH_DECODE_RF_n2087, DLX_INST_DATA_PATH_DECODE_RF_n2086, 
      DLX_INST_DATA_PATH_DECODE_RF_n2085, DLX_INST_DATA_PATH_DECODE_RF_n2084, 
      DLX_INST_DATA_PATH_DECODE_RF_n2083, DLX_INST_DATA_PATH_DECODE_RF_n2082, 
      DLX_INST_DATA_PATH_DECODE_RF_n2081, DLX_INST_DATA_PATH_DECODE_RF_n2080, 
      DLX_INST_DATA_PATH_DECODE_RF_n2079, DLX_INST_DATA_PATH_DECODE_RF_n2078, 
      DLX_INST_DATA_PATH_DECODE_RF_n2077, DLX_INST_DATA_PATH_DECODE_RF_n2076, 
      DLX_INST_DATA_PATH_DECODE_RF_n2075, DLX_INST_DATA_PATH_DECODE_RF_n2074, 
      DLX_INST_DATA_PATH_DECODE_RF_n2073, DLX_INST_DATA_PATH_DECODE_RF_n2072, 
      DLX_INST_DATA_PATH_DECODE_RF_n2071, DLX_INST_DATA_PATH_DECODE_RF_n2070, 
      DLX_INST_DATA_PATH_DECODE_RF_n2069, DLX_INST_DATA_PATH_DECODE_RF_n2068, 
      DLX_INST_DATA_PATH_DECODE_RF_n2067, DLX_INST_DATA_PATH_DECODE_RF_n2066, 
      DLX_INST_DATA_PATH_DECODE_RF_n2065, DLX_INST_DATA_PATH_DECODE_RF_n2064, 
      DLX_INST_DATA_PATH_DECODE_RF_n2063, DLX_INST_DATA_PATH_DECODE_RF_n2062, 
      DLX_INST_DATA_PATH_DECODE_RF_n2061, DLX_INST_DATA_PATH_DECODE_RF_n2060, 
      DLX_INST_DATA_PATH_DECODE_RF_n2059, DLX_INST_DATA_PATH_DECODE_RF_n2058, 
      DLX_INST_DATA_PATH_DECODE_RF_n2057, DLX_INST_DATA_PATH_DECODE_RF_n2056, 
      DLX_INST_DATA_PATH_DECODE_RF_n2055, DLX_INST_DATA_PATH_DECODE_RF_n2054, 
      DLX_INST_DATA_PATH_DECODE_RF_n2053, DLX_INST_DATA_PATH_DECODE_RF_n2052, 
      DLX_INST_DATA_PATH_DECODE_RF_n2051, DLX_INST_DATA_PATH_DECODE_RF_n2050, 
      DLX_INST_DATA_PATH_DECODE_RF_n2049, DLX_INST_DATA_PATH_DECODE_RF_n2048, 
      DLX_INST_DATA_PATH_DECODE_RF_n2047, DLX_INST_DATA_PATH_DECODE_RF_n2046, 
      DLX_INST_DATA_PATH_DECODE_RF_n2045, DLX_INST_DATA_PATH_DECODE_RF_n2044, 
      DLX_INST_DATA_PATH_DECODE_RF_n2043, DLX_INST_DATA_PATH_DECODE_RF_n2042, 
      DLX_INST_DATA_PATH_DECODE_RF_n2041, DLX_INST_DATA_PATH_DECODE_RF_n2040, 
      DLX_INST_DATA_PATH_DECODE_RF_n2039, DLX_INST_DATA_PATH_DECODE_RF_n2038, 
      DLX_INST_DATA_PATH_DECODE_RF_n2037, DLX_INST_DATA_PATH_DECODE_RF_n2036, 
      DLX_INST_DATA_PATH_DECODE_RF_n2035, DLX_INST_DATA_PATH_DECODE_RF_n2034, 
      DLX_INST_DATA_PATH_DECODE_RF_n2033, DLX_INST_DATA_PATH_DECODE_RF_n2032, 
      DLX_INST_DATA_PATH_DECODE_RF_n2031, DLX_INST_DATA_PATH_DECODE_RF_n2030, 
      DLX_INST_DATA_PATH_DECODE_RF_n2029, DLX_INST_DATA_PATH_DECODE_RF_n2028, 
      DLX_INST_DATA_PATH_DECODE_RF_n2027, DLX_INST_DATA_PATH_DECODE_RF_n2026, 
      DLX_INST_DATA_PATH_DECODE_RF_n2025, DLX_INST_DATA_PATH_DECODE_RF_n2024, 
      DLX_INST_DATA_PATH_DECODE_RF_n2023, DLX_INST_DATA_PATH_DECODE_RF_n2022, 
      DLX_INST_DATA_PATH_DECODE_RF_n2021, DLX_INST_DATA_PATH_DECODE_RF_n2020, 
      DLX_INST_DATA_PATH_DECODE_RF_n2019, DLX_INST_DATA_PATH_DECODE_RF_n2018, 
      DLX_INST_DATA_PATH_DECODE_RF_n2017, DLX_INST_DATA_PATH_DECODE_RF_n2016, 
      DLX_INST_DATA_PATH_DECODE_RF_n2015, DLX_INST_DATA_PATH_DECODE_RF_n2014, 
      DLX_INST_DATA_PATH_DECODE_RF_n2013, DLX_INST_DATA_PATH_DECODE_RF_n2012, 
      DLX_INST_DATA_PATH_DECODE_RF_n2011, DLX_INST_DATA_PATH_DECODE_RF_n2010, 
      DLX_INST_DATA_PATH_DECODE_RF_n2009, DLX_INST_DATA_PATH_DECODE_RF_n2008, 
      DLX_INST_DATA_PATH_DECODE_RF_n2007, DLX_INST_DATA_PATH_DECODE_RF_n2006, 
      DLX_INST_DATA_PATH_DECODE_RF_n2005, DLX_INST_DATA_PATH_DECODE_RF_n2004, 
      DLX_INST_DATA_PATH_DECODE_RF_n2003, DLX_INST_DATA_PATH_DECODE_RF_n2002, 
      DLX_INST_DATA_PATH_DECODE_RF_n2001, DLX_INST_DATA_PATH_DECODE_RF_n2000, 
      DLX_INST_DATA_PATH_DECODE_RF_n1999, DLX_INST_DATA_PATH_DECODE_RF_n1998, 
      DLX_INST_DATA_PATH_DECODE_RF_n1997, DLX_INST_DATA_PATH_DECODE_RF_n1996, 
      DLX_INST_DATA_PATH_DECODE_RF_n1995, DLX_INST_DATA_PATH_DECODE_RF_n1994, 
      DLX_INST_DATA_PATH_DECODE_RF_n1993, DLX_INST_DATA_PATH_DECODE_RF_n1992, 
      DLX_INST_DATA_PATH_DECODE_RF_n1991, DLX_INST_DATA_PATH_DECODE_RF_n1990, 
      DLX_INST_DATA_PATH_DECODE_RF_n1989, DLX_INST_DATA_PATH_DECODE_RF_n1988, 
      DLX_INST_DATA_PATH_DECODE_RF_n1987, DLX_INST_DATA_PATH_DECODE_RF_n1986, 
      DLX_INST_DATA_PATH_DECODE_RF_n1985, DLX_INST_DATA_PATH_DECODE_RF_n1984, 
      DLX_INST_DATA_PATH_DECODE_RF_n1983, DLX_INST_DATA_PATH_DECODE_RF_n1982, 
      DLX_INST_DATA_PATH_DECODE_RF_n1981, DLX_INST_DATA_PATH_DECODE_RF_n1980, 
      DLX_INST_DATA_PATH_DECODE_RF_n1979, DLX_INST_DATA_PATH_DECODE_RF_n1978, 
      DLX_INST_DATA_PATH_DECODE_RF_n1977, DLX_INST_DATA_PATH_DECODE_RF_n1976, 
      DLX_INST_DATA_PATH_DECODE_RF_n1975, DLX_INST_DATA_PATH_DECODE_RF_n1974, 
      DLX_INST_DATA_PATH_DECODE_RF_n1973, DLX_INST_DATA_PATH_DECODE_RF_n1972, 
      DLX_INST_DATA_PATH_DECODE_RF_n1971, DLX_INST_DATA_PATH_DECODE_RF_n1970, 
      DLX_INST_DATA_PATH_DECODE_RF_n1969, DLX_INST_DATA_PATH_DECODE_RF_n1968, 
      DLX_INST_DATA_PATH_DECODE_RF_n1967, DLX_INST_DATA_PATH_DECODE_RF_n1966, 
      DLX_INST_DATA_PATH_DECODE_RF_n1965, DLX_INST_DATA_PATH_DECODE_RF_n1964, 
      DLX_INST_DATA_PATH_DECODE_RF_n1963, DLX_INST_DATA_PATH_DECODE_RF_n1962, 
      DLX_INST_DATA_PATH_DECODE_RF_n1961, DLX_INST_DATA_PATH_DECODE_RF_n1960, 
      DLX_INST_DATA_PATH_DECODE_RF_n1959, DLX_INST_DATA_PATH_DECODE_RF_n1958, 
      DLX_INST_DATA_PATH_DECODE_RF_n1957, DLX_INST_DATA_PATH_DECODE_RF_n1956, 
      DLX_INST_DATA_PATH_DECODE_RF_n1955, DLX_INST_DATA_PATH_DECODE_RF_n1954, 
      DLX_INST_DATA_PATH_DECODE_RF_n1953, DLX_INST_DATA_PATH_DECODE_RF_n1952, 
      DLX_INST_DATA_PATH_DECODE_RF_n1951, DLX_INST_DATA_PATH_DECODE_RF_n1950, 
      DLX_INST_DATA_PATH_DECODE_RF_n1949, DLX_INST_DATA_PATH_DECODE_RF_n1948, 
      DLX_INST_DATA_PATH_DECODE_RF_n1947, DLX_INST_DATA_PATH_DECODE_RF_n1946, 
      DLX_INST_DATA_PATH_DECODE_RF_n1945, DLX_INST_DATA_PATH_DECODE_RF_n1944, 
      DLX_INST_DATA_PATH_DECODE_RF_n1943, DLX_INST_DATA_PATH_DECODE_RF_n1942, 
      DLX_INST_DATA_PATH_DECODE_RF_n1941, DLX_INST_DATA_PATH_DECODE_RF_n1940, 
      DLX_INST_DATA_PATH_DECODE_RF_n1939, DLX_INST_DATA_PATH_DECODE_RF_n1938, 
      DLX_INST_DATA_PATH_DECODE_RF_n1937, DLX_INST_DATA_PATH_DECODE_RF_n1936, 
      DLX_INST_DATA_PATH_DECODE_RF_n1935, DLX_INST_DATA_PATH_DECODE_RF_n1934, 
      DLX_INST_DATA_PATH_DECODE_RF_n1933, DLX_INST_DATA_PATH_DECODE_RF_n1932, 
      DLX_INST_DATA_PATH_DECODE_RF_n1931, DLX_INST_DATA_PATH_DECODE_RF_n1930, 
      DLX_INST_DATA_PATH_DECODE_RF_n1929, DLX_INST_DATA_PATH_DECODE_RF_n1928, 
      DLX_INST_DATA_PATH_DECODE_RF_n1927, DLX_INST_DATA_PATH_DECODE_RF_n1926, 
      DLX_INST_DATA_PATH_DECODE_RF_n1925, DLX_INST_DATA_PATH_DECODE_RF_n1924, 
      DLX_INST_DATA_PATH_DECODE_RF_n1923, DLX_INST_DATA_PATH_DECODE_RF_n1922, 
      DLX_INST_DATA_PATH_DECODE_RF_n1921, DLX_INST_DATA_PATH_DECODE_RF_n1920, 
      DLX_INST_DATA_PATH_DECODE_RF_n1919, DLX_INST_DATA_PATH_DECODE_RF_n1918, 
      DLX_INST_DATA_PATH_DECODE_RF_n1917, DLX_INST_DATA_PATH_DECODE_RF_n1916, 
      DLX_INST_DATA_PATH_DECODE_RF_n1915, DLX_INST_DATA_PATH_DECODE_RF_n1914, 
      DLX_INST_DATA_PATH_DECODE_RF_n1913, DLX_INST_DATA_PATH_DECODE_RF_n1912, 
      DLX_INST_DATA_PATH_DECODE_RF_n1911, DLX_INST_DATA_PATH_DECODE_RF_n1910, 
      DLX_INST_DATA_PATH_DECODE_RF_n1909, DLX_INST_DATA_PATH_DECODE_RF_n1908, 
      DLX_INST_DATA_PATH_DECODE_RF_n1907, DLX_INST_DATA_PATH_DECODE_RF_n1906, 
      DLX_INST_DATA_PATH_DECODE_RF_n1905, DLX_INST_DATA_PATH_DECODE_RF_n1904, 
      DLX_INST_DATA_PATH_DECODE_RF_n1903, DLX_INST_DATA_PATH_DECODE_RF_n1902, 
      DLX_INST_DATA_PATH_DECODE_RF_n1901, DLX_INST_DATA_PATH_DECODE_RF_n1900, 
      DLX_INST_DATA_PATH_DECODE_RF_n1899, DLX_INST_DATA_PATH_DECODE_RF_n1898, 
      DLX_INST_DATA_PATH_DECODE_RF_n1897, DLX_INST_DATA_PATH_DECODE_RF_n1896, 
      DLX_INST_DATA_PATH_DECODE_RF_n1895, DLX_INST_DATA_PATH_DECODE_RF_n1894, 
      DLX_INST_DATA_PATH_DECODE_RF_n1893, DLX_INST_DATA_PATH_DECODE_RF_n1892, 
      DLX_INST_DATA_PATH_DECODE_RF_n1891, DLX_INST_DATA_PATH_DECODE_RF_n1890, 
      DLX_INST_DATA_PATH_DECODE_RF_n1889, DLX_INST_DATA_PATH_DECODE_RF_n1888, 
      DLX_INST_DATA_PATH_DECODE_RF_n1887, DLX_INST_DATA_PATH_DECODE_RF_n1886, 
      DLX_INST_DATA_PATH_DECODE_RF_n1885, DLX_INST_DATA_PATH_DECODE_RF_n1884, 
      DLX_INST_DATA_PATH_DECODE_RF_n1883, DLX_INST_DATA_PATH_DECODE_RF_n1882, 
      DLX_INST_DATA_PATH_DECODE_RF_n1881, DLX_INST_DATA_PATH_DECODE_RF_n1880, 
      DLX_INST_DATA_PATH_DECODE_RF_n1879, DLX_INST_DATA_PATH_DECODE_RF_n1878, 
      DLX_INST_DATA_PATH_DECODE_RF_n1877, DLX_INST_DATA_PATH_DECODE_RF_n1876, 
      DLX_INST_DATA_PATH_DECODE_RF_n1875, DLX_INST_DATA_PATH_DECODE_RF_n1874, 
      DLX_INST_DATA_PATH_DECODE_RF_n1873, DLX_INST_DATA_PATH_DECODE_RF_n1872, 
      DLX_INST_DATA_PATH_DECODE_RF_n1871, DLX_INST_DATA_PATH_DECODE_RF_n1870, 
      DLX_INST_DATA_PATH_DECODE_RF_n1869, DLX_INST_DATA_PATH_DECODE_RF_n1868, 
      DLX_INST_DATA_PATH_DECODE_RF_n1867, DLX_INST_DATA_PATH_DECODE_RF_n1866, 
      DLX_INST_DATA_PATH_DECODE_RF_n1865, DLX_INST_DATA_PATH_DECODE_RF_n1864, 
      DLX_INST_DATA_PATH_DECODE_RF_n1863, DLX_INST_DATA_PATH_DECODE_RF_n1862, 
      DLX_INST_DATA_PATH_DECODE_RF_n1861, DLX_INST_DATA_PATH_DECODE_RF_n1860, 
      DLX_INST_DATA_PATH_DECODE_RF_n1859, DLX_INST_DATA_PATH_DECODE_RF_n1858, 
      DLX_INST_DATA_PATH_DECODE_RF_n1857, DLX_INST_DATA_PATH_DECODE_RF_n1856, 
      DLX_INST_DATA_PATH_DECODE_RF_n1855, DLX_INST_DATA_PATH_DECODE_RF_n1854, 
      DLX_INST_DATA_PATH_DECODE_RF_n1853, DLX_INST_DATA_PATH_DECODE_RF_n1852, 
      DLX_INST_DATA_PATH_DECODE_RF_n1851, DLX_INST_DATA_PATH_DECODE_RF_n1850, 
      DLX_INST_DATA_PATH_DECODE_RF_n1849, DLX_INST_DATA_PATH_DECODE_RF_n1848, 
      DLX_INST_DATA_PATH_DECODE_RF_n1847, DLX_INST_DATA_PATH_DECODE_RF_n1846, 
      DLX_INST_DATA_PATH_DECODE_RF_n1845, DLX_INST_DATA_PATH_DECODE_RF_n1844, 
      DLX_INST_DATA_PATH_DECODE_RF_n1843, DLX_INST_DATA_PATH_DECODE_RF_n1842, 
      DLX_INST_DATA_PATH_DECODE_RF_n1841, DLX_INST_DATA_PATH_DECODE_RF_n1840, 
      DLX_INST_DATA_PATH_DECODE_RF_n1839, DLX_INST_DATA_PATH_DECODE_RF_n1838, 
      DLX_INST_DATA_PATH_DECODE_RF_n1837, DLX_INST_DATA_PATH_DECODE_RF_n1836, 
      DLX_INST_DATA_PATH_DECODE_RF_n1835, DLX_INST_DATA_PATH_DECODE_RF_n1834, 
      DLX_INST_DATA_PATH_DECODE_RF_n1833, DLX_INST_DATA_PATH_DECODE_RF_n1832, 
      DLX_INST_DATA_PATH_DECODE_RF_n1831, DLX_INST_DATA_PATH_DECODE_RF_n1830, 
      DLX_INST_DATA_PATH_DECODE_RF_n1829, DLX_INST_DATA_PATH_DECODE_RF_n1828, 
      DLX_INST_DATA_PATH_DECODE_RF_n1827, DLX_INST_DATA_PATH_DECODE_RF_n1826, 
      DLX_INST_DATA_PATH_DECODE_RF_n1825, DLX_INST_DATA_PATH_DECODE_RF_n1824, 
      DLX_INST_DATA_PATH_DECODE_RF_n1823, DLX_INST_DATA_PATH_DECODE_RF_n1822, 
      DLX_INST_DATA_PATH_DECODE_RF_n1821, DLX_INST_DATA_PATH_DECODE_RF_n1820, 
      DLX_INST_DATA_PATH_DECODE_RF_n1819, DLX_INST_DATA_PATH_DECODE_RF_n1818, 
      DLX_INST_DATA_PATH_DECODE_RF_n1817, DLX_INST_DATA_PATH_DECODE_RF_n1816, 
      DLX_INST_DATA_PATH_DECODE_RF_n1815, DLX_INST_DATA_PATH_DECODE_RF_n1814, 
      DLX_INST_DATA_PATH_DECODE_RF_n1813, DLX_INST_DATA_PATH_DECODE_RF_n1812, 
      DLX_INST_DATA_PATH_DECODE_RF_n1811, DLX_INST_DATA_PATH_DECODE_RF_n1810, 
      DLX_INST_DATA_PATH_DECODE_RF_n1809, DLX_INST_DATA_PATH_DECODE_RF_n1808, 
      DLX_INST_DATA_PATH_DECODE_RF_n1807, DLX_INST_DATA_PATH_DECODE_RF_n1806, 
      DLX_INST_DATA_PATH_DECODE_RF_n1805, DLX_INST_DATA_PATH_DECODE_RF_n1804, 
      DLX_INST_DATA_PATH_DECODE_RF_n1803, DLX_INST_DATA_PATH_DECODE_RF_n1802, 
      DLX_INST_DATA_PATH_DECODE_RF_n1801, DLX_INST_DATA_PATH_DECODE_RF_n1800, 
      DLX_INST_DATA_PATH_DECODE_RF_n1799, DLX_INST_DATA_PATH_DECODE_RF_n1798, 
      DLX_INST_DATA_PATH_DECODE_RF_n1797, DLX_INST_DATA_PATH_DECODE_RF_n1796, 
      DLX_INST_DATA_PATH_DECODE_RF_n1795, DLX_INST_DATA_PATH_DECODE_RF_n1794, 
      DLX_INST_DATA_PATH_DECODE_RF_n1793, DLX_INST_DATA_PATH_DECODE_RF_n1792, 
      DLX_INST_DATA_PATH_DECODE_RF_n1791, DLX_INST_DATA_PATH_DECODE_RF_n1790, 
      DLX_INST_DATA_PATH_DECODE_RF_n1789, DLX_INST_DATA_PATH_DECODE_RF_n1788, 
      DLX_INST_DATA_PATH_DECODE_RF_n1787, DLX_INST_DATA_PATH_DECODE_RF_n1786, 
      DLX_INST_DATA_PATH_DECODE_RF_n1785, DLX_INST_DATA_PATH_DECODE_RF_n1784, 
      DLX_INST_DATA_PATH_DECODE_RF_n1783, DLX_INST_DATA_PATH_DECODE_RF_n1782, 
      DLX_INST_DATA_PATH_DECODE_RF_n1781, DLX_INST_DATA_PATH_DECODE_RF_n1780, 
      DLX_INST_DATA_PATH_DECODE_RF_n1779, DLX_INST_DATA_PATH_DECODE_RF_n1778, 
      DLX_INST_DATA_PATH_DECODE_RF_n1777, DLX_INST_DATA_PATH_DECODE_RF_n1776, 
      DLX_INST_DATA_PATH_DECODE_RF_n1775, DLX_INST_DATA_PATH_DECODE_RF_n1774, 
      DLX_INST_DATA_PATH_DECODE_RF_n1773, DLX_INST_DATA_PATH_DECODE_RF_n1772, 
      DLX_INST_DATA_PATH_DECODE_RF_n1771, DLX_INST_DATA_PATH_DECODE_RF_n1770, 
      DLX_INST_DATA_PATH_DECODE_RF_n1769, DLX_INST_DATA_PATH_DECODE_RF_n1768, 
      DLX_INST_DATA_PATH_DECODE_RF_n1767, DLX_INST_DATA_PATH_DECODE_RF_n1766, 
      DLX_INST_DATA_PATH_DECODE_RF_n1765, DLX_INST_DATA_PATH_DECODE_RF_n1764, 
      DLX_INST_DATA_PATH_DECODE_RF_n1763, DLX_INST_DATA_PATH_DECODE_RF_n1762, 
      DLX_INST_DATA_PATH_DECODE_RF_n1761, DLX_INST_DATA_PATH_DECODE_RF_n1760, 
      DLX_INST_DATA_PATH_DECODE_RF_n1759, DLX_INST_DATA_PATH_DECODE_RF_n1758, 
      DLX_INST_DATA_PATH_DECODE_RF_n1757, DLX_INST_DATA_PATH_DECODE_RF_n1756, 
      DLX_INST_DATA_PATH_DECODE_RF_n1755, DLX_INST_DATA_PATH_DECODE_RF_n1754, 
      DLX_INST_DATA_PATH_DECODE_RF_n1753, DLX_INST_DATA_PATH_DECODE_RF_n1752, 
      DLX_INST_DATA_PATH_DECODE_RF_n1751, DLX_INST_DATA_PATH_DECODE_RF_n1750, 
      DLX_INST_DATA_PATH_DECODE_RF_n1749, DLX_INST_DATA_PATH_DECODE_RF_n1748, 
      DLX_INST_DATA_PATH_DECODE_RF_n1747, DLX_INST_DATA_PATH_DECODE_RF_n1746, 
      DLX_INST_DATA_PATH_DECODE_RF_n1745, DLX_INST_DATA_PATH_DECODE_RF_n1744, 
      DLX_INST_DATA_PATH_DECODE_RF_n1743, DLX_INST_DATA_PATH_DECODE_RF_n1742, 
      DLX_INST_DATA_PATH_DECODE_RF_n1741, DLX_INST_DATA_PATH_DECODE_RF_n1740, 
      DLX_INST_DATA_PATH_DECODE_RF_n1739, DLX_INST_DATA_PATH_DECODE_RF_n1738, 
      DLX_INST_DATA_PATH_DECODE_RF_n1737, DLX_INST_DATA_PATH_DECODE_RF_n1736, 
      DLX_INST_DATA_PATH_DECODE_RF_n1735, DLX_INST_DATA_PATH_DECODE_RF_n1734, 
      DLX_INST_DATA_PATH_DECODE_RF_n1733, DLX_INST_DATA_PATH_DECODE_RF_n1732, 
      DLX_INST_DATA_PATH_DECODE_RF_n1731, DLX_INST_DATA_PATH_DECODE_RF_n1730, 
      DLX_INST_DATA_PATH_DECODE_RF_n1729, DLX_INST_DATA_PATH_DECODE_RF_n1728, 
      DLX_INST_DATA_PATH_DECODE_RF_n1727, DLX_INST_DATA_PATH_DECODE_RF_n1726, 
      DLX_INST_DATA_PATH_DECODE_RF_n1725, DLX_INST_DATA_PATH_DECODE_RF_n1724, 
      DLX_INST_DATA_PATH_DECODE_RF_n1723, DLX_INST_DATA_PATH_DECODE_RF_n1722, 
      DLX_INST_DATA_PATH_DECODE_RF_n1721, DLX_INST_DATA_PATH_DECODE_RF_n1720, 
      DLX_INST_DATA_PATH_DECODE_RF_n1719, DLX_INST_DATA_PATH_DECODE_RF_n1718, 
      DLX_INST_DATA_PATH_DECODE_RF_n1717, DLX_INST_DATA_PATH_DECODE_RF_n1716, 
      DLX_INST_DATA_PATH_DECODE_RF_n1715, DLX_INST_DATA_PATH_DECODE_RF_n1714, 
      DLX_INST_DATA_PATH_DECODE_RF_n1713, DLX_INST_DATA_PATH_DECODE_RF_n1712, 
      DLX_INST_DATA_PATH_DECODE_RF_n1711, DLX_INST_DATA_PATH_DECODE_RF_n1710, 
      DLX_INST_DATA_PATH_DECODE_RF_n1709, DLX_INST_DATA_PATH_DECODE_RF_n1708, 
      DLX_INST_DATA_PATH_DECODE_RF_n1707, DLX_INST_DATA_PATH_DECODE_RF_n1706, 
      DLX_INST_DATA_PATH_DECODE_RF_n1705, DLX_INST_DATA_PATH_DECODE_RF_n1704, 
      DLX_INST_DATA_PATH_DECODE_RF_n1703, DLX_INST_DATA_PATH_DECODE_RF_n1702, 
      DLX_INST_DATA_PATH_DECODE_RF_n1701, DLX_INST_DATA_PATH_DECODE_RF_n1700, 
      DLX_INST_DATA_PATH_DECODE_RF_n1699, DLX_INST_DATA_PATH_DECODE_RF_n1698, 
      DLX_INST_DATA_PATH_DECODE_RF_n1697, DLX_INST_DATA_PATH_DECODE_RF_n1696, 
      DLX_INST_DATA_PATH_DECODE_RF_n1695, DLX_INST_DATA_PATH_DECODE_RF_n1694, 
      DLX_INST_DATA_PATH_DECODE_RF_n1693, DLX_INST_DATA_PATH_DECODE_RF_n1692, 
      DLX_INST_DATA_PATH_DECODE_RF_n1691, DLX_INST_DATA_PATH_DECODE_RF_n1690, 
      DLX_INST_DATA_PATH_DECODE_RF_n1689, DLX_INST_DATA_PATH_DECODE_RF_n1688, 
      DLX_INST_DATA_PATH_DECODE_RF_n1687, DLX_INST_DATA_PATH_DECODE_RF_n1686, 
      DLX_INST_DATA_PATH_DECODE_RF_n1685, DLX_INST_DATA_PATH_DECODE_RF_n1684, 
      DLX_INST_DATA_PATH_DECODE_RF_n1683, DLX_INST_DATA_PATH_DECODE_RF_n1682, 
      DLX_INST_DATA_PATH_DECODE_RF_n1681, DLX_INST_DATA_PATH_DECODE_RF_n1680, 
      DLX_INST_DATA_PATH_DECODE_RF_n1679, DLX_INST_DATA_PATH_DECODE_RF_n1678, 
      DLX_INST_DATA_PATH_DECODE_RF_n1677, DLX_INST_DATA_PATH_DECODE_RF_n1676, 
      DLX_INST_DATA_PATH_DECODE_RF_n1675, DLX_INST_DATA_PATH_DECODE_RF_n1674, 
      DLX_INST_DATA_PATH_DECODE_RF_n1673, DLX_INST_DATA_PATH_DECODE_RF_n1672, 
      DLX_INST_DATA_PATH_DECODE_RF_n1671, DLX_INST_DATA_PATH_DECODE_RF_n1670, 
      DLX_INST_DATA_PATH_DECODE_RF_n1669, DLX_INST_DATA_PATH_DECODE_RF_n1668, 
      DLX_INST_DATA_PATH_DECODE_RF_n1667, DLX_INST_DATA_PATH_DECODE_RF_n1666, 
      DLX_INST_DATA_PATH_DECODE_RF_n1665, DLX_INST_DATA_PATH_DECODE_RF_n1664, 
      DLX_INST_DATA_PATH_DECODE_RF_n1663, DLX_INST_DATA_PATH_DECODE_RF_n1662, 
      DLX_INST_DATA_PATH_DECODE_RF_n1661, DLX_INST_DATA_PATH_DECODE_RF_n1660, 
      DLX_INST_DATA_PATH_DECODE_RF_n1659, DLX_INST_DATA_PATH_DECODE_RF_n1658, 
      DLX_INST_DATA_PATH_DECODE_RF_n1657, DLX_INST_DATA_PATH_DECODE_RF_n1656, 
      DLX_INST_DATA_PATH_DECODE_RF_n1655, DLX_INST_DATA_PATH_DECODE_RF_n1654, 
      DLX_INST_DATA_PATH_DECODE_RF_n1653, DLX_INST_DATA_PATH_DECODE_RF_n1652, 
      DLX_INST_DATA_PATH_DECODE_RF_n1651, DLX_INST_DATA_PATH_DECODE_RF_n1650, 
      DLX_INST_DATA_PATH_DECODE_RF_n1649, DLX_INST_DATA_PATH_DECODE_RF_n1648, 
      DLX_INST_DATA_PATH_DECODE_RF_n1647, DLX_INST_DATA_PATH_DECODE_RF_n1646, 
      DLX_INST_DATA_PATH_DECODE_RF_n1645, DLX_INST_DATA_PATH_DECODE_RF_n1644, 
      DLX_INST_DATA_PATH_DECODE_RF_n1643, DLX_INST_DATA_PATH_DECODE_RF_n1642, 
      DLX_INST_DATA_PATH_DECODE_RF_n1641, DLX_INST_DATA_PATH_DECODE_RF_n1640, 
      DLX_INST_DATA_PATH_DECODE_RF_n1639, DLX_INST_DATA_PATH_DECODE_RF_n1638, 
      DLX_INST_DATA_PATH_DECODE_RF_n1637, DLX_INST_DATA_PATH_DECODE_RF_n1636, 
      DLX_INST_DATA_PATH_DECODE_RF_n1635, DLX_INST_DATA_PATH_DECODE_RF_n1634, 
      DLX_INST_DATA_PATH_DECODE_RF_n1633, DLX_INST_DATA_PATH_DECODE_RF_n1632, 
      DLX_INST_DATA_PATH_DECODE_RF_n1631, DLX_INST_DATA_PATH_DECODE_RF_n1630, 
      DLX_INST_DATA_PATH_DECODE_RF_n1629, DLX_INST_DATA_PATH_DECODE_RF_n1628, 
      DLX_INST_DATA_PATH_DECODE_RF_n1627, DLX_INST_DATA_PATH_DECODE_RF_n1626, 
      DLX_INST_DATA_PATH_DECODE_RF_n1625, DLX_INST_DATA_PATH_DECODE_RF_n1624, 
      DLX_INST_DATA_PATH_DECODE_RF_n1623, DLX_INST_DATA_PATH_DECODE_RF_n1622, 
      DLX_INST_DATA_PATH_DECODE_RF_n1621, DLX_INST_DATA_PATH_DECODE_RF_n1620, 
      DLX_INST_DATA_PATH_DECODE_RF_n1619, DLX_INST_DATA_PATH_DECODE_RF_n1618, 
      DLX_INST_DATA_PATH_DECODE_RF_n1617, DLX_INST_DATA_PATH_DECODE_RF_n1616, 
      DLX_INST_DATA_PATH_DECODE_RF_n1615, DLX_INST_DATA_PATH_DECODE_RF_n1614, 
      DLX_INST_DATA_PATH_DECODE_RF_n1613, DLX_INST_DATA_PATH_DECODE_RF_n1612, 
      DLX_INST_DATA_PATH_DECODE_RF_n1611, DLX_INST_DATA_PATH_DECODE_RF_n1610, 
      DLX_INST_DATA_PATH_DECODE_RF_n1609, DLX_INST_DATA_PATH_DECODE_RF_n1608, 
      DLX_INST_DATA_PATH_DECODE_RF_n1607, DLX_INST_DATA_PATH_DECODE_RF_n1606, 
      DLX_INST_DATA_PATH_DECODE_RF_n1605, DLX_INST_DATA_PATH_DECODE_RF_n1604, 
      DLX_INST_DATA_PATH_DECODE_RF_n1603, DLX_INST_DATA_PATH_DECODE_RF_n1602, 
      DLX_INST_DATA_PATH_DECODE_RF_n1601, DLX_INST_DATA_PATH_DECODE_RF_n1600, 
      DLX_INST_DATA_PATH_DECODE_RF_n1599, DLX_INST_DATA_PATH_DECODE_RF_n1598, 
      DLX_INST_DATA_PATH_DECODE_RF_n1597, DLX_INST_DATA_PATH_DECODE_RF_n1596, 
      DLX_INST_DATA_PATH_DECODE_RF_n1595, DLX_INST_DATA_PATH_DECODE_RF_n1594, 
      DLX_INST_DATA_PATH_DECODE_RF_n1593, DLX_INST_DATA_PATH_DECODE_RF_n1592, 
      DLX_INST_DATA_PATH_DECODE_RF_n1591, DLX_INST_DATA_PATH_DECODE_RF_n1590, 
      DLX_INST_DATA_PATH_DECODE_RF_n1589, DLX_INST_DATA_PATH_DECODE_RF_n1588, 
      DLX_INST_DATA_PATH_DECODE_RF_n1587, DLX_INST_DATA_PATH_DECODE_RF_n1586, 
      DLX_INST_DATA_PATH_DECODE_RF_n1585, DLX_INST_DATA_PATH_DECODE_RF_n1584, 
      DLX_INST_DATA_PATH_DECODE_RF_n1583, DLX_INST_DATA_PATH_DECODE_RF_n1582, 
      DLX_INST_DATA_PATH_DECODE_RF_n1581, DLX_INST_DATA_PATH_DECODE_RF_n1580, 
      DLX_INST_DATA_PATH_DECODE_RF_n1579, DLX_INST_DATA_PATH_DECODE_RF_n1578, 
      DLX_INST_DATA_PATH_DECODE_RF_n1577, DLX_INST_DATA_PATH_DECODE_RF_n1576, 
      DLX_INST_DATA_PATH_DECODE_RF_n1575, DLX_INST_DATA_PATH_DECODE_RF_n1574, 
      DLX_INST_DATA_PATH_DECODE_RF_n1573, DLX_INST_DATA_PATH_DECODE_RF_n1572, 
      DLX_INST_DATA_PATH_DECODE_RF_n1571, DLX_INST_DATA_PATH_DECODE_RF_n1570, 
      DLX_INST_DATA_PATH_DECODE_RF_n1569, DLX_INST_DATA_PATH_DECODE_RF_n1568, 
      DLX_INST_DATA_PATH_DECODE_RF_n1567, DLX_INST_DATA_PATH_DECODE_RF_n1566, 
      DLX_INST_DATA_PATH_DECODE_RF_n1565, DLX_INST_DATA_PATH_DECODE_RF_n1564, 
      DLX_INST_DATA_PATH_DECODE_RF_n1563, DLX_INST_DATA_PATH_DECODE_RF_n1562, 
      DLX_INST_DATA_PATH_DECODE_RF_n1561, DLX_INST_DATA_PATH_DECODE_RF_n1560, 
      DLX_INST_DATA_PATH_DECODE_RF_n1559, DLX_INST_DATA_PATH_DECODE_RF_n1558, 
      DLX_INST_DATA_PATH_DECODE_RF_n1557, DLX_INST_DATA_PATH_DECODE_RF_n1556, 
      DLX_INST_DATA_PATH_DECODE_RF_n1555, DLX_INST_DATA_PATH_DECODE_RF_n1554, 
      DLX_INST_DATA_PATH_DECODE_RF_n1553, DLX_INST_DATA_PATH_DECODE_RF_n1552, 
      DLX_INST_DATA_PATH_DECODE_RF_n1551, DLX_INST_DATA_PATH_DECODE_RF_n1550, 
      DLX_INST_DATA_PATH_DECODE_RF_n1549, DLX_INST_DATA_PATH_DECODE_RF_n1548, 
      DLX_INST_DATA_PATH_DECODE_RF_n1547, DLX_INST_DATA_PATH_DECODE_RF_n1546, 
      DLX_INST_DATA_PATH_DECODE_RF_n1545, DLX_INST_DATA_PATH_DECODE_RF_n1544, 
      DLX_INST_DATA_PATH_DECODE_RF_n1543, DLX_INST_DATA_PATH_DECODE_RF_n1542, 
      DLX_INST_DATA_PATH_DECODE_RF_n1541, DLX_INST_DATA_PATH_DECODE_RF_n1540, 
      DLX_INST_DATA_PATH_DECODE_RF_n1539, DLX_INST_DATA_PATH_DECODE_RF_n1538, 
      DLX_INST_DATA_PATH_DECODE_RF_n1537, DLX_INST_DATA_PATH_DECODE_RF_n1536, 
      DLX_INST_DATA_PATH_DECODE_RF_n1535, DLX_INST_DATA_PATH_DECODE_RF_n1534, 
      DLX_INST_DATA_PATH_DECODE_RF_n1533, DLX_INST_DATA_PATH_DECODE_RF_n1532, 
      DLX_INST_DATA_PATH_DECODE_RF_n1531, DLX_INST_DATA_PATH_DECODE_RF_n1530, 
      DLX_INST_DATA_PATH_DECODE_RF_n1529, DLX_INST_DATA_PATH_DECODE_RF_n1528, 
      DLX_INST_DATA_PATH_DECODE_RF_n1527, DLX_INST_DATA_PATH_DECODE_RF_n1526, 
      DLX_INST_DATA_PATH_DECODE_RF_n1525, DLX_INST_DATA_PATH_DECODE_RF_n1524, 
      DLX_INST_DATA_PATH_DECODE_RF_n1523, DLX_INST_DATA_PATH_DECODE_RF_n1522, 
      DLX_INST_DATA_PATH_DECODE_RF_n1521, DLX_INST_DATA_PATH_DECODE_RF_n1520, 
      DLX_INST_DATA_PATH_DECODE_RF_n1519, DLX_INST_DATA_PATH_DECODE_RF_n1518, 
      DLX_INST_DATA_PATH_DECODE_RF_n1517, DLX_INST_DATA_PATH_DECODE_RF_n1516, 
      DLX_INST_DATA_PATH_DECODE_RF_n1515, DLX_INST_DATA_PATH_DECODE_RF_n1514, 
      DLX_INST_DATA_PATH_DECODE_RF_n1513, DLX_INST_DATA_PATH_DECODE_RF_n1512, 
      DLX_INST_DATA_PATH_DECODE_RF_n1511, DLX_INST_DATA_PATH_DECODE_RF_n1510, 
      DLX_INST_DATA_PATH_DECODE_RF_n1509, DLX_INST_DATA_PATH_DECODE_RF_n1508, 
      DLX_INST_DATA_PATH_DECODE_RF_n1507, DLX_INST_DATA_PATH_DECODE_RF_n1506, 
      DLX_INST_DATA_PATH_DECODE_RF_n1505, DLX_INST_DATA_PATH_DECODE_RF_n1504, 
      DLX_INST_DATA_PATH_DECODE_RF_n1503, DLX_INST_DATA_PATH_DECODE_RF_n1502, 
      DLX_INST_DATA_PATH_DECODE_RF_n1501, DLX_INST_DATA_PATH_DECODE_RF_n1500, 
      DLX_INST_DATA_PATH_DECODE_RF_n1499, DLX_INST_DATA_PATH_DECODE_RF_n1498, 
      DLX_INST_DATA_PATH_DECODE_RF_n1497, DLX_INST_DATA_PATH_DECODE_RF_n1496, 
      DLX_INST_DATA_PATH_DECODE_RF_n1495, DLX_INST_DATA_PATH_DECODE_RF_n1494, 
      DLX_INST_DATA_PATH_DECODE_RF_n1493, DLX_INST_DATA_PATH_DECODE_RF_n1492, 
      DLX_INST_DATA_PATH_DECODE_RF_n1491, DLX_INST_DATA_PATH_DECODE_RF_n1490, 
      DLX_INST_DATA_PATH_DECODE_RF_n1489, DLX_INST_DATA_PATH_DECODE_RF_n1488, 
      DLX_INST_DATA_PATH_DECODE_RF_n1487, DLX_INST_DATA_PATH_DECODE_RF_n1486, 
      DLX_INST_DATA_PATH_DECODE_RF_n1485, DLX_INST_DATA_PATH_DECODE_RF_n1484, 
      DLX_INST_DATA_PATH_DECODE_RF_n1483, DLX_INST_DATA_PATH_DECODE_RF_n1482, 
      DLX_INST_DATA_PATH_DECODE_RF_n1481, DLX_INST_DATA_PATH_DECODE_RF_n1480, 
      DLX_INST_DATA_PATH_DECODE_RF_n1479, DLX_INST_DATA_PATH_DECODE_RF_n1478, 
      DLX_INST_DATA_PATH_DECODE_RF_n1477, DLX_INST_DATA_PATH_DECODE_RF_n1476, 
      DLX_INST_DATA_PATH_DECODE_RF_n1475, DLX_INST_DATA_PATH_DECODE_RF_n1474, 
      DLX_INST_DATA_PATH_DECODE_RF_n1473, DLX_INST_DATA_PATH_DECODE_RF_n1472, 
      DLX_INST_DATA_PATH_DECODE_RF_n1471, DLX_INST_DATA_PATH_DECODE_RF_n1470, 
      DLX_INST_DATA_PATH_DECODE_RF_n1469, DLX_INST_DATA_PATH_DECODE_RF_n1468, 
      DLX_INST_DATA_PATH_DECODE_RF_n1467, DLX_INST_DATA_PATH_DECODE_RF_n1466, 
      DLX_INST_DATA_PATH_DECODE_RF_n1465, DLX_INST_DATA_PATH_DECODE_RF_n1464, 
      DLX_INST_DATA_PATH_DECODE_RF_n1463, DLX_INST_DATA_PATH_DECODE_RF_n1462, 
      DLX_INST_DATA_PATH_DECODE_RF_n1461, DLX_INST_DATA_PATH_DECODE_RF_n1460, 
      DLX_INST_DATA_PATH_DECODE_RF_n1459, DLX_INST_DATA_PATH_DECODE_RF_n1458, 
      DLX_INST_DATA_PATH_DECODE_RF_n1457, DLX_INST_DATA_PATH_DECODE_RF_n1456, 
      DLX_INST_DATA_PATH_DECODE_RF_n1455, DLX_INST_DATA_PATH_DECODE_RF_n1454, 
      DLX_INST_DATA_PATH_DECODE_RF_n1453, DLX_INST_DATA_PATH_DECODE_RF_n1452, 
      DLX_INST_DATA_PATH_DECODE_RF_n1451, DLX_INST_DATA_PATH_DECODE_RF_n1450, 
      DLX_INST_DATA_PATH_DECODE_RF_n1449, DLX_INST_DATA_PATH_DECODE_RF_n1448, 
      DLX_INST_DATA_PATH_DECODE_RF_n1447, DLX_INST_DATA_PATH_DECODE_RF_n1446, 
      DLX_INST_DATA_PATH_DECODE_RF_n1445, DLX_INST_DATA_PATH_DECODE_RF_n1444, 
      DLX_INST_DATA_PATH_DECODE_RF_n1443, DLX_INST_DATA_PATH_DECODE_RF_n1442, 
      DLX_INST_DATA_PATH_DECODE_RF_n1441, DLX_INST_DATA_PATH_DECODE_RF_n1440, 
      DLX_INST_DATA_PATH_DECODE_RF_n1439, DLX_INST_DATA_PATH_DECODE_RF_n1438, 
      DLX_INST_DATA_PATH_DECODE_RF_n1437, DLX_INST_DATA_PATH_DECODE_RF_n1436, 
      DLX_INST_DATA_PATH_DECODE_RF_n1435, DLX_INST_DATA_PATH_DECODE_RF_n1434, 
      DLX_INST_DATA_PATH_DECODE_RF_n1433, DLX_INST_DATA_PATH_DECODE_RF_n1432, 
      DLX_INST_DATA_PATH_DECODE_RF_n1431, DLX_INST_DATA_PATH_DECODE_RF_n1430, 
      DLX_INST_DATA_PATH_DECODE_RF_n1429, DLX_INST_DATA_PATH_DECODE_RF_n1428, 
      DLX_INST_DATA_PATH_DECODE_RF_n1427, DLX_INST_DATA_PATH_DECODE_RF_n1426, 
      DLX_INST_DATA_PATH_DECODE_RF_n1425, DLX_INST_DATA_PATH_DECODE_RF_n1424, 
      DLX_INST_DATA_PATH_DECODE_RF_n1423, DLX_INST_DATA_PATH_DECODE_RF_n1422, 
      DLX_INST_DATA_PATH_DECODE_RF_n1421, DLX_INST_DATA_PATH_DECODE_RF_n1420, 
      DLX_INST_DATA_PATH_DECODE_RF_n1419, DLX_INST_DATA_PATH_DECODE_RF_n1418, 
      DLX_INST_DATA_PATH_DECODE_RF_n1417, DLX_INST_DATA_PATH_DECODE_RF_n1416, 
      DLX_INST_DATA_PATH_DECODE_RF_n1415, DLX_INST_DATA_PATH_DECODE_RF_n1414, 
      DLX_INST_DATA_PATH_DECODE_RF_n1413, DLX_INST_DATA_PATH_DECODE_RF_n1412, 
      DLX_INST_DATA_PATH_DECODE_RF_n1411, DLX_INST_DATA_PATH_DECODE_RF_n1410, 
      DLX_INST_DATA_PATH_DECODE_RF_n1409, DLX_INST_DATA_PATH_DECODE_RF_n1408, 
      DLX_INST_DATA_PATH_DECODE_RF_n1407, DLX_INST_DATA_PATH_DECODE_RF_n1406, 
      DLX_INST_DATA_PATH_DECODE_RF_n1405, DLX_INST_DATA_PATH_DECODE_RF_n1404, 
      DLX_INST_DATA_PATH_DECODE_RF_n1403, DLX_INST_DATA_PATH_DECODE_RF_n1402, 
      DLX_INST_DATA_PATH_DECODE_RF_n1401, DLX_INST_DATA_PATH_DECODE_RF_n1400, 
      DLX_INST_DATA_PATH_DECODE_RF_n1399, DLX_INST_DATA_PATH_DECODE_RF_n1398, 
      DLX_INST_DATA_PATH_DECODE_RF_n1397, DLX_INST_DATA_PATH_DECODE_RF_n1396, 
      DLX_INST_DATA_PATH_DECODE_RF_n1395, DLX_INST_DATA_PATH_DECODE_RF_n1394, 
      DLX_INST_DATA_PATH_DECODE_RF_n1393, DLX_INST_DATA_PATH_DECODE_RF_n1392, 
      DLX_INST_DATA_PATH_DECODE_RF_n1391, DLX_INST_DATA_PATH_DECODE_RF_n1390, 
      DLX_INST_DATA_PATH_DECODE_RF_n1389, DLX_INST_DATA_PATH_DECODE_RF_n1388, 
      DLX_INST_DATA_PATH_DECODE_RF_n1387, DLX_INST_DATA_PATH_DECODE_RF_n1386, 
      DLX_INST_DATA_PATH_DECODE_RF_n1385, DLX_INST_DATA_PATH_DECODE_RF_n1384, 
      DLX_INST_DATA_PATH_DECODE_RF_n1383, DLX_INST_DATA_PATH_DECODE_RF_n1382, 
      DLX_INST_DATA_PATH_DECODE_RF_n1381, DLX_INST_DATA_PATH_DECODE_RF_n1380, 
      DLX_INST_DATA_PATH_DECODE_RF_n1379, DLX_INST_DATA_PATH_DECODE_RF_n1378, 
      DLX_INST_DATA_PATH_DECODE_RF_n1377, DLX_INST_DATA_PATH_DECODE_RF_n1376, 
      DLX_INST_DATA_PATH_DECODE_RF_n1375, DLX_INST_DATA_PATH_DECODE_RF_n1374, 
      DLX_INST_DATA_PATH_DECODE_RF_n1373, DLX_INST_DATA_PATH_DECODE_RF_n1372, 
      DLX_INST_DATA_PATH_DECODE_RF_n1371, DLX_INST_DATA_PATH_DECODE_RF_n1370, 
      DLX_INST_DATA_PATH_DECODE_RF_n1369, DLX_INST_DATA_PATH_DECODE_RF_n1368, 
      DLX_INST_DATA_PATH_DECODE_RF_n1367, DLX_INST_DATA_PATH_DECODE_RF_n1366, 
      DLX_INST_DATA_PATH_DECODE_RF_n1365, DLX_INST_DATA_PATH_DECODE_RF_n1364, 
      DLX_INST_DATA_PATH_DECODE_RF_n1363, DLX_INST_DATA_PATH_DECODE_RF_n1362, 
      DLX_INST_DATA_PATH_DECODE_RF_n1361, DLX_INST_DATA_PATH_DECODE_RF_n1360, 
      DLX_INST_DATA_PATH_DECODE_RF_n1359, DLX_INST_DATA_PATH_DECODE_RF_n1358, 
      DLX_INST_DATA_PATH_DECODE_RF_n1357, DLX_INST_DATA_PATH_DECODE_RF_n1356, 
      DLX_INST_DATA_PATH_DECODE_RF_n1355, DLX_INST_DATA_PATH_DECODE_RF_n1354, 
      DLX_INST_DATA_PATH_DECODE_RF_n1353, DLX_INST_DATA_PATH_DECODE_RF_n1352, 
      DLX_INST_DATA_PATH_DECODE_RF_n1351, DLX_INST_DATA_PATH_DECODE_RF_n1350, 
      DLX_INST_DATA_PATH_DECODE_RF_n1349, DLX_INST_DATA_PATH_DECODE_RF_n1348, 
      DLX_INST_DATA_PATH_DECODE_RF_n1347, DLX_INST_DATA_PATH_DECODE_RF_n1346, 
      DLX_INST_DATA_PATH_DECODE_RF_n1345, DLX_INST_DATA_PATH_DECODE_RF_n1344, 
      DLX_INST_DATA_PATH_DECODE_RF_n1343, DLX_INST_DATA_PATH_DECODE_RF_n1342, 
      DLX_INST_DATA_PATH_DECODE_RF_n1341, DLX_INST_DATA_PATH_DECODE_RF_n1340, 
      DLX_INST_DATA_PATH_DECODE_RF_n1339, DLX_INST_DATA_PATH_DECODE_RF_n1338, 
      DLX_INST_DATA_PATH_DECODE_RF_n1337, DLX_INST_DATA_PATH_DECODE_RF_n1336, 
      DLX_INST_DATA_PATH_DECODE_RF_n1335, DLX_INST_DATA_PATH_DECODE_RF_n1334, 
      DLX_INST_DATA_PATH_DECODE_RF_n1333, DLX_INST_DATA_PATH_DECODE_RF_n1332, 
      DLX_INST_DATA_PATH_DECODE_RF_n1331, DLX_INST_DATA_PATH_DECODE_RF_n1330, 
      DLX_INST_DATA_PATH_DECODE_RF_n1329, DLX_INST_DATA_PATH_DECODE_RF_n1328, 
      DLX_INST_DATA_PATH_DECODE_RF_n1327, DLX_INST_DATA_PATH_DECODE_RF_n1326, 
      DLX_INST_DATA_PATH_DECODE_RF_n1325, DLX_INST_DATA_PATH_DECODE_RF_n1324, 
      DLX_INST_DATA_PATH_DECODE_RF_n1323, DLX_INST_DATA_PATH_DECODE_RF_n1322, 
      DLX_INST_DATA_PATH_DECODE_RF_n1321, DLX_INST_DATA_PATH_DECODE_RF_n1320, 
      DLX_INST_DATA_PATH_DECODE_RF_n1319, DLX_INST_DATA_PATH_DECODE_RF_n1318, 
      DLX_INST_DATA_PATH_DECODE_RF_n1317, DLX_INST_DATA_PATH_DECODE_RF_n1316, 
      DLX_INST_DATA_PATH_DECODE_RF_n1315, DLX_INST_DATA_PATH_DECODE_RF_n1314, 
      DLX_INST_DATA_PATH_DECODE_RF_n1313, DLX_INST_DATA_PATH_DECODE_RF_n1312, 
      DLX_INST_DATA_PATH_DECODE_RF_n1311, DLX_INST_DATA_PATH_DECODE_RF_n1310, 
      DLX_INST_DATA_PATH_DECODE_RF_n1309, DLX_INST_DATA_PATH_DECODE_RF_n1308, 
      DLX_INST_DATA_PATH_DECODE_RF_n1307, DLX_INST_DATA_PATH_DECODE_RF_n1306, 
      DLX_INST_DATA_PATH_DECODE_RF_n1305, DLX_INST_DATA_PATH_DECODE_RF_n1304, 
      DLX_INST_DATA_PATH_DECODE_RF_n1303, DLX_INST_DATA_PATH_EXECUTE_n4, 
      DLX_INST_DATA_PATH_EXECUTE_n3, DLX_INST_DATA_PATH_EXECUTE_XNOR_OUT, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_0_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_1_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_2_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_3_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_4_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_5_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_6_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_7_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_8_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_9_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_10_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_11_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_12_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_13_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_14_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_15_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_16_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_17_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_18_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_19_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_20_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_21_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_22_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_23_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_24_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_25_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_26_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_27_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_28_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_29_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_30_port, 
      DLX_INST_DATA_PATH_EXECUTE_ALU_output_31_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_0_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_1_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_2_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_3_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_4_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_5_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_6_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_7_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_8_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_9_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_10_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_11_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_12_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_13_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_14_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_15_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_16_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_17_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_18_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_19_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_20_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_21_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_22_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_23_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_24_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_25_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_26_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_27_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_28_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_29_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_30_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_31_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_0_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_1_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_2_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_3_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_4_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_5_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_6_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_7_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_8_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_9_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_10_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_11_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_12_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_13_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_14_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_15_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_16_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_17_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_18_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_19_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_20_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_21_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_22_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_23_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_24_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_25_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_26_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_27_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_28_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_29_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_30_port, 
      DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_31_port, 
      DLX_INST_DATA_PATH_EXECUTE_ZERO_DEC_OUT, 
      DLX_INST_DATA_PATH_EXECUTE_Logic1_port, 
      DLX_INST_DATA_PATH_EXECUTE_zerodec_n20, 
      DLX_INST_DATA_PATH_EXECUTE_zerodec_n19, 
      DLX_INST_DATA_PATH_EXECUTE_zerodec_n18, 
      DLX_INST_DATA_PATH_EXECUTE_zerodec_n17, 
      DLX_INST_DATA_PATH_EXECUTE_zerodec_n16, 
      DLX_INST_DATA_PATH_EXECUTE_zerodec_n15, 
      DLX_INST_DATA_PATH_EXECUTE_zerodec_n14, 
      DLX_INST_DATA_PATH_EXECUTE_zerodec_n13, 
      DLX_INST_DATA_PATH_EXECUTE_zerodec_n12, 
      DLX_INST_DATA_PATH_EXECUTE_zerodec_n11, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n16, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n12, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n11, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_0_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_0_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_1_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_1_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_2_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_2_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_3_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_3_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_4_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_4_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_5_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_5_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_6_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_6_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_7_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_7_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_8_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_8_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_9_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_9_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_10_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_10_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_11_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_11_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_12_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_12_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_13_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_13_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_14_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_14_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_15_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_15_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_16_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_16_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_17_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_17_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_18_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_18_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_19_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_19_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_20_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_20_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_21_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_21_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_22_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_22_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_23_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_23_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_24_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_24_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_25_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_25_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_26_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_26_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_27_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_27_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_28_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_28_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_29_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_29_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_30_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_30_n1, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_31_n2, 
      DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_31_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_n16, DLX_INST_DATA_PATH_EXECUTE_IR3_n15, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_n14, DLX_INST_DATA_PATH_EXECUTE_IR3_n13, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_n12, DLX_INST_DATA_PATH_EXECUTE_IR3_n11, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_n10, DLX_INST_DATA_PATH_EXECUTE_IR3_n9, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_0_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_0_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_1_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_1_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_2_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_2_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_3_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_3_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_4_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_4_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_5_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_5_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_6_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_6_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_7_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_7_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_8_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_8_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_9_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_9_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_10_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_10_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_11_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_11_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_12_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_12_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_13_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_13_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_14_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_14_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_15_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_15_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_16_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_16_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_17_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_17_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_18_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_18_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_19_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_19_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_20_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_20_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_21_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_21_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_22_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_22_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_23_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_23_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_24_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_24_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_25_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_25_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_26_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_26_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_27_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_27_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_28_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_28_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_29_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_29_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_30_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_30_n1, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_31_n2, 
      DLX_INST_DATA_PATH_EXECUTE_IR3_FF_31_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_n16, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_n12, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_n11, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_0_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_0_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_1_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_1_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_2_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_2_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_3_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_3_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_4_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_4_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_5_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_5_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_6_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_6_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_7_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_7_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_8_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_8_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_9_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_9_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_10_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_10_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_11_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_11_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_12_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_12_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_13_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_13_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_14_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_14_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_15_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_15_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_16_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_16_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_17_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_17_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_18_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_18_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_19_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_19_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_20_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_20_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_21_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_21_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_22_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_22_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_23_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_23_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_24_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_24_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_25_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_25_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_26_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_26_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_27_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_27_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_28_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_28_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_29_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_29_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_30_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_30_n1, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_31_n2, 
      DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_31_n1, 
      DLX_INST_DATA_PATH_EXECUTE_COND_n4, DLX_INST_DATA_PATH_EXECUTE_COND_n3, 
      DLX_INST_DATA_PATH_MEMORY_n4, DLX_INST_DATA_PATH_MEMORY_n3, 
      DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, 
      DLX_INST_DATA_PATH_MEMORY_Logic0_port, 
      DLX_INST_DATA_PATH_MEMORY_Logic1_port, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n16, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n12, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n11, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_0_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_0_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_1_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_1_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_2_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_2_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_3_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_3_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_4_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_4_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_5_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_5_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_6_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_6_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_7_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_7_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_8_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_8_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_9_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_9_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_10_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_10_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_11_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_11_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_12_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_12_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_13_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_13_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_14_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_14_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_15_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_15_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_16_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_16_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_17_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_17_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_18_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_18_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_19_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_19_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_20_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_20_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_21_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_21_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_22_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_22_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_23_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_23_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_24_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_24_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_25_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_25_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_26_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_26_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_27_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_27_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_28_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_28_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_29_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_29_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_30_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_30_n1, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_31_n2, 
      DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_31_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_n16, DLX_INST_DATA_PATH_MEMORY_IR4_n15, 
      DLX_INST_DATA_PATH_MEMORY_IR4_n14, DLX_INST_DATA_PATH_MEMORY_IR4_n13, 
      DLX_INST_DATA_PATH_MEMORY_IR4_n12, DLX_INST_DATA_PATH_MEMORY_IR4_n11, 
      DLX_INST_DATA_PATH_MEMORY_IR4_n10, DLX_INST_DATA_PATH_MEMORY_IR4_n9, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_0_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_0_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_1_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_1_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_2_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_2_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_3_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_3_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_4_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_4_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_5_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_5_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_6_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_6_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_7_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_7_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_8_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_8_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_9_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_9_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_10_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_10_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_11_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_11_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_12_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_12_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_13_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_13_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_14_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_14_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_15_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_15_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_16_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_16_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_17_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_17_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_18_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_18_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_19_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_19_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_20_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_20_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_21_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_21_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_22_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_22_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_23_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_23_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_24_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_24_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_25_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_25_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_26_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_26_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_27_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_27_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_28_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_28_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_29_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_29_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_30_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_30_n1, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_31_n2, 
      DLX_INST_DATA_PATH_MEMORY_IR4_FF_31_n1, n_1000, n_1001, n_1002, n_1003, 
      n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, 
      n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, 
      n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, 
      n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, 
      n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, 
      n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, 
      n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, 
      n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, 
      n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, 
      n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, 
      n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, 
      n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, 
      n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, 
      n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, 
      n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, 
      n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, 
      n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, 
      n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, 
      n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, 
      n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, 
      n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, 
      n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, 
      n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, 
      n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, 
      n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, 
      n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, 
      n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, 
      n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, 
      n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, 
      n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, 
      n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, 
      n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, 
      n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, 
      n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, 
      n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, 
      n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, 
      n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, 
      n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, 
      n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, 
      n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, 
      n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, 
      n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, 
      n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, 
      n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, 
      n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, 
      n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, 
      n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, 
      n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, 
      n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, 
      n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, 
      n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, 
      n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, 
      n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, 
      n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, 
      n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, 
      n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, 
      n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, 
      n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, 
      n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, 
      n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, 
      n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, 
      n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, 
      n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, 
      n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, 
      n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, 
      n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, 
      n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, 
      n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, 
      n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, 
      n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, 
      n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, 
      n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, 
      n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, 
      n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, 
      n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, 
      n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, 
      n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, 
      n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, 
      n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, 
      n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, 
      n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, 
      n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, 
      n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, 
      n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, 
      n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, 
      n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, 
      n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, 
      n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, 
      n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, 
      n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, 
      n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, 
      n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, 
      n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, 
      n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, 
      n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, 
      n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, 
      n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, 
      n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, 
      n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, 
      n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, 
      n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, 
      n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, 
      n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, 
      n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, 
      n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, 
      n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, 
      n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, 
      n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, 
      n_1994, n_1995, n_1996 : std_logic;

begin
   
   I_RAM : IRAM port map( Rst => Rst_port_top, Addr(31) => 
                           ADDRESS_IRAM_signal_31_port, Addr(30) => 
                           ADDRESS_IRAM_signal_30_port, Addr(29) => 
                           ADDRESS_IRAM_signal_29_port, Addr(28) => 
                           ADDRESS_IRAM_signal_28_port, Addr(27) => 
                           ADDRESS_IRAM_signal_27_port, Addr(26) => 
                           ADDRESS_IRAM_signal_26_port, Addr(25) => 
                           ADDRESS_IRAM_signal_25_port, Addr(24) => 
                           ADDRESS_IRAM_signal_24_port, Addr(23) => 
                           ADDRESS_IRAM_signal_23_port, Addr(22) => 
                           ADDRESS_IRAM_signal_22_port, Addr(21) => 
                           ADDRESS_IRAM_signal_21_port, Addr(20) => 
                           ADDRESS_IRAM_signal_20_port, Addr(19) => 
                           ADDRESS_IRAM_signal_19_port, Addr(18) => 
                           ADDRESS_IRAM_signal_18_port, Addr(17) => 
                           ADDRESS_IRAM_signal_17_port, Addr(16) => 
                           ADDRESS_IRAM_signal_16_port, Addr(15) => 
                           ADDRESS_IRAM_signal_15_port, Addr(14) => 
                           ADDRESS_IRAM_signal_14_port, Addr(13) => 
                           ADDRESS_IRAM_signal_13_port, Addr(12) => 
                           ADDRESS_IRAM_signal_12_port, Addr(11) => 
                           ADDRESS_IRAM_signal_11_port, Addr(10) => 
                           ADDRESS_IRAM_signal_10_port, Addr(9) => 
                           ADDRESS_IRAM_signal_9_port, Addr(8) => 
                           ADDRESS_IRAM_signal_8_port, Addr(7) => 
                           ADDRESS_IRAM_signal_7_port, Addr(6) => 
                           ADDRESS_IRAM_signal_6_port, Addr(5) => 
                           ADDRESS_IRAM_signal_5_port, Addr(4) => 
                           ADDRESS_IRAM_signal_4_port, Addr(3) => 
                           ADDRESS_IRAM_signal_3_port, Addr(2) => 
                           ADDRESS_IRAM_signal_2_port, Addr(1) => 
                           ADDRESS_IRAM_signal_1_port, Addr(0) => 
                           ADDRESS_IRAM_signal_0_port, Dout(31) => 
                           DATA_IRAM_signal_31_port, Dout(30) => 
                           DATA_IRAM_signal_30_port, Dout(29) => 
                           DATA_IRAM_signal_29_port, Dout(28) => 
                           DATA_IRAM_signal_28_port, Dout(27) => 
                           DATA_IRAM_signal_27_port, Dout(26) => 
                           DATA_IRAM_signal_26_port, Dout(25) => 
                           DATA_IRAM_signal_25_port, Dout(24) => 
                           DATA_IRAM_signal_24_port, Dout(23) => 
                           DATA_IRAM_signal_23_port, Dout(22) => 
                           DATA_IRAM_signal_22_port, Dout(21) => 
                           DATA_IRAM_signal_21_port, Dout(20) => 
                           DATA_IRAM_signal_20_port, Dout(19) => 
                           DATA_IRAM_signal_19_port, Dout(18) => 
                           DATA_IRAM_signal_18_port, Dout(17) => 
                           DATA_IRAM_signal_17_port, Dout(16) => 
                           DATA_IRAM_signal_16_port, Dout(15) => 
                           DATA_IRAM_signal_15_port, Dout(14) => 
                           DATA_IRAM_signal_14_port, Dout(13) => 
                           DATA_IRAM_signal_13_port, Dout(12) => 
                           DATA_IRAM_signal_12_port, Dout(11) => 
                           DATA_IRAM_signal_11_port, Dout(10) => 
                           DATA_IRAM_signal_10_port, Dout(9) => 
                           DATA_IRAM_signal_9_port, Dout(8) => 
                           DATA_IRAM_signal_8_port, Dout(7) => 
                           DATA_IRAM_signal_7_port, Dout(6) => 
                           DATA_IRAM_signal_6_port, Dout(5) => 
                           DATA_IRAM_signal_5_port, Dout(4) => 
                           DATA_IRAM_signal_4_port, Dout(3) => 
                           DATA_IRAM_signal_3_port, Dout(2) => 
                           DATA_IRAM_signal_2_port, Dout(1) => 
                           DATA_IRAM_signal_1_port, Dout(0) => 
                           DATA_IRAM_signal_0_port);
   D_DRAM : dram port map( clk => Clk_port_top, w_r => n1, addr(31) => 
                           ADDRESS_DRAM_signal_31_port, addr(30) => 
                           ADDRESS_DRAM_signal_30_port, addr(29) => 
                           ADDRESS_DRAM_signal_29_port, addr(28) => 
                           ADDRESS_DRAM_signal_28_port, addr(27) => 
                           ADDRESS_DRAM_signal_27_port, addr(26) => 
                           ADDRESS_DRAM_signal_26_port, addr(25) => 
                           ADDRESS_DRAM_signal_25_port, addr(24) => 
                           ADDRESS_DRAM_signal_24_port, addr(23) => 
                           ADDRESS_DRAM_signal_23_port, addr(22) => 
                           ADDRESS_DRAM_signal_22_port, addr(21) => 
                           ADDRESS_DRAM_signal_21_port, addr(20) => 
                           ADDRESS_DRAM_signal_20_port, addr(19) => 
                           ADDRESS_DRAM_signal_19_port, addr(18) => 
                           ADDRESS_DRAM_signal_18_port, addr(17) => 
                           ADDRESS_DRAM_signal_17_port, addr(16) => 
                           ADDRESS_DRAM_signal_16_port, addr(15) => 
                           ADDRESS_DRAM_signal_15_port, addr(14) => 
                           ADDRESS_DRAM_signal_14_port, addr(13) => 
                           ADDRESS_DRAM_signal_13_port, addr(12) => 
                           ADDRESS_DRAM_signal_12_port, addr(11) => 
                           ADDRESS_DRAM_signal_11_port, addr(10) => 
                           ADDRESS_DRAM_signal_10_port, addr(9) => 
                           ADDRESS_DRAM_signal_9_port, addr(8) => 
                           ADDRESS_DRAM_signal_8_port, addr(7) => 
                           ADDRESS_DRAM_signal_7_port, addr(6) => 
                           ADDRESS_DRAM_signal_6_port, addr(5) => 
                           ADDRESS_DRAM_signal_5_port, addr(4) => 
                           ADDRESS_DRAM_signal_4_port, addr(3) => 
                           ADDRESS_DRAM_signal_3_port, addr(2) => 
                           ADDRESS_DRAM_signal_2_port, addr(1) => 
                           ADDRESS_DRAM_signal_1_port, addr(0) => 
                           ADDRESS_DRAM_signal_0_port, data_in(31) => 
                           DATAwrite_DRAM_signal_31_port, data_in(30) => 
                           DATAwrite_DRAM_signal_30_port, data_in(29) => 
                           DATAwrite_DRAM_signal_29_port, data_in(28) => 
                           DATAwrite_DRAM_signal_28_port, data_in(27) => 
                           DATAwrite_DRAM_signal_27_port, data_in(26) => 
                           DATAwrite_DRAM_signal_26_port, data_in(25) => 
                           DATAwrite_DRAM_signal_25_port, data_in(24) => 
                           DATAwrite_DRAM_signal_24_port, data_in(23) => 
                           DATAwrite_DRAM_signal_23_port, data_in(22) => 
                           DATAwrite_DRAM_signal_22_port, data_in(21) => 
                           DATAwrite_DRAM_signal_21_port, data_in(20) => 
                           DATAwrite_DRAM_signal_20_port, data_in(19) => 
                           DATAwrite_DRAM_signal_19_port, data_in(18) => 
                           DATAwrite_DRAM_signal_18_port, data_in(17) => 
                           DATAwrite_DRAM_signal_17_port, data_in(16) => 
                           DATAwrite_DRAM_signal_16_port, data_in(15) => 
                           DATAwrite_DRAM_signal_15_port, data_in(14) => 
                           DATAwrite_DRAM_signal_14_port, data_in(13) => 
                           DATAwrite_DRAM_signal_13_port, data_in(12) => 
                           DATAwrite_DRAM_signal_12_port, data_in(11) => 
                           DATAwrite_DRAM_signal_11_port, data_in(10) => 
                           DATAwrite_DRAM_signal_10_port, data_in(9) => 
                           DATAwrite_DRAM_signal_9_port, data_in(8) => 
                           DATAwrite_DRAM_signal_8_port, data_in(7) => 
                           DATAwrite_DRAM_signal_7_port, data_in(6) => 
                           DATAwrite_DRAM_signal_6_port, data_in(5) => 
                           DATAwrite_DRAM_signal_5_port, data_in(4) => 
                           DATAwrite_DRAM_signal_4_port, data_in(3) => 
                           DATAwrite_DRAM_signal_3_port, data_in(2) => 
                           DATAwrite_DRAM_signal_2_port, data_in(1) => 
                           DATAwrite_DRAM_signal_1_port, data_in(0) => 
                           DATAwrite_DRAM_signal_0_port, data_out(31) => 
                           DLX_INST_DATA_PATH_LMD_OUTs_31_port, data_out(30) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_30_port, data_out(29) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_29_port, data_out(28) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_28_port, data_out(27) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_27_port, data_out(26) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_26_port, data_out(25) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_25_port, data_out(24) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_24_port, data_out(23) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_23_port, data_out(22) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_22_port, data_out(21) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_21_port, data_out(20) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_20_port, data_out(19) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_19_port, data_out(18) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_18_port, data_out(17) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_17_port, data_out(16) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_16_port, data_out(15) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_15_port, data_out(14) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_14_port, data_out(13) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_13_port, data_out(12) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_12_port, data_out(11) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_11_port, data_out(10) =>
                           DLX_INST_DATA_PATH_LMD_OUTs_10_port, data_out(9) => 
                           DLX_INST_DATA_PATH_LMD_OUTs_9_port, data_out(8) => 
                           DLX_INST_DATA_PATH_LMD_OUTs_8_port, data_out(7) => 
                           DLX_INST_DATA_PATH_LMD_OUTs_7_port, data_out(6) => 
                           DLX_INST_DATA_PATH_LMD_OUTs_6_port, data_out(5) => 
                           DLX_INST_DATA_PATH_LMD_OUTs_5_port, data_out(4) => 
                           DLX_INST_DATA_PATH_LMD_OUTs_4_port, data_out(3) => 
                           DLX_INST_DATA_PATH_LMD_OUTs_3_port, data_out(2) => 
                           DLX_INST_DATA_PATH_LMD_OUTs_2_port, data_out(1) => 
                           DLX_INST_DATA_PATH_LMD_OUTs_1_port, data_out(0) => 
                           DLX_INST_DATA_PATH_LMD_OUTs_0_port);
   n1 <= '0';
   DLX_INST_U1 : BUF_X1 port map( A => Rst_port_top, Z => DLX_INST_n2);
   DLX_INST_IR_LATCH_EN_signal <= '1';
   DLX_INST_NPC_LATCH_EN_signal <= '1';
   DLX_INST_RegA_LATCH_EN_signal <= '0';
   DLX_INST_RegB_LATCH_EN_signal <= '0';
   DLX_INST_RegIMM_LATCH_EN_signal <= '0';
   DLX_INST_MUXA_SEL_signal <= '0';
   DLX_INST_MUXB_SEL_signal <= '0';
   DLX_INST_ALU_OUTREG_EN_signal <= '0';
   DLX_INST_EQ_COND_signal <= '0';
   DLX_INST_WE_DRAM_port <= '0';
   DLX_INST_LMD_LATCH_EN_signal <= '0';
   DLX_INST_JUMP_EN_signal <= '0';
   DLX_INST_PC_LATCH_EN_signal <= '1';
   DLX_INST_WB_MUX_SEL_signal <= '0';
   DLX_INST_RF_WE_signal <= '0';
   DLX_INST_CONTROL_UNIT_U74 : NOR3_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_28_port, A2 => 
                           DLX_INST_IR_OUT_signal_31_port, A3 => 
                           DLX_INST_IR_OUT_signal_27_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n111);
   DLX_INST_CONTROL_UNIT_U73 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_26_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n95);
   DLX_INST_CONTROL_UNIT_U72 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_29_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n65);
   DLX_INST_CONTROL_UNIT_U71 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_30_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n66);
   DLX_INST_CONTROL_UNIT_U70 : NAND4_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n111, A2 => 
                           DLX_INST_CONTROL_UNIT_n95, A3 => 
                           DLX_INST_CONTROL_UNIT_n65, A4 => 
                           DLX_INST_CONTROL_UNIT_n66, ZN => 
                           DLX_INST_CONTROL_UNIT_n69);
   DLX_INST_CONTROL_UNIT_U69 : INV_X1 port map( A => DLX_INST_CONTROL_UNIT_n69,
                           ZN => DLX_INST_CONTROL_UNIT_n76);
   DLX_INST_CONTROL_UNIT_U68 : OR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_9_port, A2 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_8_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_7_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n117);
   DLX_INST_CONTROL_UNIT_U67 : NOR4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_6_port, A2 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_4_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_10_port, A4 => 
                           DLX_INST_CONTROL_UNIT_n117, ZN => 
                           DLX_INST_CONTROL_UNIT_n77);
   DLX_INST_CONTROL_UNIT_U66 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_1_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n115);
   DLX_INST_CONTROL_UNIT_U65 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_2_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n84);
   DLX_INST_CONTROL_UNIT_U64 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_5_port, B => 
                           DLX_INST_CONTROL_UNIT_n84, Z => 
                           DLX_INST_CONTROL_UNIT_n116);
   DLX_INST_CONTROL_UNIT_U63 : NOR3_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n115, A2 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_3_port, A3 => 
                           DLX_INST_CONTROL_UNIT_n116, ZN => 
                           DLX_INST_CONTROL_UNIT_n113);
   DLX_INST_CONTROL_UNIT_U62 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_3_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n68);
   DLX_INST_CONTROL_UNIT_U61 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_5_port, A2 => 
                           DLX_INST_CONTROL_UNIT_n115, ZN => 
                           DLX_INST_CONTROL_UNIT_n81);
   DLX_INST_CONTROL_UNIT_U60 : AOI21_X1 port map( B1 => 
                           DLX_INST_CONTROL_UNIT_n68, B2 => 
                           DLX_INST_CONTROL_UNIT_n84, A => 
                           DLX_INST_CONTROL_UNIT_n81, ZN => 
                           DLX_INST_CONTROL_UNIT_n114);
   DLX_INST_CONTROL_UNIT_U59 : MUX2_X1 port map( A => 
                           DLX_INST_CONTROL_UNIT_n113, B => 
                           DLX_INST_CONTROL_UNIT_n114, S => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_0_port, Z => 
                           DLX_INST_CONTROL_UNIT_n112);
   DLX_INST_CONTROL_UNIT_U58 : NAND3_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n76, A2 => 
                           DLX_INST_CONTROL_UNIT_n77, A3 => 
                           DLX_INST_CONTROL_UNIT_n112, ZN => 
                           DLX_INST_CONTROL_UNIT_n105);
   DLX_INST_CONTROL_UNIT_U57 : NAND4_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_30_port, A2 => 
                           DLX_INST_IR_OUT_signal_29_port, A3 => 
                           DLX_INST_IR_OUT_signal_26_port, A4 => 
                           DLX_INST_CONTROL_UNIT_n111, ZN => 
                           DLX_INST_CONTROL_UNIT_n75);
   DLX_INST_CONTROL_UNIT_U56 : NAND2_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_27_port, A2 => 
                           DLX_INST_CONTROL_UNIT_n95, ZN => 
                           DLX_INST_CONTROL_UNIT_n110);
   DLX_INST_CONTROL_UNIT_U55 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_27_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n100);
   DLX_INST_CONTROL_UNIT_U54 : NAND2_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_26_port, A2 => 
                           DLX_INST_CONTROL_UNIT_n100, ZN => 
                           DLX_INST_CONTROL_UNIT_n108);
   DLX_INST_CONTROL_UNIT_U53 : MUX2_X1 port map( A => 
                           DLX_INST_CONTROL_UNIT_n110, B => 
                           DLX_INST_CONTROL_UNIT_n108, S => 
                           DLX_INST_IR_OUT_signal_29_port, Z => 
                           DLX_INST_CONTROL_UNIT_n109);
   DLX_INST_CONTROL_UNIT_U52 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_28_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n96);
   DLX_INST_CONTROL_UNIT_U51 : NAND3_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n96, A2 => 
                           DLX_INST_CONTROL_UNIT_n66, A3 => 
                           DLX_INST_IR_OUT_signal_29_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n89);
   DLX_INST_CONTROL_UNIT_U50 : OAI33_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n109, A2 => 
                           DLX_INST_CONTROL_UNIT_n66, A3 => 
                           DLX_INST_CONTROL_UNIT_n96, B1 => 
                           DLX_INST_CONTROL_UNIT_n89, B2 => 
                           DLX_INST_IR_OUT_signal_26_port, B3 => 
                           DLX_INST_CONTROL_UNIT_n100, ZN => 
                           DLX_INST_CONTROL_UNIT_n107);
   DLX_INST_CONTROL_UNIT_U49 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_31_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n72);
   DLX_INST_CONTROL_UNIT_U48 : NAND4_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_28_port, A2 => 
                           DLX_INST_IR_OUT_signal_29_port, A3 => 
                           DLX_INST_CONTROL_UNIT_n66, A4 => 
                           DLX_INST_CONTROL_UNIT_n72, ZN => 
                           DLX_INST_CONTROL_UNIT_n73);
   DLX_INST_CONTROL_UNIT_U47 : INV_X1 port map( A => DLX_INST_CONTROL_UNIT_n73,
                           ZN => DLX_INST_CONTROL_UNIT_n90);
   DLX_INST_CONTROL_UNIT_U46 : INV_X1 port map( A => DLX_INST_CONTROL_UNIT_n108
                           , ZN => DLX_INST_CONTROL_UNIT_n99);
   DLX_INST_CONTROL_UNIT_U45 : AOI22_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n107, A2 => 
                           DLX_INST_CONTROL_UNIT_n72, B1 => 
                           DLX_INST_CONTROL_UNIT_n90, B2 => 
                           DLX_INST_CONTROL_UNIT_n99, ZN => 
                           DLX_INST_CONTROL_UNIT_n106);
   DLX_INST_CONTROL_UNIT_U44 : NAND3_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n105, A2 => 
                           DLX_INST_CONTROL_UNIT_n75, A3 => 
                           DLX_INST_CONTROL_UNIT_n106, ZN => 
                           DLX_INST_CONTROL_UNIT_aluOpcode_i_0_port);
   DLX_INST_CONTROL_UNIT_U43 : NAND3_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n65, A2 => 
                           DLX_INST_CONTROL_UNIT_n66, A3 => 
                           DLX_INST_IR_OUT_signal_28_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n85);
   DLX_INST_CONTROL_UNIT_U42 : OAI211_X1 port map( C1 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_1_port, C2 => 
                           DLX_INST_CONTROL_UNIT_n84, A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_5_port, B => 
                           DLX_INST_CONTROL_UNIT_n76, ZN => 
                           DLX_INST_CONTROL_UNIT_n86);
   DLX_INST_CONTROL_UNIT_U41 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_0_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n82);
   DLX_INST_CONTROL_UNIT_U40 : XOR2_X1 port map( A => DLX_INST_CONTROL_UNIT_n82
                           , B => DLX_INST_DATA_PATH_DECODE_signExtOut_3_port, 
                           Z => DLX_INST_CONTROL_UNIT_n104);
   DLX_INST_CONTROL_UNIT_U39 : AOI21_X1 port map( B1 => 
                           DLX_INST_CONTROL_UNIT_n104, B2 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_5_port, A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_2_port, ZN => 
                           DLX_INST_CONTROL_UNIT_n103);
   DLX_INST_CONTROL_UNIT_U38 : INV_X1 port map( A => DLX_INST_CONTROL_UNIT_n103
                           , ZN => DLX_INST_CONTROL_UNIT_n101);
   DLX_INST_CONTROL_UNIT_U37 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_0_port, B2 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_3_port, A => 
                           DLX_INST_CONTROL_UNIT_n81, ZN => 
                           DLX_INST_CONTROL_UNIT_n102);
   DLX_INST_CONTROL_UNIT_U36 : AND3_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n77, A2 => 
                           DLX_INST_CONTROL_UNIT_n101, A3 => 
                           DLX_INST_CONTROL_UNIT_n102, ZN => 
                           DLX_INST_CONTROL_UNIT_n91);
   DLX_INST_CONTROL_UNIT_U35 : NOR2_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n100, A2 => 
                           DLX_INST_CONTROL_UNIT_n95, ZN => 
                           DLX_INST_CONTROL_UNIT_n71);
   DLX_INST_CONTROL_UNIT_U34 : NOR2_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_29_port, A2 => 
                           DLX_INST_CONTROL_UNIT_n71, ZN => 
                           DLX_INST_CONTROL_UNIT_n98);
   DLX_INST_CONTROL_UNIT_U33 : AOI22_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n98, A2 => 
                           DLX_INST_IR_OUT_signal_27_port, B1 => 
                           DLX_INST_CONTROL_UNIT_n99, B2 => 
                           DLX_INST_CONTROL_UNIT_n96, ZN => 
                           DLX_INST_CONTROL_UNIT_n93);
   DLX_INST_CONTROL_UNIT_U32 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_26_port, B => 
                           DLX_INST_IR_OUT_signal_27_port, S => 
                           DLX_INST_IR_OUT_signal_29_port, Z => 
                           DLX_INST_CONTROL_UNIT_n97);
   DLX_INST_CONTROL_UNIT_U31 : AOI21_X1 port map( B1 => 
                           DLX_INST_CONTROL_UNIT_n95, B2 => 
                           DLX_INST_CONTROL_UNIT_n96, A => 
                           DLX_INST_CONTROL_UNIT_n97, ZN => 
                           DLX_INST_CONTROL_UNIT_n94);
   DLX_INST_CONTROL_UNIT_U30 : MUX2_X1 port map( A => DLX_INST_CONTROL_UNIT_n93
                           , B => DLX_INST_CONTROL_UNIT_n94, S => 
                           DLX_INST_IR_OUT_signal_30_port, Z => 
                           DLX_INST_CONTROL_UNIT_n92);
   DLX_INST_CONTROL_UNIT_U29 : OAI21_X1 port map( B1 => 
                           DLX_INST_CONTROL_UNIT_n91, B2 => 
                           DLX_INST_CONTROL_UNIT_n69, A => 
                           DLX_INST_CONTROL_UNIT_n92, ZN => 
                           DLX_INST_CONTROL_UNIT_n70);
   DLX_INST_CONTROL_UNIT_U28 : AOI21_X1 port map( B1 => 
                           DLX_INST_CONTROL_UNIT_n90, B2 => 
                           DLX_INST_IR_OUT_signal_27_port, A => 
                           DLX_INST_CONTROL_UNIT_n70, ZN => 
                           DLX_INST_CONTROL_UNIT_n87);
   DLX_INST_CONTROL_UNIT_U27 : INV_X1 port map( A => DLX_INST_CONTROL_UNIT_n71,
                           ZN => DLX_INST_CONTROL_UNIT_n67);
   DLX_INST_CONTROL_UNIT_U26 : AND4_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n72, A2 => 
                           DLX_INST_CONTROL_UNIT_n67, A3 => 
                           DLX_INST_CONTROL_UNIT_n89, A4 => 
                           DLX_INST_CONTROL_UNIT_n75, ZN => 
                           DLX_INST_CONTROL_UNIT_n88);
   DLX_INST_CONTROL_UNIT_U25 : NAND4_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n85, A2 => 
                           DLX_INST_CONTROL_UNIT_n86, A3 => 
                           DLX_INST_CONTROL_UNIT_n87, A4 => 
                           DLX_INST_CONTROL_UNIT_n88, ZN => 
                           DLX_INST_CONTROL_UNIT_aluOpcode_i_1_port);
   DLX_INST_CONTROL_UNIT_U24 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_5_port, A2 => 
                           DLX_INST_CONTROL_UNIT_n82, ZN => 
                           DLX_INST_CONTROL_UNIT_n83);
   DLX_INST_CONTROL_UNIT_U23 : AOI21_X1 port map( B1 => 
                           DLX_INST_CONTROL_UNIT_n81, B2 => 
                           DLX_INST_CONTROL_UNIT_n83, A => 
                           DLX_INST_CONTROL_UNIT_n84, ZN => 
                           DLX_INST_CONTROL_UNIT_n79);
   DLX_INST_CONTROL_UNIT_U22 : NOR3_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n81, A2 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_2_port, A3 => 
                           DLX_INST_CONTROL_UNIT_n82, ZN => 
                           DLX_INST_CONTROL_UNIT_n80);
   DLX_INST_CONTROL_UNIT_U21 : MUX2_X1 port map( A => DLX_INST_CONTROL_UNIT_n79
                           , B => DLX_INST_CONTROL_UNIT_n80, S => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_3_port, Z => 
                           DLX_INST_CONTROL_UNIT_n78);
   DLX_INST_CONTROL_UNIT_U20 : NAND3_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n76, A2 => 
                           DLX_INST_CONTROL_UNIT_n77, A3 => 
                           DLX_INST_CONTROL_UNIT_n78, ZN => 
                           DLX_INST_CONTROL_UNIT_n74);
   DLX_INST_CONTROL_UNIT_U19 : OAI211_X1 port map( C1 => 
                           DLX_INST_CONTROL_UNIT_n71, C2 => 
                           DLX_INST_CONTROL_UNIT_n73, A => 
                           DLX_INST_CONTROL_UNIT_n74, B => 
                           DLX_INST_CONTROL_UNIT_n75, ZN => 
                           DLX_INST_CONTROL_UNIT_aluOpcode_i_2_port);
   DLX_INST_CONTROL_UNIT_U18 : XOR2_X1 port map( A => DLX_INST_CONTROL_UNIT_n71
                           , B => DLX_INST_CONTROL_UNIT_n72, Z => 
                           DLX_INST_CONTROL_UNIT_n60);
   DLX_INST_CONTROL_UNIT_U17 : INV_X1 port map( A => DLX_INST_CONTROL_UNIT_n70,
                           ZN => DLX_INST_CONTROL_UNIT_n61);
   DLX_INST_CONTROL_UNIT_U16 : NOR2_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n68, A2 => 
                           DLX_INST_CONTROL_UNIT_n69, ZN => 
                           DLX_INST_CONTROL_UNIT_n63);
   DLX_INST_CONTROL_UNIT_U15 : OAI21_X1 port map( B1 => 
                           DLX_INST_CONTROL_UNIT_n65, B2 => 
                           DLX_INST_CONTROL_UNIT_n66, A => 
                           DLX_INST_CONTROL_UNIT_n67, ZN => 
                           DLX_INST_CONTROL_UNIT_n64);
   DLX_INST_CONTROL_UNIT_U14 : AOI22_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n63, A2 => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_2_port, B1 => 
                           DLX_INST_IR_OUT_signal_28_port, B2 => 
                           DLX_INST_CONTROL_UNIT_n64, ZN => 
                           DLX_INST_CONTROL_UNIT_n62);
   DLX_INST_CONTROL_UNIT_U13 : NAND3_X1 port map( A1 => 
                           DLX_INST_CONTROL_UNIT_n60, A2 => 
                           DLX_INST_CONTROL_UNIT_n61, A3 => 
                           DLX_INST_CONTROL_UNIT_n62, ZN => 
                           DLX_INST_CONTROL_UNIT_aluOpcode_i_3_port);
   DLX_INST_CONTROL_UNIT_U3 : INV_X1 port map( A => DLX_INST_n2, ZN => 
                           DLX_INST_CONTROL_UNIT_n59);
   DLX_INST_CONTROL_UNIT_MUXA_SEL <= '0';
   DLX_INST_CONTROL_UNIT_MUXB_SEL <= '0';
   DLX_INST_CONTROL_UNIT_ALU_OUTREG_EN <= '0';
   DLX_INST_CONTROL_UNIT_EQ_COND <= '0';
   DLX_INST_CONTROL_UNIT_DRAM_WE <= '0';
   DLX_INST_CONTROL_UNIT_LMD_LATCH_EN <= '0';
   DLX_INST_CONTROL_UNIT_JUMP_EN <= '0';
   DLX_INST_CONTROL_UNIT_WB_MUX_SEL <= '0';
   DLX_INST_CONTROL_UNIT_RF_WE <= '0';
   DLX_INST_CONTROL_UNIT_aluOpcode1_reg_0_inst : DFFR_X1 port map( D => 
                           DLX_INST_CONTROL_UNIT_aluOpcode_i_0_port, CK => 
                           Clk_port_top, RN => DLX_INST_CONTROL_UNIT_n59, Q => 
                           DLX_INST_ALU_OPCODE_signal_3_port, QN => n_1000);
   DLX_INST_CONTROL_UNIT_aluOpcode1_reg_1_inst : DFFS_X1 port map( D => 
                           DLX_INST_CONTROL_UNIT_aluOpcode_i_1_port, CK => 
                           Clk_port_top, SN => DLX_INST_CONTROL_UNIT_n59, Q => 
                           DLX_INST_ALU_OPCODE_signal_2_port, QN => n_1001);
   DLX_INST_CONTROL_UNIT_aluOpcode1_reg_2_inst : DFFR_X1 port map( D => 
                           DLX_INST_CONTROL_UNIT_aluOpcode_i_2_port, CK => 
                           Clk_port_top, RN => DLX_INST_CONTROL_UNIT_n59, Q => 
                           DLX_INST_ALU_OPCODE_signal_1_port, QN => n_1002);
   DLX_INST_CONTROL_UNIT_aluOpcode1_reg_3_inst : DFFS_X1 port map( D => 
                           DLX_INST_CONTROL_UNIT_aluOpcode_i_3_port, CK => 
                           Clk_port_top, SN => DLX_INST_CONTROL_UNIT_n59, Q => 
                           DLX_INST_ALU_OPCODE_signal_0_port, QN => n_1003);
   DLX_INST_CONTROL_UNIT_net1651 <= '0';
   DLX_INST_CONTROL_UNIT_net1650 <= '0';
   DLX_INST_CONTROL_UNIT_net1649 <= '0';
   DLX_INST_CONTROL_UNIT_Logic1_port <= '1';
   DLX_INST_DATA_PATH_U2 : BUF_X1 port map( A => Clk_port_top, Z => 
                           DLX_INST_DATA_PATH_n4);
   DLX_INST_DATA_PATH_U1 : BUF_X1 port map( A => DLX_INST_n2, Z => 
                           DLX_INST_DATA_PATH_n3);
   DLX_INST_DATA_PATH_FETCH_U4 : BUF_X1 port map( A => DLX_INST_DATA_PATH_n4, Z
                           => DLX_INST_DATA_PATH_FETCH_n4);
   DLX_INST_DATA_PATH_FETCH_U3 : BUF_X1 port map( A => DLX_INST_DATA_PATH_n3, Z
                           => DLX_INST_DATA_PATH_FETCH_n3);
   DLX_INST_DATA_PATH_FETCH_Logic0_port <= '0';
   DLX_INST_DATA_PATH_FETCH_Logic1_port <= '1';
   DLX_INST_DATA_PATH_FETCH_ADD_U206 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_29_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n277);
   DLX_INST_DATA_PATH_FETCH_ADD_U205 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_20_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n236);
   DLX_INST_DATA_PATH_FETCH_ADD_U204 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_18_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n246);
   DLX_INST_DATA_PATH_FETCH_ADD_U203 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_14_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n312);
   DLX_INST_DATA_PATH_FETCH_ADD_U202 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_12_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n317);
   DLX_INST_DATA_PATH_FETCH_ADD_U201 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_9_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n324);
   DLX_INST_DATA_PATH_FETCH_ADD_U200 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_Logic1_port, A2 => 
                           ADDRESS_IRAM_signal_0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n240);
   DLX_INST_DATA_PATH_FETCH_ADD_U199 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n240, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n344);
   DLX_INST_DATA_PATH_FETCH_ADD_U198 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n344, B2 => 
                           ADDRESS_IRAM_signal_1_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n346);
   DLX_INST_DATA_PATH_FETCH_ADD_U197 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n346, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n345);
   DLX_INST_DATA_PATH_FETCH_ADD_U196 : OAI21_X1 port map( B1 => 
                           ADDRESS_IRAM_signal_1_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n344, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n345, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n205);
   DLX_INST_DATA_PATH_FETCH_ADD_U195 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n205, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n341);
   DLX_INST_DATA_PATH_FETCH_ADD_U194 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n341, B2 => 
                           ADDRESS_IRAM_signal_2_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n343);
   DLX_INST_DATA_PATH_FETCH_ADD_U193 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n343, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n342);
   DLX_INST_DATA_PATH_FETCH_ADD_U192 : OAI21_X1 port map( B1 => 
                           ADDRESS_IRAM_signal_2_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n341, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n342, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n195);
   DLX_INST_DATA_PATH_FETCH_ADD_U191 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n195, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n338);
   DLX_INST_DATA_PATH_FETCH_ADD_U190 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n338, B2 => 
                           ADDRESS_IRAM_signal_3_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n340);
   DLX_INST_DATA_PATH_FETCH_ADD_U189 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n340, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n339);
   DLX_INST_DATA_PATH_FETCH_ADD_U188 : OAI21_X1 port map( B1 => 
                           ADDRESS_IRAM_signal_3_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n338, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n339, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n192);
   DLX_INST_DATA_PATH_FETCH_ADD_U187 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n192, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n335);
   DLX_INST_DATA_PATH_FETCH_ADD_U186 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n335, B2 => 
                           ADDRESS_IRAM_signal_4_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n337);
   DLX_INST_DATA_PATH_FETCH_ADD_U185 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n337, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n336);
   DLX_INST_DATA_PATH_FETCH_ADD_U184 : OAI21_X1 port map( B1 => 
                           ADDRESS_IRAM_signal_4_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n335, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n336, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n332);
   DLX_INST_DATA_PATH_FETCH_ADD_U183 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_5_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n333);
   DLX_INST_DATA_PATH_FETCH_ADD_U182 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n332, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n189);
   DLX_INST_DATA_PATH_FETCH_ADD_U181 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n189, B2 => 
                           ADDRESS_IRAM_signal_5_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n334);
   DLX_INST_DATA_PATH_FETCH_ADD_U180 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n332, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n333, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n334, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n186);
   DLX_INST_DATA_PATH_FETCH_ADD_U179 : AND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n186, A2 => 
                           ADDRESS_IRAM_signal_6_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n331);
   DLX_INST_DATA_PATH_FETCH_ADD_U178 : OAI22_X1 port map( A1 => 
                           ADDRESS_IRAM_signal_6_port, A2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n186, B1 => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n331, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n183);
   DLX_INST_DATA_PATH_FETCH_ADD_U177 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_7_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n328);
   DLX_INST_DATA_PATH_FETCH_ADD_U176 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n183, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n330);
   DLX_INST_DATA_PATH_FETCH_ADD_U175 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n330, B2 => 
                           ADDRESS_IRAM_signal_7_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n329);
   DLX_INST_DATA_PATH_FETCH_ADD_U174 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n183, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n328, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n329, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n180);
   DLX_INST_DATA_PATH_FETCH_ADD_U173 : AND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n180, A2 => 
                           ADDRESS_IRAM_signal_8_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n327);
   DLX_INST_DATA_PATH_FETCH_ADD_U172 : OAI22_X1 port map( A1 => 
                           ADDRESS_IRAM_signal_8_port, A2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n180, B1 => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n327, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n177);
   DLX_INST_DATA_PATH_FETCH_ADD_U171 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n177, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n326);
   DLX_INST_DATA_PATH_FETCH_ADD_U170 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n326, B2 => 
                           ADDRESS_IRAM_signal_9_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n325);
   DLX_INST_DATA_PATH_FETCH_ADD_U169 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n324, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n177, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n325, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n271);
   DLX_INST_DATA_PATH_FETCH_ADD_U168 : AND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n271, A2 => 
                           ADDRESS_IRAM_signal_10_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n323);
   DLX_INST_DATA_PATH_FETCH_ADD_U167 : OAI22_X1 port map( A1 => 
                           ADDRESS_IRAM_signal_10_port, A2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n271, B1 => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n323, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n268);
   DLX_INST_DATA_PATH_FETCH_ADD_U166 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_11_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n320);
   DLX_INST_DATA_PATH_FETCH_ADD_U165 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n268, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n322);
   DLX_INST_DATA_PATH_FETCH_ADD_U164 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n322, B2 => 
                           ADDRESS_IRAM_signal_11_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n321);
   DLX_INST_DATA_PATH_FETCH_ADD_U163 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n268, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n320, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n321, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n319);
   DLX_INST_DATA_PATH_FETCH_ADD_U162 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n319, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n265);
   DLX_INST_DATA_PATH_FETCH_ADD_U161 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n319, B2 => 
                           ADDRESS_IRAM_signal_12_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n318);
   DLX_INST_DATA_PATH_FETCH_ADD_U160 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n317, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n265, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n318, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n262);
   DLX_INST_DATA_PATH_FETCH_ADD_U159 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n262, B2 => 
                           ADDRESS_IRAM_signal_13_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n316);
   DLX_INST_DATA_PATH_FETCH_ADD_U158 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n316, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n315);
   DLX_INST_DATA_PATH_FETCH_ADD_U157 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n262, B2 => 
                           ADDRESS_IRAM_signal_13_port, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n315, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n259);
   DLX_INST_DATA_PATH_FETCH_ADD_U156 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n259, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n314);
   DLX_INST_DATA_PATH_FETCH_ADD_U155 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n314, B2 => 
                           ADDRESS_IRAM_signal_14_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n313);
   DLX_INST_DATA_PATH_FETCH_ADD_U154 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n312, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n259, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n313, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n256);
   DLX_INST_DATA_PATH_FETCH_ADD_U153 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n256, B2 => 
                           ADDRESS_IRAM_signal_15_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n311);
   DLX_INST_DATA_PATH_FETCH_ADD_U152 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n311, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n310);
   DLX_INST_DATA_PATH_FETCH_ADD_U151 : OAI21_X1 port map( B1 => 
                           ADDRESS_IRAM_signal_15_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n256, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n310, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n253);
   DLX_INST_DATA_PATH_FETCH_ADD_U150 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_16_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n307);
   DLX_INST_DATA_PATH_FETCH_ADD_U149 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n253, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n309);
   DLX_INST_DATA_PATH_FETCH_ADD_U148 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n309, B2 => 
                           ADDRESS_IRAM_signal_16_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n308);
   DLX_INST_DATA_PATH_FETCH_ADD_U147 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n253, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n307, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n308, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n250);
   DLX_INST_DATA_PATH_FETCH_ADD_U146 : OAI21_X1 port map( B1 => 
                           ADDRESS_IRAM_signal_17_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n250, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n306);
   DLX_INST_DATA_PATH_FETCH_ADD_U145 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n306, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n305);
   DLX_INST_DATA_PATH_FETCH_ADD_U144 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n250, B2 => 
                           ADDRESS_IRAM_signal_17_port, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n305, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n303);
   DLX_INST_DATA_PATH_FETCH_ADD_U143 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n303, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n247);
   DLX_INST_DATA_PATH_FETCH_ADD_U142 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n247, B2 => 
                           ADDRESS_IRAM_signal_18_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n304);
   DLX_INST_DATA_PATH_FETCH_ADD_U141 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n246, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n303, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n304, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n243);
   DLX_INST_DATA_PATH_FETCH_ADD_U140 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n243, B2 => 
                           ADDRESS_IRAM_signal_19_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n302);
   DLX_INST_DATA_PATH_FETCH_ADD_U139 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n302, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n301);
   DLX_INST_DATA_PATH_FETCH_ADD_U138 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n243, B2 => 
                           ADDRESS_IRAM_signal_19_port, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n301, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n299);
   DLX_INST_DATA_PATH_FETCH_ADD_U137 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n299, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n237);
   DLX_INST_DATA_PATH_FETCH_ADD_U136 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n237, B2 => 
                           ADDRESS_IRAM_signal_20_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n300);
   DLX_INST_DATA_PATH_FETCH_ADD_U135 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n236, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n299, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n300, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n233);
   DLX_INST_DATA_PATH_FETCH_ADD_U134 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n233, B2 => 
                           ADDRESS_IRAM_signal_21_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n298);
   DLX_INST_DATA_PATH_FETCH_ADD_U133 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n298, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n297);
   DLX_INST_DATA_PATH_FETCH_ADD_U132 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n233, B2 => 
                           ADDRESS_IRAM_signal_21_port, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n297, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n295);
   DLX_INST_DATA_PATH_FETCH_ADD_U131 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_22_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n229);
   DLX_INST_DATA_PATH_FETCH_ADD_U130 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n295, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n230);
   DLX_INST_DATA_PATH_FETCH_ADD_U129 : OAI21_X1 port map( B1 => 
                           ADDRESS_IRAM_signal_22_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n230, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n296);
   DLX_INST_DATA_PATH_FETCH_ADD_U128 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n295, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n229, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n296, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n226);
   DLX_INST_DATA_PATH_FETCH_ADD_U127 : OR2_X1 port map( A1 => 
                           ADDRESS_IRAM_signal_23_port, A2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n226, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n294);
   DLX_INST_DATA_PATH_FETCH_ADD_U126 : AOI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n226, A2 => 
                           ADDRESS_IRAM_signal_23_port, B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n294, B2 => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n293);
   DLX_INST_DATA_PATH_FETCH_ADD_U125 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n293, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n223);
   DLX_INST_DATA_PATH_FETCH_ADD_U124 : OR2_X1 port map( A1 => 
                           ADDRESS_IRAM_signal_24_port, A2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n223, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n292);
   DLX_INST_DATA_PATH_FETCH_ADD_U123 : AOI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n223, A2 => 
                           ADDRESS_IRAM_signal_24_port, B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n292, B2 => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n289);
   DLX_INST_DATA_PATH_FETCH_ADD_U122 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_25_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n290);
   DLX_INST_DATA_PATH_FETCH_ADD_U121 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n289, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n220);
   DLX_INST_DATA_PATH_FETCH_ADD_U120 : OAI21_X1 port map( B1 => 
                           ADDRESS_IRAM_signal_25_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n220, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n291);
   DLX_INST_DATA_PATH_FETCH_ADD_U119 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n289, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n290, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n291, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n217);
   DLX_INST_DATA_PATH_FETCH_ADD_U118 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n217, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n286);
   DLX_INST_DATA_PATH_FETCH_ADD_U117 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_26_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n287);
   DLX_INST_DATA_PATH_FETCH_ADD_U116 : OAI21_X1 port map( B1 => 
                           ADDRESS_IRAM_signal_26_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n217, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n288);
   DLX_INST_DATA_PATH_FETCH_ADD_U115 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n286, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n287, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n288, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n214);
   DLX_INST_DATA_PATH_FETCH_ADD_U114 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n214, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n283);
   DLX_INST_DATA_PATH_FETCH_ADD_U113 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_27_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n284);
   DLX_INST_DATA_PATH_FETCH_ADD_U112 : OAI21_X1 port map( B1 => 
                           ADDRESS_IRAM_signal_27_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n214, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n285);
   DLX_INST_DATA_PATH_FETCH_ADD_U111 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n283, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n284, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n285, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n211);
   DLX_INST_DATA_PATH_FETCH_ADD_U110 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n211, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n280);
   DLX_INST_DATA_PATH_FETCH_ADD_U109 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_28_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n281);
   DLX_INST_DATA_PATH_FETCH_ADD_U108 : OAI21_X1 port map( B1 => 
                           ADDRESS_IRAM_signal_28_port, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n211, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n282);
   DLX_INST_DATA_PATH_FETCH_ADD_U107 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n280, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n281, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n282, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n208);
   DLX_INST_DATA_PATH_FETCH_ADD_U106 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n208, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n278);
   DLX_INST_DATA_PATH_FETCH_ADD_U105 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n208, B2 => 
                           ADDRESS_IRAM_signal_29_port, A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n279);
   DLX_INST_DATA_PATH_FETCH_ADD_U104 : AOI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n277, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n278, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n279, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n202);
   DLX_INST_DATA_PATH_FETCH_ADD_U103 : OR2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n202, A2 => 
                           ADDRESS_IRAM_signal_30_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n276);
   DLX_INST_DATA_PATH_FETCH_ADD_U102 : AOI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n202, A2 => 
                           ADDRESS_IRAM_signal_30_port, B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n276, B2 => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n198);
   DLX_INST_DATA_PATH_FETCH_ADD_U101 : INV_X1 port map( A => 
                           ADDRESS_IRAM_signal_31_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n199);
   DLX_INST_DATA_PATH_FETCH_ADD_U100 : AND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n199, A2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n198, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n274);
   DLX_INST_DATA_PATH_FETCH_ADD_U99 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n275);
   DLX_INST_DATA_PATH_FETCH_ADD_U98 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n198, A2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n199, B1 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n274, B2 => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n275, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_Co);
   DLX_INST_DATA_PATH_FETCH_ADD_U97 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic1_port, B => 
                           ADDRESS_IRAM_signal_0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n272);
   DLX_INST_DATA_PATH_FETCH_ADD_U96 : OAI21_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_FETCH_Logic1_port, B2 => 
                           ADDRESS_IRAM_signal_0_port, A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n240, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n273);
   DLX_INST_DATA_PATH_FETCH_ADD_U95 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n272, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n273, S => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_0_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U94 : XOR2_X1 port map( A => 
                           ADDRESS_IRAM_signal_10_port, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n271, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n269);
   DLX_INST_DATA_PATH_FETCH_ADD_U93 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n270);
   DLX_INST_DATA_PATH_FETCH_ADD_U92 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n269, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n270, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_10_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U91 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n266);
   DLX_INST_DATA_PATH_FETCH_ADD_U90 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n268, B => 
                           ADDRESS_IRAM_signal_11_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n267);
   DLX_INST_DATA_PATH_FETCH_ADD_U89 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n266, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n267, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_11_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U88 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n263);
   DLX_INST_DATA_PATH_FETCH_ADD_U87 : XOR2_X1 port map( A => 
                           ADDRESS_IRAM_signal_12_port, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n265, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n264);
   DLX_INST_DATA_PATH_FETCH_ADD_U86 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n263, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n264, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_12_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U85 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n260);
   DLX_INST_DATA_PATH_FETCH_ADD_U84 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n262, B => 
                           ADDRESS_IRAM_signal_13_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n261);
   DLX_INST_DATA_PATH_FETCH_ADD_U83 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n260, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n261, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_13_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U82 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n257);
   DLX_INST_DATA_PATH_FETCH_ADD_U81 : XOR2_X1 port map( A => 
                           ADDRESS_IRAM_signal_14_port, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n259, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n258);
   DLX_INST_DATA_PATH_FETCH_ADD_U80 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n257, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n258, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_14_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U79 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n254);
   DLX_INST_DATA_PATH_FETCH_ADD_U78 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n256, B => 
                           ADDRESS_IRAM_signal_15_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n255);
   DLX_INST_DATA_PATH_FETCH_ADD_U77 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n254, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n255, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_15_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U76 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n251);
   DLX_INST_DATA_PATH_FETCH_ADD_U75 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n253, B => 
                           ADDRESS_IRAM_signal_16_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n252);
   DLX_INST_DATA_PATH_FETCH_ADD_U74 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n251, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n252, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_16_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U73 : XOR2_X1 port map( A => 
                           ADDRESS_IRAM_signal_17_port, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n250, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n248);
   DLX_INST_DATA_PATH_FETCH_ADD_U72 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n249);
   DLX_INST_DATA_PATH_FETCH_ADD_U71 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n248, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n249, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_17_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U70 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n244);
   DLX_INST_DATA_PATH_FETCH_ADD_U69 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n246, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n247, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n245);
   DLX_INST_DATA_PATH_FETCH_ADD_U68 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n244, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n245, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_18_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U67 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n241);
   DLX_INST_DATA_PATH_FETCH_ADD_U66 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n243, B => 
                           ADDRESS_IRAM_signal_19_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n242);
   DLX_INST_DATA_PATH_FETCH_ADD_U65 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n241, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n242, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_19_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U64 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n238);
   DLX_INST_DATA_PATH_FETCH_ADD_U63 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n240, B => 
                           ADDRESS_IRAM_signal_1_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n239);
   DLX_INST_DATA_PATH_FETCH_ADD_U62 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n238, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n239, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_1_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U61 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n234);
   DLX_INST_DATA_PATH_FETCH_ADD_U60 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n236, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n237, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n235);
   DLX_INST_DATA_PATH_FETCH_ADD_U59 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n234, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n235, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_20_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U58 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n231);
   DLX_INST_DATA_PATH_FETCH_ADD_U57 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n233, B => 
                           ADDRESS_IRAM_signal_21_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n232);
   DLX_INST_DATA_PATH_FETCH_ADD_U56 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n231, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n232, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_21_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U55 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n227);
   DLX_INST_DATA_PATH_FETCH_ADD_U54 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n229, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n230, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n228);
   DLX_INST_DATA_PATH_FETCH_ADD_U53 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n227, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n228, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_22_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U52 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n226, B => 
                           ADDRESS_IRAM_signal_23_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n224);
   DLX_INST_DATA_PATH_FETCH_ADD_U51 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n225);
   DLX_INST_DATA_PATH_FETCH_ADD_U50 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n224, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n225, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_23_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U49 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n223, B => 
                           ADDRESS_IRAM_signal_24_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n221);
   DLX_INST_DATA_PATH_FETCH_ADD_U48 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n222);
   DLX_INST_DATA_PATH_FETCH_ADD_U47 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n221, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n222, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_24_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U46 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n220, B => 
                           ADDRESS_IRAM_signal_25_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n218);
   DLX_INST_DATA_PATH_FETCH_ADD_U45 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n219);
   DLX_INST_DATA_PATH_FETCH_ADD_U44 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n218, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n219, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_25_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U43 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n217, B => 
                           ADDRESS_IRAM_signal_26_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n215);
   DLX_INST_DATA_PATH_FETCH_ADD_U42 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n216);
   DLX_INST_DATA_PATH_FETCH_ADD_U41 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n215, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n216, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_26_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U40 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n214, B => 
                           ADDRESS_IRAM_signal_27_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n212);
   DLX_INST_DATA_PATH_FETCH_ADD_U39 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n213);
   DLX_INST_DATA_PATH_FETCH_ADD_U38 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n212, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n213, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_27_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U37 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n211, B => 
                           ADDRESS_IRAM_signal_28_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n209);
   DLX_INST_DATA_PATH_FETCH_ADD_U36 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n210);
   DLX_INST_DATA_PATH_FETCH_ADD_U35 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n209, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n210, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_28_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U34 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n208, B => 
                           ADDRESS_IRAM_signal_29_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n206);
   DLX_INST_DATA_PATH_FETCH_ADD_U33 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n207);
   DLX_INST_DATA_PATH_FETCH_ADD_U32 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n206, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n207, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_29_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U31 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n203);
   DLX_INST_DATA_PATH_FETCH_ADD_U30 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n205, B => 
                           ADDRESS_IRAM_signal_2_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n204);
   DLX_INST_DATA_PATH_FETCH_ADD_U29 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n203, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n204, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_2_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U28 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n200);
   DLX_INST_DATA_PATH_FETCH_ADD_U27 : XOR2_X1 port map( A => 
                           ADDRESS_IRAM_signal_30_port, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n202, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n201);
   DLX_INST_DATA_PATH_FETCH_ADD_U26 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n200, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n201, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_30_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U25 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n198, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n199, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n196);
   DLX_INST_DATA_PATH_FETCH_ADD_U24 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n197);
   DLX_INST_DATA_PATH_FETCH_ADD_U23 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n196, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n197, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_31_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U22 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n193);
   DLX_INST_DATA_PATH_FETCH_ADD_U21 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n195, B => 
                           ADDRESS_IRAM_signal_3_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n194);
   DLX_INST_DATA_PATH_FETCH_ADD_U20 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n193, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n194, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_3_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U19 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n190);
   DLX_INST_DATA_PATH_FETCH_ADD_U18 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n192, B => 
                           ADDRESS_IRAM_signal_4_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n191);
   DLX_INST_DATA_PATH_FETCH_ADD_U17 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n190, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n191, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_4_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U16 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n187);
   DLX_INST_DATA_PATH_FETCH_ADD_U15 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n189, B => 
                           ADDRESS_IRAM_signal_5_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n188);
   DLX_INST_DATA_PATH_FETCH_ADD_U14 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n187, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n188, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_5_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U13 : XOR2_X1 port map( A => 
                           ADDRESS_IRAM_signal_6_port, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n186, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n184);
   DLX_INST_DATA_PATH_FETCH_ADD_U12 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n185);
   DLX_INST_DATA_PATH_FETCH_ADD_U11 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n184, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n185, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_6_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U10 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n181);
   DLX_INST_DATA_PATH_FETCH_ADD_U9 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n183, B => 
                           ADDRESS_IRAM_signal_7_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n182);
   DLX_INST_DATA_PATH_FETCH_ADD_U8 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n181, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n182, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_7_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U7 : XOR2_X1 port map( A => 
                           ADDRESS_IRAM_signal_8_port, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n180, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n178);
   DLX_INST_DATA_PATH_FETCH_ADD_U6 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n179);
   DLX_INST_DATA_PATH_FETCH_ADD_U5 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n178, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n179, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_8_port);
   DLX_INST_DATA_PATH_FETCH_ADD_U4 : XNOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, B => 
                           DLX_INST_DATA_PATH_FETCH_Logic0_port, ZN => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n175);
   DLX_INST_DATA_PATH_FETCH_ADD_U3 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n177, B => 
                           ADDRESS_IRAM_signal_9_port, Z => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n176);
   DLX_INST_DATA_PATH_FETCH_ADD_U2 : XOR2_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n175, B => 
                           DLX_INST_DATA_PATH_FETCH_ADD_n176, Z => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_9_port);
   DLX_INST_DATA_PATH_FETCH_PC_U8 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_PC_n16, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_n15);
   DLX_INST_DATA_PATH_FETCH_PC_U7 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_PC_n16, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14);
   DLX_INST_DATA_PATH_FETCH_PC_U6 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_PC_n16, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13);
   DLX_INST_DATA_PATH_FETCH_PC_U5 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_PC_n12, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_n11);
   DLX_INST_DATA_PATH_FETCH_PC_U4 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_PC_n12, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10);
   DLX_INST_DATA_PATH_FETCH_PC_U3 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_PC_n12, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9);
   DLX_INST_DATA_PATH_FETCH_PC_U2 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_n4, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_n16);
   DLX_INST_DATA_PATH_FETCH_PC_U1 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_n3, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_n12);
   DLX_INST_DATA_PATH_FETCH_PC_FF_0_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_0_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_0_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_0_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_0_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n11, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_0_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_0_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_0_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_0_n2, Q => 
                           ADDRESS_IRAM_signal_0_port, QN => n_1004);
   DLX_INST_DATA_PATH_FETCH_PC_FF_1_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_1_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_1_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_1_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_1_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_1_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_1_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_1_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_1_n2, Q => 
                           ADDRESS_IRAM_signal_1_port, QN => n_1005);
   DLX_INST_DATA_PATH_FETCH_PC_FF_2_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_2_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_2_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_2_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_2_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_2_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_2_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_2_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_2_n2, Q => 
                           ADDRESS_IRAM_signal_2_port, QN => n_1006);
   DLX_INST_DATA_PATH_FETCH_PC_FF_3_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_3_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_3_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_3_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_3_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_3_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_3_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_3_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_3_n2, Q => 
                           ADDRESS_IRAM_signal_3_port, QN => n_1007);
   DLX_INST_DATA_PATH_FETCH_PC_FF_4_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_4_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_4_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_4_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_4_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_4_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_4_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_4_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_4_n2, Q => 
                           ADDRESS_IRAM_signal_4_port, QN => n_1008);
   DLX_INST_DATA_PATH_FETCH_PC_FF_5_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_5_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_5_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_5_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_5_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_5_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_5_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_5_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_5_n2, Q => 
                           ADDRESS_IRAM_signal_5_port, QN => n_1009);
   DLX_INST_DATA_PATH_FETCH_PC_FF_6_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_6_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_6_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_6_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_6_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_6_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_6_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_6_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_6_n2, Q => 
                           ADDRESS_IRAM_signal_6_port, QN => n_1010);
   DLX_INST_DATA_PATH_FETCH_PC_FF_7_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_7_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_7_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_7_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_7_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_7_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_7_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_7_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_7_n2, Q => 
                           ADDRESS_IRAM_signal_7_port, QN => n_1011);
   DLX_INST_DATA_PATH_FETCH_PC_FF_8_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_8_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_8_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_8_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_8_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_8_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_8_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_8_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_8_n2, Q => 
                           ADDRESS_IRAM_signal_8_port, QN => n_1012);
   DLX_INST_DATA_PATH_FETCH_PC_FF_9_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_9_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_9_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_9_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_9_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_9_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_9_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_9_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_9_n2, Q => 
                           ADDRESS_IRAM_signal_9_port, QN => n_1013);
   DLX_INST_DATA_PATH_FETCH_PC_FF_10_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_10_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_10_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_10_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_10_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_10_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_10_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_10_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_10_n2, Q => 
                           ADDRESS_IRAM_signal_10_port, QN => n_1014);
   DLX_INST_DATA_PATH_FETCH_PC_FF_11_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_11_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_11_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_11_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_11_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_11_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_11_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_11_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_11_n2, Q => 
                           ADDRESS_IRAM_signal_11_port, QN => n_1015);
   DLX_INST_DATA_PATH_FETCH_PC_FF_12_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_12_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_12_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_12_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_12_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n9, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_12_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_12_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_12_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_12_n2, Q => 
                           ADDRESS_IRAM_signal_12_port, QN => n_1016);
   DLX_INST_DATA_PATH_FETCH_PC_FF_13_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_13_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_13_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_13_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_13_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_13_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_13_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_13_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_13_n2, Q => 
                           ADDRESS_IRAM_signal_13_port, QN => n_1017);
   DLX_INST_DATA_PATH_FETCH_PC_FF_14_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_14_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_14_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_14_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_14_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_14_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_14_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_14_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_14_n2, Q => 
                           ADDRESS_IRAM_signal_14_port, QN => n_1018);
   DLX_INST_DATA_PATH_FETCH_PC_FF_15_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_15_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_15_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_15_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_15_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_15_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_15_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_15_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_15_n2, Q => 
                           ADDRESS_IRAM_signal_15_port, QN => n_1019);
   DLX_INST_DATA_PATH_FETCH_PC_FF_16_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_16_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_16_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_16_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_16_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_16_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_16_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_16_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_16_n2, Q => 
                           ADDRESS_IRAM_signal_16_port, QN => n_1020);
   DLX_INST_DATA_PATH_FETCH_PC_FF_17_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_17_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_17_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_17_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_17_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_17_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_17_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_17_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_17_n2, Q => 
                           ADDRESS_IRAM_signal_17_port, QN => n_1021);
   DLX_INST_DATA_PATH_FETCH_PC_FF_18_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_18_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_18_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_18_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_18_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_18_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_18_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_18_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_18_n2, Q => 
                           ADDRESS_IRAM_signal_18_port, QN => n_1022);
   DLX_INST_DATA_PATH_FETCH_PC_FF_19_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_19_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_19_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_19_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_19_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_19_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_19_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_19_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_19_n2, Q => 
                           ADDRESS_IRAM_signal_19_port, QN => n_1023);
   DLX_INST_DATA_PATH_FETCH_PC_FF_20_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_20_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_20_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_20_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_20_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_20_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_20_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_20_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_20_n2, Q => 
                           ADDRESS_IRAM_signal_20_port, QN => n_1024);
   DLX_INST_DATA_PATH_FETCH_PC_FF_21_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_21_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_21_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_21_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_21_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_21_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_21_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_21_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_21_n2, Q => 
                           ADDRESS_IRAM_signal_21_port, QN => n_1025);
   DLX_INST_DATA_PATH_FETCH_PC_FF_22_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_22_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_22_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_22_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_22_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_22_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_22_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_22_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_22_n2, Q => 
                           ADDRESS_IRAM_signal_22_port, QN => n_1026);
   DLX_INST_DATA_PATH_FETCH_PC_FF_23_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_23_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_23_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_23_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_23_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_23_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_23_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_23_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_23_n2, Q => 
                           ADDRESS_IRAM_signal_23_port, QN => n_1027);
   DLX_INST_DATA_PATH_FETCH_PC_FF_24_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_24_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_24_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_24_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_24_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n10, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_24_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_24_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_24_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_24_n2, Q => 
                           ADDRESS_IRAM_signal_24_port, QN => n_1028);
   DLX_INST_DATA_PATH_FETCH_PC_FF_25_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_25_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_25_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_25_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_25_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n11, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_25_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_25_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_25_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_25_n2, Q => 
                           ADDRESS_IRAM_signal_25_port, QN => n_1029);
   DLX_INST_DATA_PATH_FETCH_PC_FF_26_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_26_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_26_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_26_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_26_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n11, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_26_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_26_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_26_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_26_n2, Q => 
                           ADDRESS_IRAM_signal_26_port, QN => n_1030);
   DLX_INST_DATA_PATH_FETCH_PC_FF_27_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_27_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_27_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_27_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_27_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n11, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_27_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_27_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_27_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_27_n2, Q => 
                           ADDRESS_IRAM_signal_27_port, QN => n_1031);
   DLX_INST_DATA_PATH_FETCH_PC_FF_28_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_28_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_28_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_28_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_28_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n11, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_28_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_28_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_28_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_28_n2, Q => 
                           ADDRESS_IRAM_signal_28_port, QN => n_1032);
   DLX_INST_DATA_PATH_FETCH_PC_FF_29_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_29_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_29_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_29_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_29_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n11, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_29_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_29_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_29_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_29_n2, Q => 
                           ADDRESS_IRAM_signal_29_port, QN => n_1033);
   DLX_INST_DATA_PATH_FETCH_PC_FF_30_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_30_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_30_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_30_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_30_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n11, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_30_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_30_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_30_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_30_n2, Q => 
                           ADDRESS_IRAM_signal_30_port, QN => n_1034);
   DLX_INST_DATA_PATH_FETCH_PC_FF_31_U3 : MUX2_X1 port map( A => 
                           ADDRESS_IRAM_signal_31_port, B => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_31_port, S => 
                           DLX_INST_PC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_31_n1);
   DLX_INST_DATA_PATH_FETCH_PC_FF_31_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_PC_n11, A2 => 
                           DLX_INST_PC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_31_n2);
   DLX_INST_DATA_PATH_FETCH_PC_FF_31_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_31_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_PC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_PC_FF_31_n2, Q => 
                           ADDRESS_IRAM_signal_31_port, QN => n_1035);
   DLX_INST_DATA_PATH_FETCH_IR_U8 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_IR_n16, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_n15);
   DLX_INST_DATA_PATH_FETCH_IR_U7 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_IR_n16, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14);
   DLX_INST_DATA_PATH_FETCH_IR_U6 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_IR_n16, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13);
   DLX_INST_DATA_PATH_FETCH_IR_U5 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_IR_n12, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_n11);
   DLX_INST_DATA_PATH_FETCH_IR_U4 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_IR_n12, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10);
   DLX_INST_DATA_PATH_FETCH_IR_U3 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_IR_n12, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9);
   DLX_INST_DATA_PATH_FETCH_IR_U2 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_n4, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_n16);
   DLX_INST_DATA_PATH_FETCH_IR_U1 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_n3, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_n12);
   DLX_INST_DATA_PATH_FETCH_IR_FF_0_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_0_port, B => 
                           DATA_IRAM_signal_0_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_0_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_0_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_0_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_0_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_0_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_0_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_0_port, QN => 
                           n_1036);
   DLX_INST_DATA_PATH_FETCH_IR_FF_1_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_1_port, B => 
                           DATA_IRAM_signal_1_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_1_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_1_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_1_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_1_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_1_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_1_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_1_port, QN => 
                           n_1037);
   DLX_INST_DATA_PATH_FETCH_IR_FF_2_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_2_port, B => 
                           DATA_IRAM_signal_2_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_2_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_2_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_2_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_2_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_2_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_2_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_2_port, QN => 
                           n_1038);
   DLX_INST_DATA_PATH_FETCH_IR_FF_3_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_3_port, B => 
                           DATA_IRAM_signal_3_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_3_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_3_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_3_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_3_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_3_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_3_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_3_port, QN => 
                           n_1039);
   DLX_INST_DATA_PATH_FETCH_IR_FF_4_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_4_port, B => 
                           DATA_IRAM_signal_4_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_4_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_4_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_4_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_4_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_4_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_4_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_4_port, QN => 
                           n_1040);
   DLX_INST_DATA_PATH_FETCH_IR_FF_5_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_5_port, B => 
                           DATA_IRAM_signal_5_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_5_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_5_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_5_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_5_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_5_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_5_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_5_port, QN => 
                           n_1041);
   DLX_INST_DATA_PATH_FETCH_IR_FF_6_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_6_port, B => 
                           DATA_IRAM_signal_6_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_6_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_6_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_6_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_6_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_6_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_6_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_6_port, QN => 
                           n_1042);
   DLX_INST_DATA_PATH_FETCH_IR_FF_7_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_7_port, B => 
                           DATA_IRAM_signal_7_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_7_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_7_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_7_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_7_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_7_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_7_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_7_port, QN => 
                           n_1043);
   DLX_INST_DATA_PATH_FETCH_IR_FF_8_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_8_port, B => 
                           DATA_IRAM_signal_8_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_8_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_8_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_8_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_8_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_8_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_8_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_8_port, QN => 
                           n_1044);
   DLX_INST_DATA_PATH_FETCH_IR_FF_9_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_9_port, B => 
                           DATA_IRAM_signal_9_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_9_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_9_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_9_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_9_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_9_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_9_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_9_port, QN => 
                           n_1045);
   DLX_INST_DATA_PATH_FETCH_IR_FF_10_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_10_port, B => 
                           DATA_IRAM_signal_10_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_10_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_10_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_10_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_10_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_10_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_10_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_10_port, QN => 
                           n_1046);
   DLX_INST_DATA_PATH_FETCH_IR_FF_11_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_11_port, B => 
                           DATA_IRAM_signal_11_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_11_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_11_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n9, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_11_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_11_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_11_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_11_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_11_port, QN => 
                           n_1047);
   DLX_INST_DATA_PATH_FETCH_IR_FF_12_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_12_port, B => 
                           DATA_IRAM_signal_12_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_12_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_12_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_12_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_12_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_12_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_12_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_12_port, QN => 
                           n_1048);
   DLX_INST_DATA_PATH_FETCH_IR_FF_13_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_13_port, B => 
                           DATA_IRAM_signal_13_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_13_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_13_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_13_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_13_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_13_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_13_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_13_port, QN => 
                           n_1049);
   DLX_INST_DATA_PATH_FETCH_IR_FF_14_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_14_port, B => 
                           DATA_IRAM_signal_14_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_14_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_14_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_14_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_14_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_14_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_14_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_14_port, QN => 
                           n_1050);
   DLX_INST_DATA_PATH_FETCH_IR_FF_15_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, B => 
                           DATA_IRAM_signal_15_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_15_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_15_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_15_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_15_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_15_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_15_n2, Q => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, QN => 
                           n_1051);
   DLX_INST_DATA_PATH_FETCH_IR_FF_16_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_16_port, B => 
                           DATA_IRAM_signal_16_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_16_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_16_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_16_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_16_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_16_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_16_n2, Q => 
                           DLX_INST_IR_OUT_signal_16_port, QN => n_1052);
   DLX_INST_DATA_PATH_FETCH_IR_FF_17_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_17_port, B => 
                           DATA_IRAM_signal_17_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_17_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_17_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_17_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_17_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_17_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_17_n2, Q => 
                           DLX_INST_IR_OUT_signal_17_port, QN => n_1053);
   DLX_INST_DATA_PATH_FETCH_IR_FF_18_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_18_port, B => 
                           DATA_IRAM_signal_18_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_18_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_18_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_18_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_18_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_18_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_18_n2, Q => 
                           DLX_INST_IR_OUT_signal_18_port, QN => n_1054);
   DLX_INST_DATA_PATH_FETCH_IR_FF_19_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_19_port, B => 
                           DATA_IRAM_signal_19_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_19_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_19_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_19_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_19_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_19_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_19_n2, Q => 
                           DLX_INST_IR_OUT_signal_19_port, QN => n_1055);
   DLX_INST_DATA_PATH_FETCH_IR_FF_20_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_20_port, B => 
                           DATA_IRAM_signal_20_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_20_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_20_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_20_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_20_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_20_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_20_n2, Q => 
                           DLX_INST_IR_OUT_signal_20_port, QN => n_1056);
   DLX_INST_DATA_PATH_FETCH_IR_FF_21_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_21_port, B => 
                           DATA_IRAM_signal_21_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_21_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_21_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_21_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_21_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_21_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_21_n2, Q => 
                           DLX_INST_IR_OUT_signal_21_port, QN => n_1057);
   DLX_INST_DATA_PATH_FETCH_IR_FF_22_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_22_port, B => 
                           DATA_IRAM_signal_22_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_22_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_22_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_22_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_22_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_22_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_22_n2, Q => 
                           DLX_INST_IR_OUT_signal_22_port, QN => n_1058);
   DLX_INST_DATA_PATH_FETCH_IR_FF_23_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_23_port, B => 
                           DATA_IRAM_signal_23_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_23_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_23_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n10, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_23_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_23_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_23_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_23_n2, Q => 
                           DLX_INST_IR_OUT_signal_23_port, QN => n_1059);
   DLX_INST_DATA_PATH_FETCH_IR_FF_24_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_24_port, B => 
                           DATA_IRAM_signal_24_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_24_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_24_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n11, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_24_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_24_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_24_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_24_n2, Q => 
                           DLX_INST_IR_OUT_signal_24_port, QN => n_1060);
   DLX_INST_DATA_PATH_FETCH_IR_FF_25_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_25_port, B => 
                           DATA_IRAM_signal_25_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_25_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_25_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n11, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_25_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_25_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_25_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_25_n2, Q => 
                           DLX_INST_IR_OUT_signal_25_port, QN => n_1061);
   DLX_INST_DATA_PATH_FETCH_IR_FF_26_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_26_port, B => 
                           DATA_IRAM_signal_26_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_26_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_26_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n11, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_26_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_26_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_26_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_26_n2, Q => 
                           DLX_INST_IR_OUT_signal_26_port, QN => n_1062);
   DLX_INST_DATA_PATH_FETCH_IR_FF_27_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_27_port, B => 
                           DATA_IRAM_signal_27_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_27_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_27_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n11, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_27_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_27_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_27_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_27_n2, Q => 
                           DLX_INST_IR_OUT_signal_27_port, QN => n_1063);
   DLX_INST_DATA_PATH_FETCH_IR_FF_28_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_28_port, B => 
                           DATA_IRAM_signal_28_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_28_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_28_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n11, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_28_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_28_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_28_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_28_n2, Q => 
                           DLX_INST_IR_OUT_signal_28_port, QN => n_1064);
   DLX_INST_DATA_PATH_FETCH_IR_FF_29_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_29_port, B => 
                           DATA_IRAM_signal_29_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_29_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_29_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n11, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_29_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_29_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_29_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_29_n2, Q => 
                           DLX_INST_IR_OUT_signal_29_port, QN => n_1065);
   DLX_INST_DATA_PATH_FETCH_IR_FF_30_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_30_port, B => 
                           DATA_IRAM_signal_30_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_30_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_30_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n11, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_30_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_30_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_30_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_30_n2, Q => 
                           DLX_INST_IR_OUT_signal_30_port, QN => n_1066);
   DLX_INST_DATA_PATH_FETCH_IR_FF_31_U3 : MUX2_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_31_port, B => 
                           DATA_IRAM_signal_31_port, S => 
                           DLX_INST_IR_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_31_n1);
   DLX_INST_DATA_PATH_FETCH_IR_FF_31_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_IR_n11, A2 => 
                           DLX_INST_IR_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_31_n2);
   DLX_INST_DATA_PATH_FETCH_IR_FF_31_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_31_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_IR_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_IR_FF_31_n2, Q => 
                           DLX_INST_IR_OUT_signal_31_port, QN => n_1067);
   DLX_INST_DATA_PATH_FETCH_NPC_U8 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n16, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n15);
   DLX_INST_DATA_PATH_FETCH_NPC_U7 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n16, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14);
   DLX_INST_DATA_PATH_FETCH_NPC_U6 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n16, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13);
   DLX_INST_DATA_PATH_FETCH_NPC_U5 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n12, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n11);
   DLX_INST_DATA_PATH_FETCH_NPC_U4 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n12, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10);
   DLX_INST_DATA_PATH_FETCH_NPC_U3 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n12, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9);
   DLX_INST_DATA_PATH_FETCH_NPC_U2 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_n4, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n16);
   DLX_INST_DATA_PATH_FETCH_NPC_U1 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_FETCH_n3, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n12);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_0_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_0_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_0_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_0_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_0_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_0_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_0_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_0_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_0_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_0_port, QN => n_1068);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_1_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_1_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_1_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_1_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_1_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_1_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_1_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_1_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_1_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_1_port, QN => n_1069);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_2_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_2_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_2_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_2_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_2_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_2_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_2_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_2_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_2_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_2_port, QN => n_1070);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_3_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_3_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_3_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_3_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_3_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_3_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_3_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_3_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_3_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_3_port, QN => n_1071);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_4_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_4_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_4_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_4_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_4_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_4_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_4_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_4_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_4_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_4_port, QN => n_1072);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_5_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_5_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_5_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_5_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_5_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_5_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_5_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_5_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_5_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_5_port, QN => n_1073);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_6_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_6_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_6_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_6_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_6_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_6_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_6_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_6_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_6_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_6_port, QN => n_1074);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_7_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_7_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_7_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_7_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_7_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_7_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_7_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_7_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_7_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_7_port, QN => n_1075);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_8_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_8_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_8_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_8_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_8_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_8_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_8_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_8_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_8_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_8_port, QN => n_1076);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_9_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_9_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_9_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_9_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_9_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_9_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_9_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_9_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_9_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_9_port, QN => n_1077);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_10_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_10_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_10_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_10_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_10_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_10_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_10_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_10_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n13, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_10_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_10_port, QN => n_1078);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_11_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_11_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_11_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_11_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_11_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n9, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_11_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_11_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_11_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_11_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_11_port, QN => n_1079);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_12_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_12_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_12_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_12_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_12_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_12_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_12_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_12_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_12_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_12_port, QN => n_1080);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_13_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_13_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_13_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_13_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_13_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_13_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_13_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_13_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_13_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_13_port, QN => n_1081);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_14_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_14_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_14_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_14_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_14_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_14_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_14_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_14_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_14_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_14_port, QN => n_1082);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_15_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_15_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_15_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_15_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_15_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_15_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_15_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_15_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_15_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_15_port, QN => n_1083);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_16_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_16_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_16_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_16_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_16_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_16_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_16_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_16_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_16_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_16_port, QN => n_1084);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_17_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_17_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_17_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_17_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_17_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_17_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_17_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_17_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_17_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_17_port, QN => n_1085);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_18_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_18_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_18_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_18_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_18_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_18_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_18_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_18_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_18_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_18_port, QN => n_1086);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_19_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_19_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_19_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_19_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_19_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_19_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_19_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_19_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_19_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_19_port, QN => n_1087);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_20_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_20_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_20_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_20_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_20_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_20_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_20_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_20_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_20_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_20_port, QN => n_1088);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_21_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_21_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_21_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_21_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_21_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_21_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_21_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_21_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n14, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_21_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_21_port, QN => n_1089);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_22_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_22_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_22_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_22_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_22_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_22_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_22_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_22_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_22_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_22_port, QN => n_1090);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_23_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_23_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_23_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_23_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_23_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n10, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_23_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_23_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_23_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_23_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_23_port, QN => n_1091);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_24_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_24_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_24_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_24_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_24_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n11, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_24_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_24_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_24_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_24_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_24_port, QN => n_1092);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_25_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_25_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_25_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_25_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_25_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n11, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_25_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_25_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_25_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_25_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_25_port, QN => n_1093);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_26_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_26_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_26_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_26_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_26_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n11, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_26_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_26_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_26_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_26_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_26_port, QN => n_1094);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_27_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_27_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_27_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_27_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_27_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n11, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_27_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_27_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_27_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_27_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_27_port, QN => n_1095);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_28_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_28_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_28_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_28_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_28_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n11, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_28_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_28_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_28_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_28_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_28_port, QN => n_1096);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_29_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_29_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_29_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_29_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_29_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n11, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_29_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_29_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_29_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_29_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_29_port, QN => n_1097);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_30_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_30_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_30_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_30_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_30_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n11, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_30_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_30_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_30_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_30_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_30_port, QN => n_1098);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_31_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC_OUTs_31_port, B => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_31_port, S => 
                           DLX_INST_NPC_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_31_n1);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_31_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n11, A2 => 
                           DLX_INST_NPC_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_31_n2);
   DLX_INST_DATA_PATH_FETCH_NPC_FF_31_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_31_n1, CK => 
                           DLX_INST_DATA_PATH_FETCH_NPC_n15, RN => 
                           DLX_INST_DATA_PATH_FETCH_NPC_FF_31_n2, Q => 
                           DLX_INST_DATA_PATH_NPC_OUTs_31_port, QN => n_1099);
   DLX_INST_DATA_PATH_DECODE_U10 : OR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_IR_OUT4s_31_port, A2 => 
                           DLX_INST_DATA_PATH_IR_OUT4s_30_port, A3 => 
                           DLX_INST_DATA_PATH_IR_OUT4s_29_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_n13);
   DLX_INST_DATA_PATH_DECODE_U9 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_16_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT4s_11_port, S => 
                           DLX_INST_DATA_PATH_DECODE_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_n1);
   DLX_INST_DATA_PATH_DECODE_U8 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_17_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT4s_12_port, S => 
                           DLX_INST_DATA_PATH_DECODE_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_n2);
   DLX_INST_DATA_PATH_DECODE_U7 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_18_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT4s_13_port, S => 
                           DLX_INST_DATA_PATH_DECODE_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_n3);
   DLX_INST_DATA_PATH_DECODE_U6 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_19_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT4s_14_port, S => 
                           DLX_INST_DATA_PATH_DECODE_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_n4);
   DLX_INST_DATA_PATH_DECODE_U5 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_20_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT4s_15_port, S => 
                           DLX_INST_DATA_PATH_DECODE_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_n5);
   DLX_INST_DATA_PATH_DECODE_U4 : BUF_X1 port map( A => DLX_INST_DATA_PATH_n4, 
                           Z => DLX_INST_DATA_PATH_DECODE_n11);
   DLX_INST_DATA_PATH_DECODE_U3 : BUF_X1 port map( A => DLX_INST_DATA_PATH_n3, 
                           Z => DLX_INST_DATA_PATH_DECODE_n10);
   DLX_INST_DATA_PATH_DECODE_U2 : NOR4_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_IR_OUT4s_28_port, A2 => 
                           DLX_INST_DATA_PATH_IR_OUT4s_27_port, A3 => 
                           DLX_INST_DATA_PATH_IR_OUT4s_26_port, A4 => 
                           DLX_INST_DATA_PATH_DECODE_n13, ZN => 
                           DLX_INST_DATA_PATH_DECODE_n12);
   DLX_INST_DATA_PATH_DECODE_Logic1_port <= '1';
   DLX_INST_DATA_PATH_DECODE_NPC2_U8 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n16, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n15);
   DLX_INST_DATA_PATH_DECODE_NPC2_U7 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n16, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14);
   DLX_INST_DATA_PATH_DECODE_NPC2_U6 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n16, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13);
   DLX_INST_DATA_PATH_DECODE_NPC2_U5 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n11);
   DLX_INST_DATA_PATH_DECODE_NPC2_U4 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10);
   DLX_INST_DATA_PATH_DECODE_NPC2_U3 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9);
   DLX_INST_DATA_PATH_DECODE_NPC2_U2 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n11, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n16);
   DLX_INST_DATA_PATH_DECODE_NPC2_U1 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n10, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n12);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_0_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_0_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_0_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_0_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_0_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_0_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_0_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_0_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_0_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_0_port, QN => n_1100);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_1_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_1_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_1_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_1_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_1_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_1_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_1_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_1_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_1_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_1_port, QN => n_1101);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_2_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_2_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_2_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_2_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_2_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_2_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_2_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_2_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_2_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_2_port, QN => n_1102);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_3_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_3_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_3_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_3_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_3_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_3_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_3_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_3_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_3_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_3_port, QN => n_1103);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_4_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_4_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_4_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_4_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_4_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_4_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_4_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_4_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_4_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_4_port, QN => n_1104);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_5_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_5_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_5_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_5_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_5_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_5_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_5_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_5_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_5_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_5_port, QN => n_1105);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_6_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_6_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_6_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_6_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_6_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_6_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_6_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_6_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_6_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_6_port, QN => n_1106);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_7_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_7_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_7_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_7_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_7_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_7_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_7_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_7_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_7_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_7_port, QN => n_1107);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_8_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_8_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_8_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_8_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_8_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_8_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_8_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_8_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_8_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_8_port, QN => n_1108);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_9_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_9_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_9_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_9_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_9_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_9_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_9_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_9_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_9_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_9_port, QN => n_1109);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_10_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_10_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_10_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_10_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_10_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_10_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_10_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_10_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_10_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_10_port, QN => n_1110);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_11_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_11_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_11_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_11_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_11_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_11_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_11_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_11_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_11_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_11_port, QN => n_1111);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_12_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_12_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_12_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_12_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_12_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_12_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_12_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_12_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_12_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_12_port, QN => n_1112);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_13_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_13_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_13_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_13_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_13_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_13_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_13_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_13_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_13_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_13_port, QN => n_1113);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_14_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_14_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_14_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_14_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_14_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_14_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_14_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_14_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_14_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_14_port, QN => n_1114);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_15_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_15_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_15_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_15_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_15_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_15_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_15_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_15_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_15_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_15_port, QN => n_1115);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_16_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_16_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_16_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_16_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_16_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_16_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_16_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_16_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_16_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_16_port, QN => n_1116);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_17_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_17_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_17_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_17_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_17_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_17_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_17_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_17_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_17_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_17_port, QN => n_1117);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_18_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_18_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_18_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_18_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_18_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_18_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_18_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_18_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_18_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_18_port, QN => n_1118);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_19_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_19_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_19_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_19_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_19_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_19_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_19_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_19_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_19_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_19_port, QN => n_1119);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_20_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_20_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_20_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_20_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_20_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_20_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_20_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_20_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_20_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_20_port, QN => n_1120);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_21_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_21_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_21_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_21_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_21_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_21_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_21_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_21_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_21_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_21_port, QN => n_1121);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_22_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_22_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_22_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_22_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_22_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_22_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_22_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_22_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_22_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_22_port, QN => n_1122);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_23_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_23_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_23_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_23_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_23_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_23_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_23_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_23_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_23_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_23_port, QN => n_1123);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_24_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_24_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_24_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_24_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_24_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_24_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_24_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_24_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_24_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_24_port, QN => n_1124);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_25_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_25_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_25_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_25_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_25_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_25_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_25_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_25_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_25_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_25_port, QN => n_1125);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_26_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_26_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_26_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_26_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_26_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_26_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_26_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_26_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_26_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_26_port, QN => n_1126);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_27_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_27_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_27_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_27_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_27_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_27_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_27_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_27_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_27_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_27_port, QN => n_1127);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_28_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_28_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_28_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_28_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_28_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_28_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_28_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_28_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_28_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_28_port, QN => n_1128);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_29_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_29_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_29_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_29_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_29_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_29_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_29_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_29_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_29_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_29_port, QN => n_1129);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_30_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_30_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_30_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_30_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_30_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_30_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_30_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_30_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_30_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_30_port, QN => n_1130);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_31_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_31_port, B => 
                           DLX_INST_DATA_PATH_NPC_OUTs_31_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_31_n1);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_31_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_31_n2);
   DLX_INST_DATA_PATH_DECODE_NPC2_FF_31_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_31_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_NPC2_FF_31_n2, Q => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_31_port, QN => n_1131);
   DLX_INST_DATA_PATH_DECODE_Imm_U8 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n16, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n15);
   DLX_INST_DATA_PATH_DECODE_Imm_U7 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n16, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14);
   DLX_INST_DATA_PATH_DECODE_Imm_U6 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n16, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13);
   DLX_INST_DATA_PATH_DECODE_Imm_U5 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n11);
   DLX_INST_DATA_PATH_DECODE_Imm_U4 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10);
   DLX_INST_DATA_PATH_DECODE_Imm_U3 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9);
   DLX_INST_DATA_PATH_DECODE_Imm_U2 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n11, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n16);
   DLX_INST_DATA_PATH_DECODE_Imm_U1 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n10, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n12);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_0_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_0_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_0_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_0_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_0_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_0_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_0_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_0_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_0_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_0_port, QN => n_1132);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_1_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_1_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_1_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_1_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_1_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_1_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_1_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_1_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_1_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_1_port, QN => n_1133);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_2_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_2_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_2_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_2_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_2_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_2_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_2_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_2_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_2_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_2_port, QN => n_1134);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_3_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_3_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_3_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_3_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_3_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_3_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_3_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_3_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_3_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_3_port, QN => n_1135);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_4_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_4_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_4_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_4_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_4_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_4_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_4_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_4_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_4_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_4_port, QN => n_1136);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_5_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_5_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_5_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_5_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_5_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_5_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_5_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_5_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_5_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_5_port, QN => n_1137);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_6_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_6_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_6_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_6_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_6_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_6_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_6_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_6_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_6_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_6_port, QN => n_1138);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_7_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_7_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_7_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_7_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_7_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_7_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_7_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_7_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_7_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_7_port, QN => n_1139);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_8_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_8_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_8_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_8_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_8_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_8_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_8_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_8_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_8_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_8_port, QN => n_1140);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_9_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_9_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_9_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_9_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_9_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_9_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_9_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_9_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_9_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_9_port, QN => n_1141);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_10_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_10_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_10_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_10_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_10_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_10_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_10_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_10_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_10_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_10_port, QN => n_1142);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_11_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_11_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_11_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_11_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_11_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n9, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_11_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_11_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_11_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_11_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_11_port, QN => n_1143);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_12_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_12_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_12_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_12_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_12_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_12_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_12_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_12_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_12_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_12_port, QN => n_1144);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_13_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_13_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_13_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_13_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_13_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_13_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_13_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_13_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_13_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_13_port, QN => n_1145);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_14_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_14_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_14_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_14_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_14_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_14_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_14_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_14_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_14_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_14_port, QN => n_1146);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_15_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_15_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_15_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_15_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_15_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_15_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_15_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_15_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_15_port, QN => n_1147);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_16_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_16_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_16_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_16_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_16_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_16_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_16_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_16_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_16_port, QN => n_1148);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_17_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_17_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_17_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_17_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_17_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_17_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_17_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_17_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_17_port, QN => n_1149);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_18_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_18_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_18_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_18_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_18_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_18_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_18_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_18_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_18_port, QN => n_1150);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_19_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_19_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_19_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_19_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_19_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_19_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_19_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_19_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_19_port, QN => n_1151);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_20_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_20_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_20_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_20_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_20_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_20_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_20_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_20_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_20_port, QN => n_1152);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_21_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_21_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_21_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_21_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_21_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_21_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_21_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_21_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_21_port, QN => n_1153);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_22_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_22_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_22_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_22_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_22_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_22_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_22_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_22_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_22_port, QN => n_1154);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_23_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_23_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_23_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_23_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n10, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_23_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_23_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_23_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_23_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_23_port, QN => n_1155);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_24_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_24_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_24_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_24_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n11, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_24_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_24_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_24_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_24_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_24_port, QN => n_1156);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_25_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_25_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_25_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_25_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n11, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_25_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_25_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_25_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_25_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_25_port, QN => n_1157);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_26_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_26_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_26_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_26_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n11, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_26_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_26_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_26_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_26_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_26_port, QN => n_1158);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_27_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_27_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_27_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_27_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n11, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_27_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_27_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_27_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_27_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_27_port, QN => n_1159);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_28_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_28_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_28_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_28_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n11, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_28_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_28_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_28_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_28_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_28_port, QN => n_1160);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_29_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_29_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_29_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_29_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n11, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_29_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_29_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_29_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_29_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_29_port, QN => n_1161);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_30_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_30_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_30_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_30_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n11, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_30_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_30_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_30_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_30_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_30_port, QN => n_1162);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_31_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_Imm_outs_31_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_RegIMM_LATCH_EN_signal, Z => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_31_n1);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_31_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n11, A2 => 
                           DLX_INST_RegIMM_LATCH_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_31_n2);
   DLX_INST_DATA_PATH_DECODE_Imm_FF_31_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_31_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_Imm_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_Imm_FF_31_n2, Q => 
                           DLX_INST_DATA_PATH_Imm_outs_31_port, QN => n_1163);
   DLX_INST_DATA_PATH_DECODE_IR2_U8 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n16, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n15);
   DLX_INST_DATA_PATH_DECODE_IR2_U7 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n16, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14);
   DLX_INST_DATA_PATH_DECODE_IR2_U6 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n16, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13);
   DLX_INST_DATA_PATH_DECODE_IR2_U5 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n11);
   DLX_INST_DATA_PATH_DECODE_IR2_U4 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10);
   DLX_INST_DATA_PATH_DECODE_IR2_U3 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n12, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9);
   DLX_INST_DATA_PATH_DECODE_IR2_U2 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n11, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n16);
   DLX_INST_DATA_PATH_DECODE_IR2_U1 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n10, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n12);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_0_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_0_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_0_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_0_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_0_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_0_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_0_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_0_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_0_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_0_port, QN => n_1164);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_1_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_1_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_1_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_1_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_1_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_1_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_1_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_1_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_1_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_1_port, QN => n_1165);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_2_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_2_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_2_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_2_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_2_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_2_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_2_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_2_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_2_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_2_port, QN => n_1166);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_3_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_3_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_3_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_3_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_3_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_3_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_3_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_3_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_3_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_3_port, QN => n_1167);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_4_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_4_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_4_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_4_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_4_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_4_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_4_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_4_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_4_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_4_port, QN => n_1168);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_5_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_5_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_5_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_5_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_5_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_5_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_5_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_5_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_5_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_5_port, QN => n_1169);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_6_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_6_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_6_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_6_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_6_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_6_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_6_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_6_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_6_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_6_port, QN => n_1170);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_7_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_7_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_7_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_7_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_7_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_7_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_7_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_7_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_7_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_7_port, QN => n_1171);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_8_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_8_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_8_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_8_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_8_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_8_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_8_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_8_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_8_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_8_port, QN => n_1172);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_9_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_9_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_9_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_9_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_9_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_9_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_9_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_9_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_9_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_9_port, QN => n_1173);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_10_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_10_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_10_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_10_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_10_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_10_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_10_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_10_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n13, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_10_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_10_port, QN => n_1174);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_11_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_11_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_11_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_11_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_11_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n9, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_11_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_11_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_11_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_11_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_11_port, QN => n_1175);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_12_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_12_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_12_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_12_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_12_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_12_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_12_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_12_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_12_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_12_port, QN => n_1176);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_13_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_13_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_13_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_13_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_13_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_13_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_13_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_13_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_13_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_13_port, QN => n_1177);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_14_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_14_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_14_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_14_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_14_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_14_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_14_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_14_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_14_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_14_port, QN => n_1178);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_15_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_15_port, B => 
                           DLX_INST_DATA_PATH_DECODE_signExtOut_31_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_15_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_15_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_15_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_15_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_15_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_15_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_15_port, QN => n_1179);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_16_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_16_port, B => 
                           DLX_INST_IR_OUT_signal_16_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_16_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_16_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_16_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_16_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_16_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_16_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_16_port, QN => n_1180);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_17_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_17_port, B => 
                           DLX_INST_IR_OUT_signal_17_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_17_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_17_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_17_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_17_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_17_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_17_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_17_port, QN => n_1181);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_18_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_18_port, B => 
                           DLX_INST_IR_OUT_signal_18_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_18_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_18_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_18_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_18_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_18_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_18_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_18_port, QN => n_1182);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_19_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_19_port, B => 
                           DLX_INST_IR_OUT_signal_19_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_19_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_19_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_19_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_19_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_19_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_19_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_19_port, QN => n_1183);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_20_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_20_port, B => 
                           DLX_INST_IR_OUT_signal_20_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_20_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_20_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_20_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_20_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_20_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_20_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_20_port, QN => n_1184);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_21_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_21_port, B => 
                           DLX_INST_IR_OUT_signal_21_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_21_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_21_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_21_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_21_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_21_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n14, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_21_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_21_port, QN => n_1185);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_22_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_22_port, B => 
                           DLX_INST_IR_OUT_signal_22_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_22_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_22_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_22_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_22_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_22_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_22_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_22_port, QN => n_1186);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_23_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_23_port, B => 
                           DLX_INST_IR_OUT_signal_23_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_23_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_23_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n10, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_23_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_23_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_23_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_23_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_23_port, QN => n_1187);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_24_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_24_port, B => 
                           DLX_INST_IR_OUT_signal_24_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_24_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_24_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_24_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_24_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_24_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_24_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_24_port, QN => n_1188);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_25_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_25_port, B => 
                           DLX_INST_IR_OUT_signal_25_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_25_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_25_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_25_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_25_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_25_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_25_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_25_port, QN => n_1189);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_26_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_26_port, B => 
                           DLX_INST_IR_OUT_signal_26_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_26_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_26_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_26_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_26_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_26_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_26_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_26_port, QN => n_1190);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_27_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_27_port, B => 
                           DLX_INST_IR_OUT_signal_27_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_27_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_27_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_27_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_27_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_27_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_27_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_27_port, QN => n_1191);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_28_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_28_port, B => 
                           DLX_INST_IR_OUT_signal_28_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_28_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_28_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_28_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_28_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_28_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_28_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_28_port, QN => n_1192);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_29_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_29_port, B => 
                           DLX_INST_IR_OUT_signal_29_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_29_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_29_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_29_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_29_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_29_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_29_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_29_port, QN => n_1193);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_30_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_30_port, B => 
                           DLX_INST_IR_OUT_signal_30_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_30_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_30_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_30_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_30_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_30_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_30_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_30_port, QN => n_1194);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_31_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT2s_31_port, B => 
                           DLX_INST_IR_OUT_signal_31_port, S => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_31_n1);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_31_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n11, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_31_n2);
   DLX_INST_DATA_PATH_DECODE_IR2_FF_31_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_31_n1, CK => 
                           DLX_INST_DATA_PATH_DECODE_IR2_n15, RN => 
                           DLX_INST_DATA_PATH_DECODE_IR2_FF_31_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT2s_31_port, QN => n_1195);
   DLX_INST_DATA_PATH_DECODE_RF_U2543 : AND2_X1 port map( A1 => 
                           DLX_INST_RF_WE_signal, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6586);
   DLX_INST_DATA_PATH_DECODE_RF_U2542 : AND3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_n4, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6586, A3 => 
                           DLX_INST_DATA_PATH_DECODE_n5, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6623);
   DLX_INST_DATA_PATH_DECODE_RF_U2541 : AND3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_n2, A2 => 
                           DLX_INST_DATA_PATH_DECODE_n1, A3 => 
                           DLX_INST_DATA_PATH_DECODE_n3, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6583);
   DLX_INST_DATA_PATH_DECODE_RF_U2540 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4676, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1303);
   DLX_INST_DATA_PATH_DECODE_RF_U2539 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4675, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1304);
   DLX_INST_DATA_PATH_DECODE_RF_U2538 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4674, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1305);
   DLX_INST_DATA_PATH_DECODE_RF_U2537 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4673, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1306);
   DLX_INST_DATA_PATH_DECODE_RF_U2536 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4672, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1307);
   DLX_INST_DATA_PATH_DECODE_RF_U2535 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4671, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1308);
   DLX_INST_DATA_PATH_DECODE_RF_U2534 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4670, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1309);
   DLX_INST_DATA_PATH_DECODE_RF_U2533 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4669, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1310);
   DLX_INST_DATA_PATH_DECODE_RF_U2532 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4668, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1311);
   DLX_INST_DATA_PATH_DECODE_RF_U2531 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4667, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1312);
   DLX_INST_DATA_PATH_DECODE_RF_U2530 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4666, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1313);
   DLX_INST_DATA_PATH_DECODE_RF_U2529 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4665, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1314);
   DLX_INST_DATA_PATH_DECODE_RF_U2528 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4664, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1315);
   DLX_INST_DATA_PATH_DECODE_RF_U2527 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4663, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1316);
   DLX_INST_DATA_PATH_DECODE_RF_U2526 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4662, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1317);
   DLX_INST_DATA_PATH_DECODE_RF_U2525 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4661, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1318);
   DLX_INST_DATA_PATH_DECODE_RF_U2524 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4660, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1319);
   DLX_INST_DATA_PATH_DECODE_RF_U2523 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4659, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1320);
   DLX_INST_DATA_PATH_DECODE_RF_U2522 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4658, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1321);
   DLX_INST_DATA_PATH_DECODE_RF_U2521 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4657, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1322);
   DLX_INST_DATA_PATH_DECODE_RF_U2520 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4656, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1323);
   DLX_INST_DATA_PATH_DECODE_RF_U2519 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4655, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1324);
   DLX_INST_DATA_PATH_DECODE_RF_U2518 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4654, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1325);
   DLX_INST_DATA_PATH_DECODE_RF_U2517 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4653, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1326);
   DLX_INST_DATA_PATH_DECODE_RF_U2516 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4652, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1327);
   DLX_INST_DATA_PATH_DECODE_RF_U2515 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4651, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1328);
   DLX_INST_DATA_PATH_DECODE_RF_U2514 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4650, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1329);
   DLX_INST_DATA_PATH_DECODE_RF_U2513 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4649, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1330);
   DLX_INST_DATA_PATH_DECODE_RF_U2512 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4648, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1331);
   DLX_INST_DATA_PATH_DECODE_RF_U2511 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4647, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1332);
   DLX_INST_DATA_PATH_DECODE_RF_U2510 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4646, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1333);
   DLX_INST_DATA_PATH_DECODE_RF_U2509 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4645, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1334);
   DLX_INST_DATA_PATH_DECODE_RF_U2508 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n1, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6626);
   DLX_INST_DATA_PATH_DECODE_RF_U2507 : AND3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_n2, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6626, A3 => 
                           DLX_INST_DATA_PATH_DECODE_n3, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6580);
   DLX_INST_DATA_PATH_DECODE_RF_U2506 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5188, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1335);
   DLX_INST_DATA_PATH_DECODE_RF_U2505 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5187, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1336);
   DLX_INST_DATA_PATH_DECODE_RF_U2504 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5186, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1337);
   DLX_INST_DATA_PATH_DECODE_RF_U2503 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5185, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1338);
   DLX_INST_DATA_PATH_DECODE_RF_U2502 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5184, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1339);
   DLX_INST_DATA_PATH_DECODE_RF_U2501 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5183, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1340);
   DLX_INST_DATA_PATH_DECODE_RF_U2500 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5182, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1341);
   DLX_INST_DATA_PATH_DECODE_RF_U2499 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5181, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1342);
   DLX_INST_DATA_PATH_DECODE_RF_U2498 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5180, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1343);
   DLX_INST_DATA_PATH_DECODE_RF_U2497 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5179, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1344);
   DLX_INST_DATA_PATH_DECODE_RF_U2496 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5178, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1345);
   DLX_INST_DATA_PATH_DECODE_RF_U2495 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5177, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1346);
   DLX_INST_DATA_PATH_DECODE_RF_U2494 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5176, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1347);
   DLX_INST_DATA_PATH_DECODE_RF_U2493 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5175, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1348);
   DLX_INST_DATA_PATH_DECODE_RF_U2492 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5174, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1349);
   DLX_INST_DATA_PATH_DECODE_RF_U2491 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5173, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1350);
   DLX_INST_DATA_PATH_DECODE_RF_U2490 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5172, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1351);
   DLX_INST_DATA_PATH_DECODE_RF_U2489 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5171, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1352);
   DLX_INST_DATA_PATH_DECODE_RF_U2488 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5170, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1353);
   DLX_INST_DATA_PATH_DECODE_RF_U2487 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5169, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1354);
   DLX_INST_DATA_PATH_DECODE_RF_U2486 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5168, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1355);
   DLX_INST_DATA_PATH_DECODE_RF_U2485 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5167, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1356);
   DLX_INST_DATA_PATH_DECODE_RF_U2484 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5166, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1357);
   DLX_INST_DATA_PATH_DECODE_RF_U2483 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5165, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1358);
   DLX_INST_DATA_PATH_DECODE_RF_U2482 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5164, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1359);
   DLX_INST_DATA_PATH_DECODE_RF_U2481 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5163, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1360);
   DLX_INST_DATA_PATH_DECODE_RF_U2480 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5162, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1361);
   DLX_INST_DATA_PATH_DECODE_RF_U2479 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5161, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1362);
   DLX_INST_DATA_PATH_DECODE_RF_U2478 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5160, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1363);
   DLX_INST_DATA_PATH_DECODE_RF_U2477 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5159, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1364);
   DLX_INST_DATA_PATH_DECODE_RF_U2476 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5158, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1365);
   DLX_INST_DATA_PATH_DECODE_RF_U2475 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5157, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1366);
   DLX_INST_DATA_PATH_DECODE_RF_U2474 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n2, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6629);
   DLX_INST_DATA_PATH_DECODE_RF_U2473 : AND3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_n1, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6629, A3 => 
                           DLX_INST_DATA_PATH_DECODE_n3, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6577);
   DLX_INST_DATA_PATH_DECODE_RF_U2472 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4418, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1367);
   DLX_INST_DATA_PATH_DECODE_RF_U2471 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4417, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1368);
   DLX_INST_DATA_PATH_DECODE_RF_U2470 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4416, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1369);
   DLX_INST_DATA_PATH_DECODE_RF_U2469 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4415, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1370);
   DLX_INST_DATA_PATH_DECODE_RF_U2468 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4414, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1371);
   DLX_INST_DATA_PATH_DECODE_RF_U2467 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4413, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1372);
   DLX_INST_DATA_PATH_DECODE_RF_U2466 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4412, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1373);
   DLX_INST_DATA_PATH_DECODE_RF_U2465 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4411, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1374);
   DLX_INST_DATA_PATH_DECODE_RF_U2464 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4410, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1375);
   DLX_INST_DATA_PATH_DECODE_RF_U2463 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4409, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1376);
   DLX_INST_DATA_PATH_DECODE_RF_U2462 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4408, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1377);
   DLX_INST_DATA_PATH_DECODE_RF_U2461 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4407, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1378);
   DLX_INST_DATA_PATH_DECODE_RF_U2460 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4406, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1379);
   DLX_INST_DATA_PATH_DECODE_RF_U2459 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4405, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1380);
   DLX_INST_DATA_PATH_DECODE_RF_U2458 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4404, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1381);
   DLX_INST_DATA_PATH_DECODE_RF_U2457 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4403, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1382);
   DLX_INST_DATA_PATH_DECODE_RF_U2456 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4402, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1383);
   DLX_INST_DATA_PATH_DECODE_RF_U2455 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4401, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1384);
   DLX_INST_DATA_PATH_DECODE_RF_U2454 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4400, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1385);
   DLX_INST_DATA_PATH_DECODE_RF_U2453 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4399, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1386);
   DLX_INST_DATA_PATH_DECODE_RF_U2452 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4398, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1387);
   DLX_INST_DATA_PATH_DECODE_RF_U2451 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4397, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1388);
   DLX_INST_DATA_PATH_DECODE_RF_U2450 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4396, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1389);
   DLX_INST_DATA_PATH_DECODE_RF_U2449 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4395, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1390);
   DLX_INST_DATA_PATH_DECODE_RF_U2448 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4394, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1391);
   DLX_INST_DATA_PATH_DECODE_RF_U2447 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4393, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1392);
   DLX_INST_DATA_PATH_DECODE_RF_U2446 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4392, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1393);
   DLX_INST_DATA_PATH_DECODE_RF_U2445 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4391, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1394);
   DLX_INST_DATA_PATH_DECODE_RF_U2444 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4390, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1395);
   DLX_INST_DATA_PATH_DECODE_RF_U2443 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4389, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1396);
   DLX_INST_DATA_PATH_DECODE_RF_U2442 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1397);
   DLX_INST_DATA_PATH_DECODE_RF_U2441 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4387, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1398);
   DLX_INST_DATA_PATH_DECODE_RF_U2440 : AND3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6626, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6629, A3 => 
                           DLX_INST_DATA_PATH_DECODE_n3, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6574);
   DLX_INST_DATA_PATH_DECODE_RF_U2439 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4644, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1399);
   DLX_INST_DATA_PATH_DECODE_RF_U2438 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4643, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1400);
   DLX_INST_DATA_PATH_DECODE_RF_U2437 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4642, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1401);
   DLX_INST_DATA_PATH_DECODE_RF_U2436 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4641, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1402);
   DLX_INST_DATA_PATH_DECODE_RF_U2435 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4640, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1403);
   DLX_INST_DATA_PATH_DECODE_RF_U2434 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4639, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1404);
   DLX_INST_DATA_PATH_DECODE_RF_U2433 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4638, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1405);
   DLX_INST_DATA_PATH_DECODE_RF_U2432 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4637, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1406);
   DLX_INST_DATA_PATH_DECODE_RF_U2431 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4636, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1407);
   DLX_INST_DATA_PATH_DECODE_RF_U2430 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4635, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1408);
   DLX_INST_DATA_PATH_DECODE_RF_U2429 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4634, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1409);
   DLX_INST_DATA_PATH_DECODE_RF_U2428 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4633, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1410);
   DLX_INST_DATA_PATH_DECODE_RF_U2427 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4632, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1411);
   DLX_INST_DATA_PATH_DECODE_RF_U2426 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4631, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1412);
   DLX_INST_DATA_PATH_DECODE_RF_U2425 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4630, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1413);
   DLX_INST_DATA_PATH_DECODE_RF_U2424 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4629, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1414);
   DLX_INST_DATA_PATH_DECODE_RF_U2423 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4628, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1415);
   DLX_INST_DATA_PATH_DECODE_RF_U2422 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4627, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1416);
   DLX_INST_DATA_PATH_DECODE_RF_U2421 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4626, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1417);
   DLX_INST_DATA_PATH_DECODE_RF_U2420 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4625, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1418);
   DLX_INST_DATA_PATH_DECODE_RF_U2419 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4624, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1419);
   DLX_INST_DATA_PATH_DECODE_RF_U2418 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4623, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1420);
   DLX_INST_DATA_PATH_DECODE_RF_U2417 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4622, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1421);
   DLX_INST_DATA_PATH_DECODE_RF_U2416 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4621, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1422);
   DLX_INST_DATA_PATH_DECODE_RF_U2415 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4620, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1423);
   DLX_INST_DATA_PATH_DECODE_RF_U2414 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4619, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1424);
   DLX_INST_DATA_PATH_DECODE_RF_U2413 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4618, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1425);
   DLX_INST_DATA_PATH_DECODE_RF_U2412 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4617, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1426);
   DLX_INST_DATA_PATH_DECODE_RF_U2411 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4616, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1427);
   DLX_INST_DATA_PATH_DECODE_RF_U2410 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4615, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1428);
   DLX_INST_DATA_PATH_DECODE_RF_U2409 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4614, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1429);
   DLX_INST_DATA_PATH_DECODE_RF_U2408 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4613, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1430);
   DLX_INST_DATA_PATH_DECODE_RF_U2407 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6626, A2 => 
                           DLX_INST_DATA_PATH_DECODE_n3, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6629, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6571);
   DLX_INST_DATA_PATH_DECODE_RF_U2406 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4386, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1431);
   DLX_INST_DATA_PATH_DECODE_RF_U2405 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4385, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1432);
   DLX_INST_DATA_PATH_DECODE_RF_U2404 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4384, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1433);
   DLX_INST_DATA_PATH_DECODE_RF_U2403 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4383, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1434);
   DLX_INST_DATA_PATH_DECODE_RF_U2402 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1435);
   DLX_INST_DATA_PATH_DECODE_RF_U2401 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4381, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1436);
   DLX_INST_DATA_PATH_DECODE_RF_U2400 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4380, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1437);
   DLX_INST_DATA_PATH_DECODE_RF_U2399 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4379, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1438);
   DLX_INST_DATA_PATH_DECODE_RF_U2398 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4378, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1439);
   DLX_INST_DATA_PATH_DECODE_RF_U2397 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1440);
   DLX_INST_DATA_PATH_DECODE_RF_U2396 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4376, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1441);
   DLX_INST_DATA_PATH_DECODE_RF_U2395 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4375, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1442);
   DLX_INST_DATA_PATH_DECODE_RF_U2394 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4374, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1443);
   DLX_INST_DATA_PATH_DECODE_RF_U2393 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4373, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1444);
   DLX_INST_DATA_PATH_DECODE_RF_U2392 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4372, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1445);
   DLX_INST_DATA_PATH_DECODE_RF_U2391 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1446);
   DLX_INST_DATA_PATH_DECODE_RF_U2390 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4370, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1447);
   DLX_INST_DATA_PATH_DECODE_RF_U2389 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4369, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1448);
   DLX_INST_DATA_PATH_DECODE_RF_U2388 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4368, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1449);
   DLX_INST_DATA_PATH_DECODE_RF_U2387 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4367, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1450);
   DLX_INST_DATA_PATH_DECODE_RF_U2386 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4366, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1451);
   DLX_INST_DATA_PATH_DECODE_RF_U2385 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4365, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1452);
   DLX_INST_DATA_PATH_DECODE_RF_U2384 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4364, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1453);
   DLX_INST_DATA_PATH_DECODE_RF_U2383 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4363, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1454);
   DLX_INST_DATA_PATH_DECODE_RF_U2382 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1455);
   DLX_INST_DATA_PATH_DECODE_RF_U2381 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4361, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1456);
   DLX_INST_DATA_PATH_DECODE_RF_U2380 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4360, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1457);
   DLX_INST_DATA_PATH_DECODE_RF_U2379 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4359, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1458);
   DLX_INST_DATA_PATH_DECODE_RF_U2378 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1459);
   DLX_INST_DATA_PATH_DECODE_RF_U2377 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1460);
   DLX_INST_DATA_PATH_DECODE_RF_U2376 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4356, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1461);
   DLX_INST_DATA_PATH_DECODE_RF_U2375 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4355, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1462);
   DLX_INST_DATA_PATH_DECODE_RF_U2374 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_n1, A2 => 
                           DLX_INST_DATA_PATH_DECODE_n3, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6629, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6568);
   DLX_INST_DATA_PATH_DECODE_RF_U2373 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4964, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1463);
   DLX_INST_DATA_PATH_DECODE_RF_U2372 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4963, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1464);
   DLX_INST_DATA_PATH_DECODE_RF_U2371 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4962, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1465);
   DLX_INST_DATA_PATH_DECODE_RF_U2370 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1466);
   DLX_INST_DATA_PATH_DECODE_RF_U2369 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4960, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1467);
   DLX_INST_DATA_PATH_DECODE_RF_U2368 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4959, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1468);
   DLX_INST_DATA_PATH_DECODE_RF_U2367 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4958, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1469);
   DLX_INST_DATA_PATH_DECODE_RF_U2366 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4957, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1470);
   DLX_INST_DATA_PATH_DECODE_RF_U2365 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4956, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1471);
   DLX_INST_DATA_PATH_DECODE_RF_U2364 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4955, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1472);
   DLX_INST_DATA_PATH_DECODE_RF_U2363 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4954, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1473);
   DLX_INST_DATA_PATH_DECODE_RF_U2362 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4953, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1474);
   DLX_INST_DATA_PATH_DECODE_RF_U2361 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1475);
   DLX_INST_DATA_PATH_DECODE_RF_U2360 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4951, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1476);
   DLX_INST_DATA_PATH_DECODE_RF_U2359 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4950, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1477);
   DLX_INST_DATA_PATH_DECODE_RF_U2358 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4949, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1478);
   DLX_INST_DATA_PATH_DECODE_RF_U2357 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4948, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1479);
   DLX_INST_DATA_PATH_DECODE_RF_U2356 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1480);
   DLX_INST_DATA_PATH_DECODE_RF_U2355 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4946, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1481);
   DLX_INST_DATA_PATH_DECODE_RF_U2354 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4945, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1482);
   DLX_INST_DATA_PATH_DECODE_RF_U2353 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4944, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1483);
   DLX_INST_DATA_PATH_DECODE_RF_U2352 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4943, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1484);
   DLX_INST_DATA_PATH_DECODE_RF_U2351 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1485);
   DLX_INST_DATA_PATH_DECODE_RF_U2350 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4941, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1486);
   DLX_INST_DATA_PATH_DECODE_RF_U2349 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4940, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1487);
   DLX_INST_DATA_PATH_DECODE_RF_U2348 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4939, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1488);
   DLX_INST_DATA_PATH_DECODE_RF_U2347 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4938, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1489);
   DLX_INST_DATA_PATH_DECODE_RF_U2346 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1490);
   DLX_INST_DATA_PATH_DECODE_RF_U2345 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4936, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1491);
   DLX_INST_DATA_PATH_DECODE_RF_U2344 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4935, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1492);
   DLX_INST_DATA_PATH_DECODE_RF_U2343 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4934, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1493);
   DLX_INST_DATA_PATH_DECODE_RF_U2342 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4933, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1494);
   DLX_INST_DATA_PATH_DECODE_RF_U2341 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_n2, A2 => 
                           DLX_INST_DATA_PATH_DECODE_n3, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6626, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6565);
   DLX_INST_DATA_PATH_DECODE_RF_U2340 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4354, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1495);
   DLX_INST_DATA_PATH_DECODE_RF_U2339 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4353, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1496);
   DLX_INST_DATA_PATH_DECODE_RF_U2338 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1497);
   DLX_INST_DATA_PATH_DECODE_RF_U2337 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4351, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1498);
   DLX_INST_DATA_PATH_DECODE_RF_U2336 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4350, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1499);
   DLX_INST_DATA_PATH_DECODE_RF_U2335 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4349, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1500);
   DLX_INST_DATA_PATH_DECODE_RF_U2334 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4348, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1501);
   DLX_INST_DATA_PATH_DECODE_RF_U2333 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1502);
   DLX_INST_DATA_PATH_DECODE_RF_U2332 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4346, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1503);
   DLX_INST_DATA_PATH_DECODE_RF_U2331 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4345, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1504);
   DLX_INST_DATA_PATH_DECODE_RF_U2330 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4344, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1505);
   DLX_INST_DATA_PATH_DECODE_RF_U2329 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4343, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1506);
   DLX_INST_DATA_PATH_DECODE_RF_U2328 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4342, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1507);
   DLX_INST_DATA_PATH_DECODE_RF_U2327 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4341, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1508);
   DLX_INST_DATA_PATH_DECODE_RF_U2326 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4340, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1509);
   DLX_INST_DATA_PATH_DECODE_RF_U2325 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4339, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1510);
   DLX_INST_DATA_PATH_DECODE_RF_U2324 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4338, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1511);
   DLX_INST_DATA_PATH_DECODE_RF_U2323 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4337, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1512);
   DLX_INST_DATA_PATH_DECODE_RF_U2322 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4336, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1513);
   DLX_INST_DATA_PATH_DECODE_RF_U2321 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4335, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1514);
   DLX_INST_DATA_PATH_DECODE_RF_U2320 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4334, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1515);
   DLX_INST_DATA_PATH_DECODE_RF_U2319 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4333, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1516);
   DLX_INST_DATA_PATH_DECODE_RF_U2318 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4332, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1517);
   DLX_INST_DATA_PATH_DECODE_RF_U2317 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4331, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1518);
   DLX_INST_DATA_PATH_DECODE_RF_U2316 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4330, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1519);
   DLX_INST_DATA_PATH_DECODE_RF_U2315 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4329, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1520);
   DLX_INST_DATA_PATH_DECODE_RF_U2314 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4328, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1521);
   DLX_INST_DATA_PATH_DECODE_RF_U2313 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4327, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1522);
   DLX_INST_DATA_PATH_DECODE_RF_U2312 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4326, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1523);
   DLX_INST_DATA_PATH_DECODE_RF_U2311 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4325, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1524);
   DLX_INST_DATA_PATH_DECODE_RF_U2310 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4324, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1525);
   DLX_INST_DATA_PATH_DECODE_RF_U2309 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4323, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1526);
   DLX_INST_DATA_PATH_DECODE_RF_U2308 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_n2, A2 => 
                           DLX_INST_DATA_PATH_DECODE_n3, A3 => 
                           DLX_INST_DATA_PATH_DECODE_n1, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6561);
   DLX_INST_DATA_PATH_DECODE_RF_U2307 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4612, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1527);
   DLX_INST_DATA_PATH_DECODE_RF_U2306 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4611, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1528);
   DLX_INST_DATA_PATH_DECODE_RF_U2305 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4610, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1529);
   DLX_INST_DATA_PATH_DECODE_RF_U2304 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4609, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1530);
   DLX_INST_DATA_PATH_DECODE_RF_U2303 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4608, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1531);
   DLX_INST_DATA_PATH_DECODE_RF_U2302 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4607, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1532);
   DLX_INST_DATA_PATH_DECODE_RF_U2301 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4606, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1533);
   DLX_INST_DATA_PATH_DECODE_RF_U2300 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4605, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1534);
   DLX_INST_DATA_PATH_DECODE_RF_U2299 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4604, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1535);
   DLX_INST_DATA_PATH_DECODE_RF_U2298 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4603, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1536);
   DLX_INST_DATA_PATH_DECODE_RF_U2297 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4602, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1537);
   DLX_INST_DATA_PATH_DECODE_RF_U2296 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4601, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1538);
   DLX_INST_DATA_PATH_DECODE_RF_U2295 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4600, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1539);
   DLX_INST_DATA_PATH_DECODE_RF_U2294 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4599, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1540);
   DLX_INST_DATA_PATH_DECODE_RF_U2293 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4598, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1541);
   DLX_INST_DATA_PATH_DECODE_RF_U2292 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4597, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1542);
   DLX_INST_DATA_PATH_DECODE_RF_U2291 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4596, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1543);
   DLX_INST_DATA_PATH_DECODE_RF_U2290 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4595, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1544);
   DLX_INST_DATA_PATH_DECODE_RF_U2289 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4594, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1545);
   DLX_INST_DATA_PATH_DECODE_RF_U2288 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4593, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1546);
   DLX_INST_DATA_PATH_DECODE_RF_U2287 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4592, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1547);
   DLX_INST_DATA_PATH_DECODE_RF_U2286 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4591, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1548);
   DLX_INST_DATA_PATH_DECODE_RF_U2285 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4590, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1549);
   DLX_INST_DATA_PATH_DECODE_RF_U2284 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4589, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1550);
   DLX_INST_DATA_PATH_DECODE_RF_U2283 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4588, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1551);
   DLX_INST_DATA_PATH_DECODE_RF_U2282 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4587, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1552);
   DLX_INST_DATA_PATH_DECODE_RF_U2281 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4586, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1553);
   DLX_INST_DATA_PATH_DECODE_RF_U2280 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4585, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1554);
   DLX_INST_DATA_PATH_DECODE_RF_U2279 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4584, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1555);
   DLX_INST_DATA_PATH_DECODE_RF_U2278 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4583, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1556);
   DLX_INST_DATA_PATH_DECODE_RF_U2277 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4582, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1557);
   DLX_INST_DATA_PATH_DECODE_RF_U2276 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4581, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1558);
   DLX_INST_DATA_PATH_DECODE_RF_U2275 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n4, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6584);
   DLX_INST_DATA_PATH_DECODE_RF_U2274 : AND3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6586, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6584, A3 => 
                           DLX_INST_DATA_PATH_DECODE_n5, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6606);
   DLX_INST_DATA_PATH_DECODE_RF_U2273 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4580, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1559);
   DLX_INST_DATA_PATH_DECODE_RF_U2272 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4579, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1560);
   DLX_INST_DATA_PATH_DECODE_RF_U2271 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4578, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1561);
   DLX_INST_DATA_PATH_DECODE_RF_U2270 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4577, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1562);
   DLX_INST_DATA_PATH_DECODE_RF_U2269 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4576, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1563);
   DLX_INST_DATA_PATH_DECODE_RF_U2268 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4575, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1564);
   DLX_INST_DATA_PATH_DECODE_RF_U2267 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4574, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1565);
   DLX_INST_DATA_PATH_DECODE_RF_U2266 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4573, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1566);
   DLX_INST_DATA_PATH_DECODE_RF_U2265 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4572, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1567);
   DLX_INST_DATA_PATH_DECODE_RF_U2264 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4571, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1568);
   DLX_INST_DATA_PATH_DECODE_RF_U2263 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4570, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1569);
   DLX_INST_DATA_PATH_DECODE_RF_U2262 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4569, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1570);
   DLX_INST_DATA_PATH_DECODE_RF_U2261 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4568, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1571);
   DLX_INST_DATA_PATH_DECODE_RF_U2260 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4567, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1572);
   DLX_INST_DATA_PATH_DECODE_RF_U2259 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4566, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1573);
   DLX_INST_DATA_PATH_DECODE_RF_U2258 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4565, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1574);
   DLX_INST_DATA_PATH_DECODE_RF_U2257 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4564, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1575);
   DLX_INST_DATA_PATH_DECODE_RF_U2256 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4563, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1576);
   DLX_INST_DATA_PATH_DECODE_RF_U2255 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4562, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1577);
   DLX_INST_DATA_PATH_DECODE_RF_U2254 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4561, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1578);
   DLX_INST_DATA_PATH_DECODE_RF_U2253 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4560, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1579);
   DLX_INST_DATA_PATH_DECODE_RF_U2252 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4559, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1580);
   DLX_INST_DATA_PATH_DECODE_RF_U2251 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4558, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1581);
   DLX_INST_DATA_PATH_DECODE_RF_U2250 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4557, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1582);
   DLX_INST_DATA_PATH_DECODE_RF_U2249 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4556, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1583);
   DLX_INST_DATA_PATH_DECODE_RF_U2248 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4555, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1584);
   DLX_INST_DATA_PATH_DECODE_RF_U2247 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4554, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1585);
   DLX_INST_DATA_PATH_DECODE_RF_U2246 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4553, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1586);
   DLX_INST_DATA_PATH_DECODE_RF_U2245 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4552, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1587);
   DLX_INST_DATA_PATH_DECODE_RF_U2244 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4551, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1588);
   DLX_INST_DATA_PATH_DECODE_RF_U2243 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4550, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1589);
   DLX_INST_DATA_PATH_DECODE_RF_U2242 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4549, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1590);
   DLX_INST_DATA_PATH_DECODE_RF_U2241 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4932, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1591);
   DLX_INST_DATA_PATH_DECODE_RF_U2240 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4931, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1592);
   DLX_INST_DATA_PATH_DECODE_RF_U2239 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4930, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1593);
   DLX_INST_DATA_PATH_DECODE_RF_U2238 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4929, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1594);
   DLX_INST_DATA_PATH_DECODE_RF_U2237 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4928, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1595);
   DLX_INST_DATA_PATH_DECODE_RF_U2236 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4927, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1596);
   DLX_INST_DATA_PATH_DECODE_RF_U2235 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4926, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1597);
   DLX_INST_DATA_PATH_DECODE_RF_U2234 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4925, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1598);
   DLX_INST_DATA_PATH_DECODE_RF_U2233 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4924, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1599);
   DLX_INST_DATA_PATH_DECODE_RF_U2232 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4923, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1600);
   DLX_INST_DATA_PATH_DECODE_RF_U2231 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4922, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1601);
   DLX_INST_DATA_PATH_DECODE_RF_U2230 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4921, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1602);
   DLX_INST_DATA_PATH_DECODE_RF_U2229 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4920, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1603);
   DLX_INST_DATA_PATH_DECODE_RF_U2228 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4919, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1604);
   DLX_INST_DATA_PATH_DECODE_RF_U2227 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4918, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1605);
   DLX_INST_DATA_PATH_DECODE_RF_U2226 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4917, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1606);
   DLX_INST_DATA_PATH_DECODE_RF_U2225 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4916, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1607);
   DLX_INST_DATA_PATH_DECODE_RF_U2224 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4915, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1608);
   DLX_INST_DATA_PATH_DECODE_RF_U2223 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4914, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1609);
   DLX_INST_DATA_PATH_DECODE_RF_U2222 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4913, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1610);
   DLX_INST_DATA_PATH_DECODE_RF_U2221 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4912, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1611);
   DLX_INST_DATA_PATH_DECODE_RF_U2220 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4911, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1612);
   DLX_INST_DATA_PATH_DECODE_RF_U2219 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4910, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1613);
   DLX_INST_DATA_PATH_DECODE_RF_U2218 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4909, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1614);
   DLX_INST_DATA_PATH_DECODE_RF_U2217 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4908, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1615);
   DLX_INST_DATA_PATH_DECODE_RF_U2216 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4907, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1616);
   DLX_INST_DATA_PATH_DECODE_RF_U2215 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4906, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1617);
   DLX_INST_DATA_PATH_DECODE_RF_U2214 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4905, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1618);
   DLX_INST_DATA_PATH_DECODE_RF_U2213 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4904, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1619);
   DLX_INST_DATA_PATH_DECODE_RF_U2212 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4903, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1620);
   DLX_INST_DATA_PATH_DECODE_RF_U2211 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4902, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1621);
   DLX_INST_DATA_PATH_DECODE_RF_U2210 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4901, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1622);
   DLX_INST_DATA_PATH_DECODE_RF_U2209 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4322, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1623);
   DLX_INST_DATA_PATH_DECODE_RF_U2208 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4321, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1624);
   DLX_INST_DATA_PATH_DECODE_RF_U2207 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4320, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1625);
   DLX_INST_DATA_PATH_DECODE_RF_U2206 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4319, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1626);
   DLX_INST_DATA_PATH_DECODE_RF_U2205 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4318, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1627);
   DLX_INST_DATA_PATH_DECODE_RF_U2204 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4317, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1628);
   DLX_INST_DATA_PATH_DECODE_RF_U2203 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4316, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1629);
   DLX_INST_DATA_PATH_DECODE_RF_U2202 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4315, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1630);
   DLX_INST_DATA_PATH_DECODE_RF_U2201 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4314, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1631);
   DLX_INST_DATA_PATH_DECODE_RF_U2200 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4313, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1632);
   DLX_INST_DATA_PATH_DECODE_RF_U2199 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4312, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1633);
   DLX_INST_DATA_PATH_DECODE_RF_U2198 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4311, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1634);
   DLX_INST_DATA_PATH_DECODE_RF_U2197 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4310, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1635);
   DLX_INST_DATA_PATH_DECODE_RF_U2196 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4309, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1636);
   DLX_INST_DATA_PATH_DECODE_RF_U2195 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4308, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1637);
   DLX_INST_DATA_PATH_DECODE_RF_U2194 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4307, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1638);
   DLX_INST_DATA_PATH_DECODE_RF_U2193 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4306, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1639);
   DLX_INST_DATA_PATH_DECODE_RF_U2192 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4305, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1640);
   DLX_INST_DATA_PATH_DECODE_RF_U2191 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4304, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1641);
   DLX_INST_DATA_PATH_DECODE_RF_U2190 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4303, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1642);
   DLX_INST_DATA_PATH_DECODE_RF_U2189 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4302, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1643);
   DLX_INST_DATA_PATH_DECODE_RF_U2188 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4301, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1644);
   DLX_INST_DATA_PATH_DECODE_RF_U2187 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4300, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1645);
   DLX_INST_DATA_PATH_DECODE_RF_U2186 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4299, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1646);
   DLX_INST_DATA_PATH_DECODE_RF_U2185 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4298, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1647);
   DLX_INST_DATA_PATH_DECODE_RF_U2184 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4297, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1648);
   DLX_INST_DATA_PATH_DECODE_RF_U2183 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4296, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1649);
   DLX_INST_DATA_PATH_DECODE_RF_U2182 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4295, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1650);
   DLX_INST_DATA_PATH_DECODE_RF_U2181 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4294, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1651);
   DLX_INST_DATA_PATH_DECODE_RF_U2180 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4293, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1652);
   DLX_INST_DATA_PATH_DECODE_RF_U2179 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4292, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1653);
   DLX_INST_DATA_PATH_DECODE_RF_U2178 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4291, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1654);
   DLX_INST_DATA_PATH_DECODE_RF_U2177 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4290, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1655);
   DLX_INST_DATA_PATH_DECODE_RF_U2176 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4289, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1656);
   DLX_INST_DATA_PATH_DECODE_RF_U2175 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4288, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1657);
   DLX_INST_DATA_PATH_DECODE_RF_U2174 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4287, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1658);
   DLX_INST_DATA_PATH_DECODE_RF_U2173 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4286, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1659);
   DLX_INST_DATA_PATH_DECODE_RF_U2172 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4285, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1660);
   DLX_INST_DATA_PATH_DECODE_RF_U2171 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4284, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1661);
   DLX_INST_DATA_PATH_DECODE_RF_U2170 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4283, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1662);
   DLX_INST_DATA_PATH_DECODE_RF_U2169 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4282, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1663);
   DLX_INST_DATA_PATH_DECODE_RF_U2168 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4281, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1664);
   DLX_INST_DATA_PATH_DECODE_RF_U2167 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4280, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1665);
   DLX_INST_DATA_PATH_DECODE_RF_U2166 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4279, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1666);
   DLX_INST_DATA_PATH_DECODE_RF_U2165 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4278, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1667);
   DLX_INST_DATA_PATH_DECODE_RF_U2164 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4277, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1668);
   DLX_INST_DATA_PATH_DECODE_RF_U2163 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4276, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1669);
   DLX_INST_DATA_PATH_DECODE_RF_U2162 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4275, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1670);
   DLX_INST_DATA_PATH_DECODE_RF_U2161 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4274, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1671);
   DLX_INST_DATA_PATH_DECODE_RF_U2160 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4273, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1672);
   DLX_INST_DATA_PATH_DECODE_RF_U2159 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4272, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1673);
   DLX_INST_DATA_PATH_DECODE_RF_U2158 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4271, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1674);
   DLX_INST_DATA_PATH_DECODE_RF_U2157 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4270, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1675);
   DLX_INST_DATA_PATH_DECODE_RF_U2156 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4269, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1676);
   DLX_INST_DATA_PATH_DECODE_RF_U2155 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4268, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1677);
   DLX_INST_DATA_PATH_DECODE_RF_U2154 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4267, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1678);
   DLX_INST_DATA_PATH_DECODE_RF_U2153 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4266, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1679);
   DLX_INST_DATA_PATH_DECODE_RF_U2152 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4265, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1680);
   DLX_INST_DATA_PATH_DECODE_RF_U2151 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4264, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1681);
   DLX_INST_DATA_PATH_DECODE_RF_U2150 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4263, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1682);
   DLX_INST_DATA_PATH_DECODE_RF_U2149 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4262, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1683);
   DLX_INST_DATA_PATH_DECODE_RF_U2148 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4261, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1684);
   DLX_INST_DATA_PATH_DECODE_RF_U2147 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4260, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1685);
   DLX_INST_DATA_PATH_DECODE_RF_U2146 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4259, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1686);
   DLX_INST_DATA_PATH_DECODE_RF_U2145 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4900, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1687);
   DLX_INST_DATA_PATH_DECODE_RF_U2144 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4899, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1688);
   DLX_INST_DATA_PATH_DECODE_RF_U2143 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4898, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1689);
   DLX_INST_DATA_PATH_DECODE_RF_U2142 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4897, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1690);
   DLX_INST_DATA_PATH_DECODE_RF_U2141 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4896, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1691);
   DLX_INST_DATA_PATH_DECODE_RF_U2140 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4895, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1692);
   DLX_INST_DATA_PATH_DECODE_RF_U2139 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4894, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1693);
   DLX_INST_DATA_PATH_DECODE_RF_U2138 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4893, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1694);
   DLX_INST_DATA_PATH_DECODE_RF_U2137 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4892, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1695);
   DLX_INST_DATA_PATH_DECODE_RF_U2136 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4891, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1696);
   DLX_INST_DATA_PATH_DECODE_RF_U2135 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4890, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1697);
   DLX_INST_DATA_PATH_DECODE_RF_U2134 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4889, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1698);
   DLX_INST_DATA_PATH_DECODE_RF_U2133 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4888, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1699);
   DLX_INST_DATA_PATH_DECODE_RF_U2132 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4887, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1700);
   DLX_INST_DATA_PATH_DECODE_RF_U2131 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4886, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1701);
   DLX_INST_DATA_PATH_DECODE_RF_U2130 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4885, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1702);
   DLX_INST_DATA_PATH_DECODE_RF_U2129 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4884, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1703);
   DLX_INST_DATA_PATH_DECODE_RF_U2128 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4883, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1704);
   DLX_INST_DATA_PATH_DECODE_RF_U2127 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4882, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1705);
   DLX_INST_DATA_PATH_DECODE_RF_U2126 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4881, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1706);
   DLX_INST_DATA_PATH_DECODE_RF_U2125 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4880, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1707);
   DLX_INST_DATA_PATH_DECODE_RF_U2124 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4879, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1708);
   DLX_INST_DATA_PATH_DECODE_RF_U2123 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4878, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1709);
   DLX_INST_DATA_PATH_DECODE_RF_U2122 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4877, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1710);
   DLX_INST_DATA_PATH_DECODE_RF_U2121 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4876, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1711);
   DLX_INST_DATA_PATH_DECODE_RF_U2120 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4875, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1712);
   DLX_INST_DATA_PATH_DECODE_RF_U2119 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4874, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1713);
   DLX_INST_DATA_PATH_DECODE_RF_U2118 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4873, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1714);
   DLX_INST_DATA_PATH_DECODE_RF_U2117 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4872, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1715);
   DLX_INST_DATA_PATH_DECODE_RF_U2116 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4871, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1716);
   DLX_INST_DATA_PATH_DECODE_RF_U2115 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4870, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1717);
   DLX_INST_DATA_PATH_DECODE_RF_U2114 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4869, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1718);
   DLX_INST_DATA_PATH_DECODE_RF_U2113 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5156, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1719);
   DLX_INST_DATA_PATH_DECODE_RF_U2112 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5155, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1720);
   DLX_INST_DATA_PATH_DECODE_RF_U2111 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5154, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1721);
   DLX_INST_DATA_PATH_DECODE_RF_U2110 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5153, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1722);
   DLX_INST_DATA_PATH_DECODE_RF_U2109 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5152, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1723);
   DLX_INST_DATA_PATH_DECODE_RF_U2108 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5151, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1724);
   DLX_INST_DATA_PATH_DECODE_RF_U2107 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5150, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1725);
   DLX_INST_DATA_PATH_DECODE_RF_U2106 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5149, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1726);
   DLX_INST_DATA_PATH_DECODE_RF_U2105 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5148, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1727);
   DLX_INST_DATA_PATH_DECODE_RF_U2104 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5147, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1728);
   DLX_INST_DATA_PATH_DECODE_RF_U2103 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5146, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1729);
   DLX_INST_DATA_PATH_DECODE_RF_U2102 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5145, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1730);
   DLX_INST_DATA_PATH_DECODE_RF_U2101 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5144, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1731);
   DLX_INST_DATA_PATH_DECODE_RF_U2100 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5143, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1732);
   DLX_INST_DATA_PATH_DECODE_RF_U2099 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5142, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1733);
   DLX_INST_DATA_PATH_DECODE_RF_U2098 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5141, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1734);
   DLX_INST_DATA_PATH_DECODE_RF_U2097 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5140, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1735);
   DLX_INST_DATA_PATH_DECODE_RF_U2096 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5139, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1736);
   DLX_INST_DATA_PATH_DECODE_RF_U2095 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5138, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1737);
   DLX_INST_DATA_PATH_DECODE_RF_U2094 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5137, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1738);
   DLX_INST_DATA_PATH_DECODE_RF_U2093 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5136, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1739);
   DLX_INST_DATA_PATH_DECODE_RF_U2092 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5135, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1740);
   DLX_INST_DATA_PATH_DECODE_RF_U2091 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5134, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1741);
   DLX_INST_DATA_PATH_DECODE_RF_U2090 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5133, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1742);
   DLX_INST_DATA_PATH_DECODE_RF_U2089 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5132, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1743);
   DLX_INST_DATA_PATH_DECODE_RF_U2088 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5131, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1744);
   DLX_INST_DATA_PATH_DECODE_RF_U2087 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5130, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1745);
   DLX_INST_DATA_PATH_DECODE_RF_U2086 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5129, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1746);
   DLX_INST_DATA_PATH_DECODE_RF_U2085 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5128, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1747);
   DLX_INST_DATA_PATH_DECODE_RF_U2084 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5127, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1748);
   DLX_INST_DATA_PATH_DECODE_RF_U2083 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5126, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1749);
   DLX_INST_DATA_PATH_DECODE_RF_U2082 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5125, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1750);
   DLX_INST_DATA_PATH_DECODE_RF_U2081 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4548, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1751);
   DLX_INST_DATA_PATH_DECODE_RF_U2080 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4547, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1752);
   DLX_INST_DATA_PATH_DECODE_RF_U2079 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4546, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1753);
   DLX_INST_DATA_PATH_DECODE_RF_U2078 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4545, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1754);
   DLX_INST_DATA_PATH_DECODE_RF_U2077 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4544, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1755);
   DLX_INST_DATA_PATH_DECODE_RF_U2076 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4543, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1756);
   DLX_INST_DATA_PATH_DECODE_RF_U2075 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4542, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1757);
   DLX_INST_DATA_PATH_DECODE_RF_U2074 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4541, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1758);
   DLX_INST_DATA_PATH_DECODE_RF_U2073 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4540, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1759);
   DLX_INST_DATA_PATH_DECODE_RF_U2072 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4539, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1760);
   DLX_INST_DATA_PATH_DECODE_RF_U2071 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4538, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1761);
   DLX_INST_DATA_PATH_DECODE_RF_U2070 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4537, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1762);
   DLX_INST_DATA_PATH_DECODE_RF_U2069 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4536, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1763);
   DLX_INST_DATA_PATH_DECODE_RF_U2068 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4535, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1764);
   DLX_INST_DATA_PATH_DECODE_RF_U2067 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4534, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1765);
   DLX_INST_DATA_PATH_DECODE_RF_U2066 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4533, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1766);
   DLX_INST_DATA_PATH_DECODE_RF_U2065 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4532, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1767);
   DLX_INST_DATA_PATH_DECODE_RF_U2064 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4531, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1768);
   DLX_INST_DATA_PATH_DECODE_RF_U2063 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4530, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1769);
   DLX_INST_DATA_PATH_DECODE_RF_U2062 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4529, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1770);
   DLX_INST_DATA_PATH_DECODE_RF_U2061 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4528, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1771);
   DLX_INST_DATA_PATH_DECODE_RF_U2060 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4527, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1772);
   DLX_INST_DATA_PATH_DECODE_RF_U2059 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4526, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1773);
   DLX_INST_DATA_PATH_DECODE_RF_U2058 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4525, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1774);
   DLX_INST_DATA_PATH_DECODE_RF_U2057 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4524, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1775);
   DLX_INST_DATA_PATH_DECODE_RF_U2056 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4523, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1776);
   DLX_INST_DATA_PATH_DECODE_RF_U2055 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4522, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1777);
   DLX_INST_DATA_PATH_DECODE_RF_U2054 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4521, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1778);
   DLX_INST_DATA_PATH_DECODE_RF_U2053 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4520, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1779);
   DLX_INST_DATA_PATH_DECODE_RF_U2052 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4519, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1780);
   DLX_INST_DATA_PATH_DECODE_RF_U2051 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4518, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1781);
   DLX_INST_DATA_PATH_DECODE_RF_U2050 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4517, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1782);
   DLX_INST_DATA_PATH_DECODE_RF_U2049 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5124, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1783);
   DLX_INST_DATA_PATH_DECODE_RF_U2048 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5123, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1784);
   DLX_INST_DATA_PATH_DECODE_RF_U2047 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5122, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1785);
   DLX_INST_DATA_PATH_DECODE_RF_U2046 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5121, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1786);
   DLX_INST_DATA_PATH_DECODE_RF_U2045 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5120, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1787);
   DLX_INST_DATA_PATH_DECODE_RF_U2044 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5119, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1788);
   DLX_INST_DATA_PATH_DECODE_RF_U2043 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5118, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1789);
   DLX_INST_DATA_PATH_DECODE_RF_U2042 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5117, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1790);
   DLX_INST_DATA_PATH_DECODE_RF_U2041 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5116, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1791);
   DLX_INST_DATA_PATH_DECODE_RF_U2040 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5115, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1792);
   DLX_INST_DATA_PATH_DECODE_RF_U2039 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5114, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1793);
   DLX_INST_DATA_PATH_DECODE_RF_U2038 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5113, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1794);
   DLX_INST_DATA_PATH_DECODE_RF_U2037 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5112, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1795);
   DLX_INST_DATA_PATH_DECODE_RF_U2036 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5111, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1796);
   DLX_INST_DATA_PATH_DECODE_RF_U2035 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5110, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1797);
   DLX_INST_DATA_PATH_DECODE_RF_U2034 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5109, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1798);
   DLX_INST_DATA_PATH_DECODE_RF_U2033 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5108, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1799);
   DLX_INST_DATA_PATH_DECODE_RF_U2032 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5107, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1800);
   DLX_INST_DATA_PATH_DECODE_RF_U2031 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5106, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1801);
   DLX_INST_DATA_PATH_DECODE_RF_U2030 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5105, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1802);
   DLX_INST_DATA_PATH_DECODE_RF_U2029 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5104, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1803);
   DLX_INST_DATA_PATH_DECODE_RF_U2028 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5103, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1804);
   DLX_INST_DATA_PATH_DECODE_RF_U2027 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5102, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1805);
   DLX_INST_DATA_PATH_DECODE_RF_U2026 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5101, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1806);
   DLX_INST_DATA_PATH_DECODE_RF_U2025 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5100, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1807);
   DLX_INST_DATA_PATH_DECODE_RF_U2024 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5099, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1808);
   DLX_INST_DATA_PATH_DECODE_RF_U2023 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5098, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1809);
   DLX_INST_DATA_PATH_DECODE_RF_U2022 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5097, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1810);
   DLX_INST_DATA_PATH_DECODE_RF_U2021 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5096, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1811);
   DLX_INST_DATA_PATH_DECODE_RF_U2020 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5095, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1812);
   DLX_INST_DATA_PATH_DECODE_RF_U2019 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5094, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1813);
   DLX_INST_DATA_PATH_DECODE_RF_U2018 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5093, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1814);
   DLX_INST_DATA_PATH_DECODE_RF_U2017 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n5, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6585);
   DLX_INST_DATA_PATH_DECODE_RF_U2016 : AND3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6586, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6585, A3 => 
                           DLX_INST_DATA_PATH_DECODE_n4, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6589);
   DLX_INST_DATA_PATH_DECODE_RF_U2015 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4868, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1815);
   DLX_INST_DATA_PATH_DECODE_RF_U2014 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4867, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1816);
   DLX_INST_DATA_PATH_DECODE_RF_U2013 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4866, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1817);
   DLX_INST_DATA_PATH_DECODE_RF_U2012 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4865, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1818);
   DLX_INST_DATA_PATH_DECODE_RF_U2011 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4864, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1819);
   DLX_INST_DATA_PATH_DECODE_RF_U2010 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4863, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1820);
   DLX_INST_DATA_PATH_DECODE_RF_U2009 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4862, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1821);
   DLX_INST_DATA_PATH_DECODE_RF_U2008 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4861, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1822);
   DLX_INST_DATA_PATH_DECODE_RF_U2007 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4860, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1823);
   DLX_INST_DATA_PATH_DECODE_RF_U2006 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4859, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1824);
   DLX_INST_DATA_PATH_DECODE_RF_U2005 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4858, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1825);
   DLX_INST_DATA_PATH_DECODE_RF_U2004 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4857, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1826);
   DLX_INST_DATA_PATH_DECODE_RF_U2003 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4856, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1827);
   DLX_INST_DATA_PATH_DECODE_RF_U2002 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4855, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1828);
   DLX_INST_DATA_PATH_DECODE_RF_U2001 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4854, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1829);
   DLX_INST_DATA_PATH_DECODE_RF_U2000 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4853, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1830);
   DLX_INST_DATA_PATH_DECODE_RF_U1999 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4852, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1831);
   DLX_INST_DATA_PATH_DECODE_RF_U1998 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4851, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1832);
   DLX_INST_DATA_PATH_DECODE_RF_U1997 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4850, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1833);
   DLX_INST_DATA_PATH_DECODE_RF_U1996 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4849, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1834);
   DLX_INST_DATA_PATH_DECODE_RF_U1995 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4848, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1835);
   DLX_INST_DATA_PATH_DECODE_RF_U1994 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4847, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1836);
   DLX_INST_DATA_PATH_DECODE_RF_U1993 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4846, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1837);
   DLX_INST_DATA_PATH_DECODE_RF_U1992 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4845, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1838);
   DLX_INST_DATA_PATH_DECODE_RF_U1991 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4844, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1839);
   DLX_INST_DATA_PATH_DECODE_RF_U1990 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4843, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1840);
   DLX_INST_DATA_PATH_DECODE_RF_U1989 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4842, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1841);
   DLX_INST_DATA_PATH_DECODE_RF_U1988 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4841, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1842);
   DLX_INST_DATA_PATH_DECODE_RF_U1987 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4840, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1843);
   DLX_INST_DATA_PATH_DECODE_RF_U1986 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4839, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1844);
   DLX_INST_DATA_PATH_DECODE_RF_U1985 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4838, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1845);
   DLX_INST_DATA_PATH_DECODE_RF_U1984 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4837, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1846);
   DLX_INST_DATA_PATH_DECODE_RF_U1983 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4482, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1847);
   DLX_INST_DATA_PATH_DECODE_RF_U1982 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4481, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1848);
   DLX_INST_DATA_PATH_DECODE_RF_U1981 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4480, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1849);
   DLX_INST_DATA_PATH_DECODE_RF_U1980 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4479, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1850);
   DLX_INST_DATA_PATH_DECODE_RF_U1979 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4478, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1851);
   DLX_INST_DATA_PATH_DECODE_RF_U1978 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4477, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1852);
   DLX_INST_DATA_PATH_DECODE_RF_U1977 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4476, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1853);
   DLX_INST_DATA_PATH_DECODE_RF_U1976 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4475, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1854);
   DLX_INST_DATA_PATH_DECODE_RF_U1975 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4474, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1855);
   DLX_INST_DATA_PATH_DECODE_RF_U1974 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4473, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1856);
   DLX_INST_DATA_PATH_DECODE_RF_U1973 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4472, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1857);
   DLX_INST_DATA_PATH_DECODE_RF_U1972 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4471, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1858);
   DLX_INST_DATA_PATH_DECODE_RF_U1971 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4470, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1859);
   DLX_INST_DATA_PATH_DECODE_RF_U1970 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4469, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1860);
   DLX_INST_DATA_PATH_DECODE_RF_U1969 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4468, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1861);
   DLX_INST_DATA_PATH_DECODE_RF_U1968 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4467, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1862);
   DLX_INST_DATA_PATH_DECODE_RF_U1967 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4466, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1863);
   DLX_INST_DATA_PATH_DECODE_RF_U1966 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4465, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1864);
   DLX_INST_DATA_PATH_DECODE_RF_U1965 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4464, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1865);
   DLX_INST_DATA_PATH_DECODE_RF_U1964 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4463, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1866);
   DLX_INST_DATA_PATH_DECODE_RF_U1963 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4462, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1867);
   DLX_INST_DATA_PATH_DECODE_RF_U1962 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4461, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1868);
   DLX_INST_DATA_PATH_DECODE_RF_U1961 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4460, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1869);
   DLX_INST_DATA_PATH_DECODE_RF_U1960 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4459, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1870);
   DLX_INST_DATA_PATH_DECODE_RF_U1959 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4458, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1871);
   DLX_INST_DATA_PATH_DECODE_RF_U1958 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4457, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1872);
   DLX_INST_DATA_PATH_DECODE_RF_U1957 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4456, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1873);
   DLX_INST_DATA_PATH_DECODE_RF_U1956 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4455, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1874);
   DLX_INST_DATA_PATH_DECODE_RF_U1955 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4454, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1875);
   DLX_INST_DATA_PATH_DECODE_RF_U1954 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4453, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1876);
   DLX_INST_DATA_PATH_DECODE_RF_U1953 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4452, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1877);
   DLX_INST_DATA_PATH_DECODE_RF_U1952 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4451, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1878);
   DLX_INST_DATA_PATH_DECODE_RF_U1951 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4740, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1879);
   DLX_INST_DATA_PATH_DECODE_RF_U1950 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4739, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1880);
   DLX_INST_DATA_PATH_DECODE_RF_U1949 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4738, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1881);
   DLX_INST_DATA_PATH_DECODE_RF_U1948 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4737, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1882);
   DLX_INST_DATA_PATH_DECODE_RF_U1947 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4736, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1883);
   DLX_INST_DATA_PATH_DECODE_RF_U1946 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4735, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1884);
   DLX_INST_DATA_PATH_DECODE_RF_U1945 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4734, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1885);
   DLX_INST_DATA_PATH_DECODE_RF_U1944 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4733, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1886);
   DLX_INST_DATA_PATH_DECODE_RF_U1943 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4732, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1887);
   DLX_INST_DATA_PATH_DECODE_RF_U1942 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4731, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1888);
   DLX_INST_DATA_PATH_DECODE_RF_U1941 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4730, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1889);
   DLX_INST_DATA_PATH_DECODE_RF_U1940 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4729, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1890);
   DLX_INST_DATA_PATH_DECODE_RF_U1939 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4728, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1891);
   DLX_INST_DATA_PATH_DECODE_RF_U1938 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4727, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1892);
   DLX_INST_DATA_PATH_DECODE_RF_U1937 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4726, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1893);
   DLX_INST_DATA_PATH_DECODE_RF_U1936 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4725, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1894);
   DLX_INST_DATA_PATH_DECODE_RF_U1935 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4724, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1895);
   DLX_INST_DATA_PATH_DECODE_RF_U1934 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4723, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1896);
   DLX_INST_DATA_PATH_DECODE_RF_U1933 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4722, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1897);
   DLX_INST_DATA_PATH_DECODE_RF_U1932 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4721, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1898);
   DLX_INST_DATA_PATH_DECODE_RF_U1931 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4720, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1899);
   DLX_INST_DATA_PATH_DECODE_RF_U1930 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4719, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1900);
   DLX_INST_DATA_PATH_DECODE_RF_U1929 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4718, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1901);
   DLX_INST_DATA_PATH_DECODE_RF_U1928 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4717, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1902);
   DLX_INST_DATA_PATH_DECODE_RF_U1927 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4716, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1903);
   DLX_INST_DATA_PATH_DECODE_RF_U1926 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4715, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1904);
   DLX_INST_DATA_PATH_DECODE_RF_U1925 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4714, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1905);
   DLX_INST_DATA_PATH_DECODE_RF_U1924 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4713, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1906);
   DLX_INST_DATA_PATH_DECODE_RF_U1923 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4712, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1907);
   DLX_INST_DATA_PATH_DECODE_RF_U1922 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4711, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1908);
   DLX_INST_DATA_PATH_DECODE_RF_U1921 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4710, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1909);
   DLX_INST_DATA_PATH_DECODE_RF_U1920 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4709, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1910);
   DLX_INST_DATA_PATH_DECODE_RF_U1919 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5092, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1911);
   DLX_INST_DATA_PATH_DECODE_RF_U1918 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5091, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1912);
   DLX_INST_DATA_PATH_DECODE_RF_U1917 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5090, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1913);
   DLX_INST_DATA_PATH_DECODE_RF_U1916 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5089, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1914);
   DLX_INST_DATA_PATH_DECODE_RF_U1915 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5088, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1915);
   DLX_INST_DATA_PATH_DECODE_RF_U1914 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5087, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1916);
   DLX_INST_DATA_PATH_DECODE_RF_U1913 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5086, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1917);
   DLX_INST_DATA_PATH_DECODE_RF_U1912 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5085, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1918);
   DLX_INST_DATA_PATH_DECODE_RF_U1911 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5084, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1919);
   DLX_INST_DATA_PATH_DECODE_RF_U1910 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5083, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1920);
   DLX_INST_DATA_PATH_DECODE_RF_U1909 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5082, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1921);
   DLX_INST_DATA_PATH_DECODE_RF_U1908 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5081, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1922);
   DLX_INST_DATA_PATH_DECODE_RF_U1907 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5080, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1923);
   DLX_INST_DATA_PATH_DECODE_RF_U1906 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5079, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1924);
   DLX_INST_DATA_PATH_DECODE_RF_U1905 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5078, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1925);
   DLX_INST_DATA_PATH_DECODE_RF_U1904 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5077, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1926);
   DLX_INST_DATA_PATH_DECODE_RF_U1903 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5076, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1927);
   DLX_INST_DATA_PATH_DECODE_RF_U1902 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5075, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1928);
   DLX_INST_DATA_PATH_DECODE_RF_U1901 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5074, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1929);
   DLX_INST_DATA_PATH_DECODE_RF_U1900 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5073, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1930);
   DLX_INST_DATA_PATH_DECODE_RF_U1899 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5072, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1931);
   DLX_INST_DATA_PATH_DECODE_RF_U1898 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5071, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1932);
   DLX_INST_DATA_PATH_DECODE_RF_U1897 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5070, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1933);
   DLX_INST_DATA_PATH_DECODE_RF_U1896 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5069, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1934);
   DLX_INST_DATA_PATH_DECODE_RF_U1895 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5068, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1935);
   DLX_INST_DATA_PATH_DECODE_RF_U1894 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5067, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1936);
   DLX_INST_DATA_PATH_DECODE_RF_U1893 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5066, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1937);
   DLX_INST_DATA_PATH_DECODE_RF_U1892 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5065, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1938);
   DLX_INST_DATA_PATH_DECODE_RF_U1891 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5064, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1939);
   DLX_INST_DATA_PATH_DECODE_RF_U1890 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5063, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1940);
   DLX_INST_DATA_PATH_DECODE_RF_U1889 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5062, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1941);
   DLX_INST_DATA_PATH_DECODE_RF_U1888 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5061, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1942);
   DLX_INST_DATA_PATH_DECODE_RF_U1887 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5060, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1943);
   DLX_INST_DATA_PATH_DECODE_RF_U1886 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5059, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1944);
   DLX_INST_DATA_PATH_DECODE_RF_U1885 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5058, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1945);
   DLX_INST_DATA_PATH_DECODE_RF_U1884 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5057, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1946);
   DLX_INST_DATA_PATH_DECODE_RF_U1883 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5056, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1947);
   DLX_INST_DATA_PATH_DECODE_RF_U1882 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5055, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1948);
   DLX_INST_DATA_PATH_DECODE_RF_U1881 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5054, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1949);
   DLX_INST_DATA_PATH_DECODE_RF_U1880 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5053, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1950);
   DLX_INST_DATA_PATH_DECODE_RF_U1879 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5052, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1951);
   DLX_INST_DATA_PATH_DECODE_RF_U1878 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5051, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1952);
   DLX_INST_DATA_PATH_DECODE_RF_U1877 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5050, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1953);
   DLX_INST_DATA_PATH_DECODE_RF_U1876 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5049, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1954);
   DLX_INST_DATA_PATH_DECODE_RF_U1875 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5048, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1955);
   DLX_INST_DATA_PATH_DECODE_RF_U1874 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5047, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1956);
   DLX_INST_DATA_PATH_DECODE_RF_U1873 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5046, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1957);
   DLX_INST_DATA_PATH_DECODE_RF_U1872 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5045, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1958);
   DLX_INST_DATA_PATH_DECODE_RF_U1871 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5044, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1959);
   DLX_INST_DATA_PATH_DECODE_RF_U1870 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5043, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1960);
   DLX_INST_DATA_PATH_DECODE_RF_U1869 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5042, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1961);
   DLX_INST_DATA_PATH_DECODE_RF_U1868 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5041, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1962);
   DLX_INST_DATA_PATH_DECODE_RF_U1867 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5040, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1963);
   DLX_INST_DATA_PATH_DECODE_RF_U1866 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5039, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1964);
   DLX_INST_DATA_PATH_DECODE_RF_U1865 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5038, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1965);
   DLX_INST_DATA_PATH_DECODE_RF_U1864 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5037, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1966);
   DLX_INST_DATA_PATH_DECODE_RF_U1863 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5036, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1967);
   DLX_INST_DATA_PATH_DECODE_RF_U1862 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5035, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1968);
   DLX_INST_DATA_PATH_DECODE_RF_U1861 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5034, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1969);
   DLX_INST_DATA_PATH_DECODE_RF_U1860 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5033, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1970);
   DLX_INST_DATA_PATH_DECODE_RF_U1859 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5032, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1971);
   DLX_INST_DATA_PATH_DECODE_RF_U1858 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5031, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1972);
   DLX_INST_DATA_PATH_DECODE_RF_U1857 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5030, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1973);
   DLX_INST_DATA_PATH_DECODE_RF_U1856 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5029, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1974);
   DLX_INST_DATA_PATH_DECODE_RF_U1855 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4226, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1975);
   DLX_INST_DATA_PATH_DECODE_RF_U1854 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4225, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1976);
   DLX_INST_DATA_PATH_DECODE_RF_U1853 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4224, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1977);
   DLX_INST_DATA_PATH_DECODE_RF_U1852 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4223, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1978);
   DLX_INST_DATA_PATH_DECODE_RF_U1851 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4222, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1979);
   DLX_INST_DATA_PATH_DECODE_RF_U1850 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4221, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1980);
   DLX_INST_DATA_PATH_DECODE_RF_U1849 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4220, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1981);
   DLX_INST_DATA_PATH_DECODE_RF_U1848 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4219, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1982);
   DLX_INST_DATA_PATH_DECODE_RF_U1847 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4218, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1983);
   DLX_INST_DATA_PATH_DECODE_RF_U1846 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4217, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1984);
   DLX_INST_DATA_PATH_DECODE_RF_U1845 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4216, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1985);
   DLX_INST_DATA_PATH_DECODE_RF_U1844 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4215, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1986);
   DLX_INST_DATA_PATH_DECODE_RF_U1843 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4214, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1987);
   DLX_INST_DATA_PATH_DECODE_RF_U1842 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4213, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1988);
   DLX_INST_DATA_PATH_DECODE_RF_U1841 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4212, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1989);
   DLX_INST_DATA_PATH_DECODE_RF_U1840 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4211, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1990);
   DLX_INST_DATA_PATH_DECODE_RF_U1839 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4210, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1991);
   DLX_INST_DATA_PATH_DECODE_RF_U1838 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4209, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1992);
   DLX_INST_DATA_PATH_DECODE_RF_U1837 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4208, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1993);
   DLX_INST_DATA_PATH_DECODE_RF_U1836 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4207, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1994);
   DLX_INST_DATA_PATH_DECODE_RF_U1835 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4206, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1995);
   DLX_INST_DATA_PATH_DECODE_RF_U1834 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4205, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1996);
   DLX_INST_DATA_PATH_DECODE_RF_U1833 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4204, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1997);
   DLX_INST_DATA_PATH_DECODE_RF_U1832 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4203, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1998);
   DLX_INST_DATA_PATH_DECODE_RF_U1831 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4202, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n1999);
   DLX_INST_DATA_PATH_DECODE_RF_U1830 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4201, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2000);
   DLX_INST_DATA_PATH_DECODE_RF_U1829 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4200, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2001);
   DLX_INST_DATA_PATH_DECODE_RF_U1828 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4199, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2002);
   DLX_INST_DATA_PATH_DECODE_RF_U1827 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4198, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2003);
   DLX_INST_DATA_PATH_DECODE_RF_U1826 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4197, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2004);
   DLX_INST_DATA_PATH_DECODE_RF_U1825 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4196, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2005);
   DLX_INST_DATA_PATH_DECODE_RF_U1824 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4195, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2006);
   DLX_INST_DATA_PATH_DECODE_RF_U1823 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4258, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2007);
   DLX_INST_DATA_PATH_DECODE_RF_U1822 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4257, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2008);
   DLX_INST_DATA_PATH_DECODE_RF_U1821 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4256, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2009);
   DLX_INST_DATA_PATH_DECODE_RF_U1820 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4255, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2010);
   DLX_INST_DATA_PATH_DECODE_RF_U1819 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4254, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2011);
   DLX_INST_DATA_PATH_DECODE_RF_U1818 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4253, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2012);
   DLX_INST_DATA_PATH_DECODE_RF_U1817 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4252, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2013);
   DLX_INST_DATA_PATH_DECODE_RF_U1816 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4251, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2014);
   DLX_INST_DATA_PATH_DECODE_RF_U1815 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4250, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2015);
   DLX_INST_DATA_PATH_DECODE_RF_U1814 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4249, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2016);
   DLX_INST_DATA_PATH_DECODE_RF_U1813 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4248, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2017);
   DLX_INST_DATA_PATH_DECODE_RF_U1812 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4247, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2018);
   DLX_INST_DATA_PATH_DECODE_RF_U1811 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4246, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2019);
   DLX_INST_DATA_PATH_DECODE_RF_U1810 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4245, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2020);
   DLX_INST_DATA_PATH_DECODE_RF_U1809 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4244, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2021);
   DLX_INST_DATA_PATH_DECODE_RF_U1808 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4243, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2022);
   DLX_INST_DATA_PATH_DECODE_RF_U1807 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4242, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2023);
   DLX_INST_DATA_PATH_DECODE_RF_U1806 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4241, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2024);
   DLX_INST_DATA_PATH_DECODE_RF_U1805 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4240, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2025);
   DLX_INST_DATA_PATH_DECODE_RF_U1804 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4239, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2026);
   DLX_INST_DATA_PATH_DECODE_RF_U1803 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4238, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2027);
   DLX_INST_DATA_PATH_DECODE_RF_U1802 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4237, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2028);
   DLX_INST_DATA_PATH_DECODE_RF_U1801 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4236, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2029);
   DLX_INST_DATA_PATH_DECODE_RF_U1800 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4235, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2030);
   DLX_INST_DATA_PATH_DECODE_RF_U1799 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4234, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2031);
   DLX_INST_DATA_PATH_DECODE_RF_U1798 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4233, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2032);
   DLX_INST_DATA_PATH_DECODE_RF_U1797 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4232, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2033);
   DLX_INST_DATA_PATH_DECODE_RF_U1796 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4231, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2034);
   DLX_INST_DATA_PATH_DECODE_RF_U1795 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4230, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2035);
   DLX_INST_DATA_PATH_DECODE_RF_U1794 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4229, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2036);
   DLX_INST_DATA_PATH_DECODE_RF_U1793 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4228, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2037);
   DLX_INST_DATA_PATH_DECODE_RF_U1792 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4227, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2038);
   DLX_INST_DATA_PATH_DECODE_RF_U1791 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4836, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2039);
   DLX_INST_DATA_PATH_DECODE_RF_U1790 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4835, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2040);
   DLX_INST_DATA_PATH_DECODE_RF_U1789 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4834, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2041);
   DLX_INST_DATA_PATH_DECODE_RF_U1788 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4833, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2042);
   DLX_INST_DATA_PATH_DECODE_RF_U1787 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4832, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2043);
   DLX_INST_DATA_PATH_DECODE_RF_U1786 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4831, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2044);
   DLX_INST_DATA_PATH_DECODE_RF_U1785 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4830, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2045);
   DLX_INST_DATA_PATH_DECODE_RF_U1784 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4829, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2046);
   DLX_INST_DATA_PATH_DECODE_RF_U1783 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4828, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2047);
   DLX_INST_DATA_PATH_DECODE_RF_U1782 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4827, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2048);
   DLX_INST_DATA_PATH_DECODE_RF_U1781 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4826, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2049);
   DLX_INST_DATA_PATH_DECODE_RF_U1780 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4825, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2050);
   DLX_INST_DATA_PATH_DECODE_RF_U1779 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4824, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2051);
   DLX_INST_DATA_PATH_DECODE_RF_U1778 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4823, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2052);
   DLX_INST_DATA_PATH_DECODE_RF_U1777 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4822, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2053);
   DLX_INST_DATA_PATH_DECODE_RF_U1776 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4821, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2054);
   DLX_INST_DATA_PATH_DECODE_RF_U1775 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4820, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2055);
   DLX_INST_DATA_PATH_DECODE_RF_U1774 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4819, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2056);
   DLX_INST_DATA_PATH_DECODE_RF_U1773 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4818, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2057);
   DLX_INST_DATA_PATH_DECODE_RF_U1772 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4817, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2058);
   DLX_INST_DATA_PATH_DECODE_RF_U1771 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4816, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2059);
   DLX_INST_DATA_PATH_DECODE_RF_U1770 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4815, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2060);
   DLX_INST_DATA_PATH_DECODE_RF_U1769 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4814, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2061);
   DLX_INST_DATA_PATH_DECODE_RF_U1768 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4813, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2062);
   DLX_INST_DATA_PATH_DECODE_RF_U1767 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4812, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2063);
   DLX_INST_DATA_PATH_DECODE_RF_U1766 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4811, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2064);
   DLX_INST_DATA_PATH_DECODE_RF_U1765 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4810, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2065);
   DLX_INST_DATA_PATH_DECODE_RF_U1764 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4809, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2066);
   DLX_INST_DATA_PATH_DECODE_RF_U1763 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4808, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2067);
   DLX_INST_DATA_PATH_DECODE_RF_U1762 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4807, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2068);
   DLX_INST_DATA_PATH_DECODE_RF_U1761 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4806, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2069);
   DLX_INST_DATA_PATH_DECODE_RF_U1760 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4805, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2070);
   DLX_INST_DATA_PATH_DECODE_RF_U1759 : AND3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6584, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6585, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6586, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6562);
   DLX_INST_DATA_PATH_DECODE_RF_U1758 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4450, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2071);
   DLX_INST_DATA_PATH_DECODE_RF_U1757 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4449, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2072);
   DLX_INST_DATA_PATH_DECODE_RF_U1756 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4448, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2073);
   DLX_INST_DATA_PATH_DECODE_RF_U1755 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4447, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2074);
   DLX_INST_DATA_PATH_DECODE_RF_U1754 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4446, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2075);
   DLX_INST_DATA_PATH_DECODE_RF_U1753 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4445, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2076);
   DLX_INST_DATA_PATH_DECODE_RF_U1752 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4444, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2077);
   DLX_INST_DATA_PATH_DECODE_RF_U1751 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4443, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2078);
   DLX_INST_DATA_PATH_DECODE_RF_U1750 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4442, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2079);
   DLX_INST_DATA_PATH_DECODE_RF_U1749 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4441, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2080);
   DLX_INST_DATA_PATH_DECODE_RF_U1748 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4440, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2081);
   DLX_INST_DATA_PATH_DECODE_RF_U1747 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4439, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2082);
   DLX_INST_DATA_PATH_DECODE_RF_U1746 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4438, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2083);
   DLX_INST_DATA_PATH_DECODE_RF_U1745 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4437, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2084);
   DLX_INST_DATA_PATH_DECODE_RF_U1744 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4436, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2085);
   DLX_INST_DATA_PATH_DECODE_RF_U1743 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4435, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2086);
   DLX_INST_DATA_PATH_DECODE_RF_U1742 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4434, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2087);
   DLX_INST_DATA_PATH_DECODE_RF_U1741 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4433, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2088);
   DLX_INST_DATA_PATH_DECODE_RF_U1740 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4432, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2089);
   DLX_INST_DATA_PATH_DECODE_RF_U1739 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4431, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2090);
   DLX_INST_DATA_PATH_DECODE_RF_U1738 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4430, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2091);
   DLX_INST_DATA_PATH_DECODE_RF_U1737 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4429, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2092);
   DLX_INST_DATA_PATH_DECODE_RF_U1736 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4428, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2093);
   DLX_INST_DATA_PATH_DECODE_RF_U1735 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4427, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2094);
   DLX_INST_DATA_PATH_DECODE_RF_U1734 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4426, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2095);
   DLX_INST_DATA_PATH_DECODE_RF_U1733 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4425, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2096);
   DLX_INST_DATA_PATH_DECODE_RF_U1732 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4424, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2097);
   DLX_INST_DATA_PATH_DECODE_RF_U1731 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4423, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2098);
   DLX_INST_DATA_PATH_DECODE_RF_U1730 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4422, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2099);
   DLX_INST_DATA_PATH_DECODE_RF_U1729 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4421, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2100);
   DLX_INST_DATA_PATH_DECODE_RF_U1728 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4420, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2101);
   DLX_INST_DATA_PATH_DECODE_RF_U1727 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4419, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2102);
   DLX_INST_DATA_PATH_DECODE_RF_U1726 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4708, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2103);
   DLX_INST_DATA_PATH_DECODE_RF_U1725 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4707, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2104);
   DLX_INST_DATA_PATH_DECODE_RF_U1724 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4706, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2105);
   DLX_INST_DATA_PATH_DECODE_RF_U1723 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4705, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2106);
   DLX_INST_DATA_PATH_DECODE_RF_U1722 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4704, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2107);
   DLX_INST_DATA_PATH_DECODE_RF_U1721 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4703, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2108);
   DLX_INST_DATA_PATH_DECODE_RF_U1720 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4702, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2109);
   DLX_INST_DATA_PATH_DECODE_RF_U1719 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4701, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2110);
   DLX_INST_DATA_PATH_DECODE_RF_U1718 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4700, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2111);
   DLX_INST_DATA_PATH_DECODE_RF_U1717 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4699, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2112);
   DLX_INST_DATA_PATH_DECODE_RF_U1716 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4698, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2113);
   DLX_INST_DATA_PATH_DECODE_RF_U1715 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4697, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2114);
   DLX_INST_DATA_PATH_DECODE_RF_U1714 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4696, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2115);
   DLX_INST_DATA_PATH_DECODE_RF_U1713 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4695, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2116);
   DLX_INST_DATA_PATH_DECODE_RF_U1712 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4694, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2117);
   DLX_INST_DATA_PATH_DECODE_RF_U1711 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4693, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2118);
   DLX_INST_DATA_PATH_DECODE_RF_U1710 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4692, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2119);
   DLX_INST_DATA_PATH_DECODE_RF_U1709 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4691, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2120);
   DLX_INST_DATA_PATH_DECODE_RF_U1708 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4690, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2121);
   DLX_INST_DATA_PATH_DECODE_RF_U1707 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4689, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2122);
   DLX_INST_DATA_PATH_DECODE_RF_U1706 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4688, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2123);
   DLX_INST_DATA_PATH_DECODE_RF_U1705 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4687, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2124);
   DLX_INST_DATA_PATH_DECODE_RF_U1704 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4686, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2125);
   DLX_INST_DATA_PATH_DECODE_RF_U1703 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4685, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2126);
   DLX_INST_DATA_PATH_DECODE_RF_U1702 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4684, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2127);
   DLX_INST_DATA_PATH_DECODE_RF_U1701 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4683, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2128);
   DLX_INST_DATA_PATH_DECODE_RF_U1700 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4682, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2129);
   DLX_INST_DATA_PATH_DECODE_RF_U1699 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4681, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2130);
   DLX_INST_DATA_PATH_DECODE_RF_U1698 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4680, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2131);
   DLX_INST_DATA_PATH_DECODE_RF_U1697 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4679, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2132);
   DLX_INST_DATA_PATH_DECODE_RF_U1696 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4678, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2133);
   DLX_INST_DATA_PATH_DECODE_RF_U1695 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4677, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2134);
   DLX_INST_DATA_PATH_DECODE_RF_U1694 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4194, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2135);
   DLX_INST_DATA_PATH_DECODE_RF_U1693 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4193, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2136);
   DLX_INST_DATA_PATH_DECODE_RF_U1692 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4192, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2137);
   DLX_INST_DATA_PATH_DECODE_RF_U1691 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4191, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2138);
   DLX_INST_DATA_PATH_DECODE_RF_U1690 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4190, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2139);
   DLX_INST_DATA_PATH_DECODE_RF_U1689 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4189, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2140);
   DLX_INST_DATA_PATH_DECODE_RF_U1688 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4188, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2141);
   DLX_INST_DATA_PATH_DECODE_RF_U1687 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4187, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2142);
   DLX_INST_DATA_PATH_DECODE_RF_U1686 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4186, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2143);
   DLX_INST_DATA_PATH_DECODE_RF_U1685 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4185, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2144);
   DLX_INST_DATA_PATH_DECODE_RF_U1684 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4184, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2145);
   DLX_INST_DATA_PATH_DECODE_RF_U1683 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4183, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2146);
   DLX_INST_DATA_PATH_DECODE_RF_U1682 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4182, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2147);
   DLX_INST_DATA_PATH_DECODE_RF_U1681 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4181, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2148);
   DLX_INST_DATA_PATH_DECODE_RF_U1680 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4180, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2149);
   DLX_INST_DATA_PATH_DECODE_RF_U1679 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4179, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2150);
   DLX_INST_DATA_PATH_DECODE_RF_U1678 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4178, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2151);
   DLX_INST_DATA_PATH_DECODE_RF_U1677 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4177, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2152);
   DLX_INST_DATA_PATH_DECODE_RF_U1676 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4176, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2153);
   DLX_INST_DATA_PATH_DECODE_RF_U1675 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4175, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2154);
   DLX_INST_DATA_PATH_DECODE_RF_U1674 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4174, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2155);
   DLX_INST_DATA_PATH_DECODE_RF_U1673 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4173, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2156);
   DLX_INST_DATA_PATH_DECODE_RF_U1672 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4172, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2157);
   DLX_INST_DATA_PATH_DECODE_RF_U1671 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4171, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2158);
   DLX_INST_DATA_PATH_DECODE_RF_U1670 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4170, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2159);
   DLX_INST_DATA_PATH_DECODE_RF_U1669 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4169, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2160);
   DLX_INST_DATA_PATH_DECODE_RF_U1668 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4168, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2161);
   DLX_INST_DATA_PATH_DECODE_RF_U1667 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4167, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2162);
   DLX_INST_DATA_PATH_DECODE_RF_U1666 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4166, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2163);
   DLX_INST_DATA_PATH_DECODE_RF_U1665 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4165, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2164);
   DLX_INST_DATA_PATH_DECODE_RF_U1664 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4164, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2165);
   DLX_INST_DATA_PATH_DECODE_RF_U1663 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4163, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2166);
   DLX_INST_DATA_PATH_DECODE_RF_U1662 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4804, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2167);
   DLX_INST_DATA_PATH_DECODE_RF_U1661 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4803, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2168);
   DLX_INST_DATA_PATH_DECODE_RF_U1660 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4802, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2169);
   DLX_INST_DATA_PATH_DECODE_RF_U1659 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4801, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2170);
   DLX_INST_DATA_PATH_DECODE_RF_U1658 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4800, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2171);
   DLX_INST_DATA_PATH_DECODE_RF_U1657 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4799, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2172);
   DLX_INST_DATA_PATH_DECODE_RF_U1656 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4798, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2173);
   DLX_INST_DATA_PATH_DECODE_RF_U1655 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4797, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2174);
   DLX_INST_DATA_PATH_DECODE_RF_U1654 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4796, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2175);
   DLX_INST_DATA_PATH_DECODE_RF_U1653 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4795, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2176);
   DLX_INST_DATA_PATH_DECODE_RF_U1652 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4794, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2177);
   DLX_INST_DATA_PATH_DECODE_RF_U1651 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4793, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2178);
   DLX_INST_DATA_PATH_DECODE_RF_U1650 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4792, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2179);
   DLX_INST_DATA_PATH_DECODE_RF_U1649 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4791, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2180);
   DLX_INST_DATA_PATH_DECODE_RF_U1648 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4790, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2181);
   DLX_INST_DATA_PATH_DECODE_RF_U1647 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4789, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2182);
   DLX_INST_DATA_PATH_DECODE_RF_U1646 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4788, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2183);
   DLX_INST_DATA_PATH_DECODE_RF_U1645 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4787, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2184);
   DLX_INST_DATA_PATH_DECODE_RF_U1644 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4786, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2185);
   DLX_INST_DATA_PATH_DECODE_RF_U1643 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4785, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2186);
   DLX_INST_DATA_PATH_DECODE_RF_U1642 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4784, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2187);
   DLX_INST_DATA_PATH_DECODE_RF_U1641 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4783, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2188);
   DLX_INST_DATA_PATH_DECODE_RF_U1640 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4782, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2189);
   DLX_INST_DATA_PATH_DECODE_RF_U1639 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4781, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2190);
   DLX_INST_DATA_PATH_DECODE_RF_U1638 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4780, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2191);
   DLX_INST_DATA_PATH_DECODE_RF_U1637 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4779, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2192);
   DLX_INST_DATA_PATH_DECODE_RF_U1636 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4778, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2193);
   DLX_INST_DATA_PATH_DECODE_RF_U1635 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4777, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2194);
   DLX_INST_DATA_PATH_DECODE_RF_U1634 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4776, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2195);
   DLX_INST_DATA_PATH_DECODE_RF_U1633 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4775, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2196);
   DLX_INST_DATA_PATH_DECODE_RF_U1632 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4774, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2197);
   DLX_INST_DATA_PATH_DECODE_RF_U1631 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4773, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2198);
   DLX_INST_DATA_PATH_DECODE_RF_U1630 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4772, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2199);
   DLX_INST_DATA_PATH_DECODE_RF_U1629 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4771, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2200);
   DLX_INST_DATA_PATH_DECODE_RF_U1628 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4770, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2201);
   DLX_INST_DATA_PATH_DECODE_RF_U1627 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4769, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2202);
   DLX_INST_DATA_PATH_DECODE_RF_U1626 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4768, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2203);
   DLX_INST_DATA_PATH_DECODE_RF_U1625 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4767, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2204);
   DLX_INST_DATA_PATH_DECODE_RF_U1624 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4766, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2205);
   DLX_INST_DATA_PATH_DECODE_RF_U1623 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4765, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2206);
   DLX_INST_DATA_PATH_DECODE_RF_U1622 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4764, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2207);
   DLX_INST_DATA_PATH_DECODE_RF_U1621 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4763, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2208);
   DLX_INST_DATA_PATH_DECODE_RF_U1620 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4762, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2209);
   DLX_INST_DATA_PATH_DECODE_RF_U1619 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4761, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2210);
   DLX_INST_DATA_PATH_DECODE_RF_U1618 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4760, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2211);
   DLX_INST_DATA_PATH_DECODE_RF_U1617 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4759, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2212);
   DLX_INST_DATA_PATH_DECODE_RF_U1616 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4758, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2213);
   DLX_INST_DATA_PATH_DECODE_RF_U1615 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4757, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2214);
   DLX_INST_DATA_PATH_DECODE_RF_U1614 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4756, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2215);
   DLX_INST_DATA_PATH_DECODE_RF_U1613 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4755, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2216);
   DLX_INST_DATA_PATH_DECODE_RF_U1612 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4754, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2217);
   DLX_INST_DATA_PATH_DECODE_RF_U1611 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4753, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2218);
   DLX_INST_DATA_PATH_DECODE_RF_U1610 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4752, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2219);
   DLX_INST_DATA_PATH_DECODE_RF_U1609 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4751, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2220);
   DLX_INST_DATA_PATH_DECODE_RF_U1608 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4750, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2221);
   DLX_INST_DATA_PATH_DECODE_RF_U1607 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4749, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2222);
   DLX_INST_DATA_PATH_DECODE_RF_U1606 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4748, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2223);
   DLX_INST_DATA_PATH_DECODE_RF_U1605 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4747, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2224);
   DLX_INST_DATA_PATH_DECODE_RF_U1604 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4746, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2225);
   DLX_INST_DATA_PATH_DECODE_RF_U1603 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4745, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2226);
   DLX_INST_DATA_PATH_DECODE_RF_U1602 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4744, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2227);
   DLX_INST_DATA_PATH_DECODE_RF_U1601 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4743, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2228);
   DLX_INST_DATA_PATH_DECODE_RF_U1600 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4742, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2229);
   DLX_INST_DATA_PATH_DECODE_RF_U1599 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4741, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2230);
   DLX_INST_DATA_PATH_DECODE_RF_U1598 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5028, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2231);
   DLX_INST_DATA_PATH_DECODE_RF_U1597 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5027, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2232);
   DLX_INST_DATA_PATH_DECODE_RF_U1596 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5026, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2233);
   DLX_INST_DATA_PATH_DECODE_RF_U1595 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5025, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2234);
   DLX_INST_DATA_PATH_DECODE_RF_U1594 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5024, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2235);
   DLX_INST_DATA_PATH_DECODE_RF_U1593 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5023, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2236);
   DLX_INST_DATA_PATH_DECODE_RF_U1592 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5022, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2237);
   DLX_INST_DATA_PATH_DECODE_RF_U1591 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5021, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2238);
   DLX_INST_DATA_PATH_DECODE_RF_U1590 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5020, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2239);
   DLX_INST_DATA_PATH_DECODE_RF_U1589 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5019, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2240);
   DLX_INST_DATA_PATH_DECODE_RF_U1588 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5018, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2241);
   DLX_INST_DATA_PATH_DECODE_RF_U1587 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5017, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2242);
   DLX_INST_DATA_PATH_DECODE_RF_U1586 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5016, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2243);
   DLX_INST_DATA_PATH_DECODE_RF_U1585 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5015, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2244);
   DLX_INST_DATA_PATH_DECODE_RF_U1584 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5014, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2245);
   DLX_INST_DATA_PATH_DECODE_RF_U1583 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5013, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2246);
   DLX_INST_DATA_PATH_DECODE_RF_U1582 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5012, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2247);
   DLX_INST_DATA_PATH_DECODE_RF_U1581 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5011, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2248);
   DLX_INST_DATA_PATH_DECODE_RF_U1580 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5010, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2249);
   DLX_INST_DATA_PATH_DECODE_RF_U1579 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5009, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2250);
   DLX_INST_DATA_PATH_DECODE_RF_U1578 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5008, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2251);
   DLX_INST_DATA_PATH_DECODE_RF_U1577 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5007, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2252);
   DLX_INST_DATA_PATH_DECODE_RF_U1576 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5006, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2253);
   DLX_INST_DATA_PATH_DECODE_RF_U1575 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5005, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2254);
   DLX_INST_DATA_PATH_DECODE_RF_U1574 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5004, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2255);
   DLX_INST_DATA_PATH_DECODE_RF_U1573 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5003, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2256);
   DLX_INST_DATA_PATH_DECODE_RF_U1572 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5002, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2257);
   DLX_INST_DATA_PATH_DECODE_RF_U1571 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5001, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2258);
   DLX_INST_DATA_PATH_DECODE_RF_U1570 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5000, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2259);
   DLX_INST_DATA_PATH_DECODE_RF_U1569 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4999, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2260);
   DLX_INST_DATA_PATH_DECODE_RF_U1568 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4998, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2261);
   DLX_INST_DATA_PATH_DECODE_RF_U1567 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4997, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2262);
   DLX_INST_DATA_PATH_DECODE_RF_U1566 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4996, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2263);
   DLX_INST_DATA_PATH_DECODE_RF_U1565 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4995, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2264);
   DLX_INST_DATA_PATH_DECODE_RF_U1564 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4994, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2265);
   DLX_INST_DATA_PATH_DECODE_RF_U1563 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4993, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2266);
   DLX_INST_DATA_PATH_DECODE_RF_U1562 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4992, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2267);
   DLX_INST_DATA_PATH_DECODE_RF_U1561 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4991, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2268);
   DLX_INST_DATA_PATH_DECODE_RF_U1560 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4990, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2269);
   DLX_INST_DATA_PATH_DECODE_RF_U1559 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4989, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2270);
   DLX_INST_DATA_PATH_DECODE_RF_U1558 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4988, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2271);
   DLX_INST_DATA_PATH_DECODE_RF_U1557 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4987, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2272);
   DLX_INST_DATA_PATH_DECODE_RF_U1556 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4986, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2273);
   DLX_INST_DATA_PATH_DECODE_RF_U1555 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4985, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2274);
   DLX_INST_DATA_PATH_DECODE_RF_U1554 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4984, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2275);
   DLX_INST_DATA_PATH_DECODE_RF_U1553 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4983, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2276);
   DLX_INST_DATA_PATH_DECODE_RF_U1552 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4982, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2277);
   DLX_INST_DATA_PATH_DECODE_RF_U1551 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4981, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2278);
   DLX_INST_DATA_PATH_DECODE_RF_U1550 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4980, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2279);
   DLX_INST_DATA_PATH_DECODE_RF_U1549 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4979, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2280);
   DLX_INST_DATA_PATH_DECODE_RF_U1548 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2281);
   DLX_INST_DATA_PATH_DECODE_RF_U1547 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4977, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2282);
   DLX_INST_DATA_PATH_DECODE_RF_U1546 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4976, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2283);
   DLX_INST_DATA_PATH_DECODE_RF_U1545 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4975, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2284);
   DLX_INST_DATA_PATH_DECODE_RF_U1544 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4974, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2285);
   DLX_INST_DATA_PATH_DECODE_RF_U1543 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4973, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2286);
   DLX_INST_DATA_PATH_DECODE_RF_U1542 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2287);
   DLX_INST_DATA_PATH_DECODE_RF_U1541 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4971, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2288);
   DLX_INST_DATA_PATH_DECODE_RF_U1540 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4970, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2289);
   DLX_INST_DATA_PATH_DECODE_RF_U1539 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4969, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2290);
   DLX_INST_DATA_PATH_DECODE_RF_U1538 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4968, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2291);
   DLX_INST_DATA_PATH_DECODE_RF_U1537 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2292);
   DLX_INST_DATA_PATH_DECODE_RF_U1536 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4966, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2293);
   DLX_INST_DATA_PATH_DECODE_RF_U1535 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4965, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2294);
   DLX_INST_DATA_PATH_DECODE_RF_U1534 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4516, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2295);
   DLX_INST_DATA_PATH_DECODE_RF_U1533 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4515, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2296);
   DLX_INST_DATA_PATH_DECODE_RF_U1532 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4514, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2297);
   DLX_INST_DATA_PATH_DECODE_RF_U1531 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4513, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2298);
   DLX_INST_DATA_PATH_DECODE_RF_U1530 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4512, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2299);
   DLX_INST_DATA_PATH_DECODE_RF_U1529 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4511, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2300);
   DLX_INST_DATA_PATH_DECODE_RF_U1528 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4510, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2301);
   DLX_INST_DATA_PATH_DECODE_RF_U1527 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4509, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2302);
   DLX_INST_DATA_PATH_DECODE_RF_U1526 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4508, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2303);
   DLX_INST_DATA_PATH_DECODE_RF_U1525 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4507, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2304);
   DLX_INST_DATA_PATH_DECODE_RF_U1524 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4506, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2305);
   DLX_INST_DATA_PATH_DECODE_RF_U1523 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4505, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2306);
   DLX_INST_DATA_PATH_DECODE_RF_U1522 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4504, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2307);
   DLX_INST_DATA_PATH_DECODE_RF_U1521 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4503, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2308);
   DLX_INST_DATA_PATH_DECODE_RF_U1520 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4502, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2309);
   DLX_INST_DATA_PATH_DECODE_RF_U1519 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4501, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2310);
   DLX_INST_DATA_PATH_DECODE_RF_U1518 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4500, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2311);
   DLX_INST_DATA_PATH_DECODE_RF_U1517 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4499, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2312);
   DLX_INST_DATA_PATH_DECODE_RF_U1516 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4498, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2313);
   DLX_INST_DATA_PATH_DECODE_RF_U1515 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4497, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2314);
   DLX_INST_DATA_PATH_DECODE_RF_U1514 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4496, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2315);
   DLX_INST_DATA_PATH_DECODE_RF_U1513 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4495, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2316);
   DLX_INST_DATA_PATH_DECODE_RF_U1512 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4494, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2317);
   DLX_INST_DATA_PATH_DECODE_RF_U1511 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4493, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2318);
   DLX_INST_DATA_PATH_DECODE_RF_U1510 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4492, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2319);
   DLX_INST_DATA_PATH_DECODE_RF_U1509 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4491, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2320);
   DLX_INST_DATA_PATH_DECODE_RF_U1508 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4490, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2321);
   DLX_INST_DATA_PATH_DECODE_RF_U1507 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4489, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2322);
   DLX_INST_DATA_PATH_DECODE_RF_U1506 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4488, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2323);
   DLX_INST_DATA_PATH_DECODE_RF_U1505 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4487, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2324);
   DLX_INST_DATA_PATH_DECODE_RF_U1504 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4486, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2325);
   DLX_INST_DATA_PATH_DECODE_RF_U1503 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4485, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2326);
   DLX_INST_DATA_PATH_DECODE_RF_U1502 : NOR2_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_20_port, A2 => 
                           DLX_INST_IR_OUT_signal_19_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6518);
   DLX_INST_DATA_PATH_DECODE_RF_U1501 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_18_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6524);
   DLX_INST_DATA_PATH_DECODE_RF_U1500 : NOR3_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_16_port, A2 => 
                           DLX_INST_IR_OUT_signal_17_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6524, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6498);
   DLX_INST_DATA_PATH_DECODE_RF_U1499 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_19_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6526);
   DLX_INST_DATA_PATH_DECODE_RF_U1498 : NOR2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6526, A2 => 
                           DLX_INST_IR_OUT_signal_20_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6519);
   DLX_INST_DATA_PATH_DECODE_RF_U1497 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_17_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6523);
   DLX_INST_DATA_PATH_DECODE_RF_U1496 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_16_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6521);
   DLX_INST_DATA_PATH_DECODE_RF_U1495 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6524, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6523, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6521, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6506);
   DLX_INST_DATA_PATH_DECODE_RF_U1494 : AND2_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_20_port, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6526, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6509);
   DLX_INST_DATA_PATH_DECODE_RF_U1493 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6524, A2 => 
                           DLX_INST_IR_OUT_signal_17_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6521, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6504);
   DLX_INST_DATA_PATH_DECODE_RF_U1492 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4580, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4322, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6525);
   DLX_INST_DATA_PATH_DECODE_RF_U1491 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6767, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6863, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6525, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6513);
   DLX_INST_DATA_PATH_DECODE_RF_U1490 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6523, A2 => 
                           DLX_INST_IR_OUT_signal_18_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6521, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6508);
   DLX_INST_DATA_PATH_DECODE_RF_U1489 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6523, A2 => 
                           DLX_INST_IR_OUT_signal_16_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6524, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6502);
   DLX_INST_DATA_PATH_DECODE_RF_U1488 : NOR3_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_16_port, A2 => 
                           DLX_INST_IR_OUT_signal_18_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6523, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6507);
   DLX_INST_DATA_PATH_DECODE_RF_U1487 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4708, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4226, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4482, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6522);
   DLX_INST_DATA_PATH_DECODE_RF_U1486 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6735, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6831, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6522, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6514);
   DLX_INST_DATA_PATH_DECODE_RF_U1485 : NOR3_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_17_port, A2 => 
                           DLX_INST_IR_OUT_signal_18_port, A3 => 
                           DLX_INST_IR_OUT_signal_16_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6501);
   DLX_INST_DATA_PATH_DECODE_RF_U1484 : NOR3_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_17_port, A2 => 
                           DLX_INST_IR_OUT_signal_18_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6521, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6500);
   DLX_INST_DATA_PATH_DECODE_RF_U1483 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4516, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4258, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6520);
   DLX_INST_DATA_PATH_DECODE_RF_U1482 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6799, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6703, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6520, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6515);
   DLX_INST_DATA_PATH_DECODE_RF_U1481 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4740, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4194, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4450, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6517);
   DLX_INST_DATA_PATH_DECODE_RF_U1480 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6895, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6671, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6517, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6516);
   DLX_INST_DATA_PATH_DECODE_RF_U1479 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6513, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6514, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6515, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6516, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6511);
   DLX_INST_DATA_PATH_DECODE_RF_U1478 : AND3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, A2 => 
                           DLX_INST_IR_OUT_signal_20_port, A3 => 
                           DLX_INST_IR_OUT_signal_19_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6505);
   DLX_INST_DATA_PATH_DECODE_RF_U1477 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4644, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4386, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6512);
   DLX_INST_DATA_PATH_DECODE_RF_U1476 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6511, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_0_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6512, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6493);
   DLX_INST_DATA_PATH_DECODE_RF_U1475 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4612, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4354, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6510);
   DLX_INST_DATA_PATH_DECODE_RF_U1474 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7055, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7087, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6510, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6494);
   DLX_INST_DATA_PATH_DECODE_RF_U1473 : AND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6509, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6499);
   DLX_INST_DATA_PATH_DECODE_RF_U1472 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4676, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4418, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6503);
   DLX_INST_DATA_PATH_DECODE_RF_U1471 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6927, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6991, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6503, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6495);
   DLX_INST_DATA_PATH_DECODE_RF_U1470 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4548, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4290, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6497);
   DLX_INST_DATA_PATH_DECODE_RF_U1469 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7023, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6959, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6497, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6496);
   DLX_INST_DATA_PATH_DECODE_RF_U1468 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6493, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6494, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6495, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6496, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4099);
   DLX_INST_DATA_PATH_DECODE_RF_U1467 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4579, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4321, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6492);
   DLX_INST_DATA_PATH_DECODE_RF_U1466 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6766, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6862, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6492, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6485);
   DLX_INST_DATA_PATH_DECODE_RF_U1465 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4707, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4225, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4481, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6491);
   DLX_INST_DATA_PATH_DECODE_RF_U1464 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6734, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6830, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6491, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6486);
   DLX_INST_DATA_PATH_DECODE_RF_U1463 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4515, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4257, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6490);
   DLX_INST_DATA_PATH_DECODE_RF_U1462 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6798, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6702, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6490, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6487);
   DLX_INST_DATA_PATH_DECODE_RF_U1461 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4739, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4193, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4449, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6489);
   DLX_INST_DATA_PATH_DECODE_RF_U1460 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6894, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6670, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6489, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6488);
   DLX_INST_DATA_PATH_DECODE_RF_U1459 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6485, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6486, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6487, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6488, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6483);
   DLX_INST_DATA_PATH_DECODE_RF_U1458 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4643, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4385, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6484);
   DLX_INST_DATA_PATH_DECODE_RF_U1457 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6483, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_1_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6484, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6476);
   DLX_INST_DATA_PATH_DECODE_RF_U1456 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4611, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4353, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6482);
   DLX_INST_DATA_PATH_DECODE_RF_U1455 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7054, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7086, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6482, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6477);
   DLX_INST_DATA_PATH_DECODE_RF_U1454 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4675, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4417, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6481);
   DLX_INST_DATA_PATH_DECODE_RF_U1453 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6926, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6990, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6481, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6478);
   DLX_INST_DATA_PATH_DECODE_RF_U1452 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4547, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4289, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6480);
   DLX_INST_DATA_PATH_DECODE_RF_U1451 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7022, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6958, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6480, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6479);
   DLX_INST_DATA_PATH_DECODE_RF_U1450 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6476, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6477, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6478, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6479, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4100);
   DLX_INST_DATA_PATH_DECODE_RF_U1449 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4578, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4320, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6475);
   DLX_INST_DATA_PATH_DECODE_RF_U1448 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6765, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6861, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6475, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6468);
   DLX_INST_DATA_PATH_DECODE_RF_U1447 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4706, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4224, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4480, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6474);
   DLX_INST_DATA_PATH_DECODE_RF_U1446 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6733, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6829, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6474, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6469);
   DLX_INST_DATA_PATH_DECODE_RF_U1445 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4514, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4256, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6473);
   DLX_INST_DATA_PATH_DECODE_RF_U1444 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6797, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6701, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6473, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6470);
   DLX_INST_DATA_PATH_DECODE_RF_U1443 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4738, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4192, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4448, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6472);
   DLX_INST_DATA_PATH_DECODE_RF_U1442 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6893, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6669, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6472, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6471);
   DLX_INST_DATA_PATH_DECODE_RF_U1441 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6468, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6469, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6470, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6471, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6466);
   DLX_INST_DATA_PATH_DECODE_RF_U1440 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4642, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4384, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6467);
   DLX_INST_DATA_PATH_DECODE_RF_U1439 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6466, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_2_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6467, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6459);
   DLX_INST_DATA_PATH_DECODE_RF_U1438 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4610, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6465);
   DLX_INST_DATA_PATH_DECODE_RF_U1437 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7053, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7085, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6465, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6460);
   DLX_INST_DATA_PATH_DECODE_RF_U1436 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4674, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4416, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6464);
   DLX_INST_DATA_PATH_DECODE_RF_U1435 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6925, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6989, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6464, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6461);
   DLX_INST_DATA_PATH_DECODE_RF_U1434 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4546, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4288, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6463);
   DLX_INST_DATA_PATH_DECODE_RF_U1433 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7021, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6957, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6463, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6462);
   DLX_INST_DATA_PATH_DECODE_RF_U1432 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6459, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6460, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6461, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6462, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4101);
   DLX_INST_DATA_PATH_DECODE_RF_U1431 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4577, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4319, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6458);
   DLX_INST_DATA_PATH_DECODE_RF_U1430 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6764, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6860, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6458, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6451);
   DLX_INST_DATA_PATH_DECODE_RF_U1429 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4705, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4223, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4479, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6457);
   DLX_INST_DATA_PATH_DECODE_RF_U1428 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6732, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6828, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6457, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6452);
   DLX_INST_DATA_PATH_DECODE_RF_U1427 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4513, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4255, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6456);
   DLX_INST_DATA_PATH_DECODE_RF_U1426 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6796, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6700, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6456, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6453);
   DLX_INST_DATA_PATH_DECODE_RF_U1425 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4737, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4191, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4447, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6455);
   DLX_INST_DATA_PATH_DECODE_RF_U1424 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6892, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6668, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6455, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6454);
   DLX_INST_DATA_PATH_DECODE_RF_U1423 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6451, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6452, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6453, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6454, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6449);
   DLX_INST_DATA_PATH_DECODE_RF_U1422 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4641, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4383, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6450);
   DLX_INST_DATA_PATH_DECODE_RF_U1421 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6449, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_3_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6450, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6442);
   DLX_INST_DATA_PATH_DECODE_RF_U1420 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4609, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4351, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6448);
   DLX_INST_DATA_PATH_DECODE_RF_U1419 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7052, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7084, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6448, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6443);
   DLX_INST_DATA_PATH_DECODE_RF_U1418 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4673, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4415, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6447);
   DLX_INST_DATA_PATH_DECODE_RF_U1417 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6924, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6988, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6447, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6444);
   DLX_INST_DATA_PATH_DECODE_RF_U1416 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4545, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4287, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6446);
   DLX_INST_DATA_PATH_DECODE_RF_U1415 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7020, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6956, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6446, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6445);
   DLX_INST_DATA_PATH_DECODE_RF_U1414 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6442, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6443, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6444, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6445, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4102);
   DLX_INST_DATA_PATH_DECODE_RF_U1413 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4576, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4318, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6441);
   DLX_INST_DATA_PATH_DECODE_RF_U1412 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6763, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6859, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6441, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6434);
   DLX_INST_DATA_PATH_DECODE_RF_U1411 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4704, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4222, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4478, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6440);
   DLX_INST_DATA_PATH_DECODE_RF_U1410 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6731, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6827, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6440, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6435);
   DLX_INST_DATA_PATH_DECODE_RF_U1409 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4512, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4254, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6439);
   DLX_INST_DATA_PATH_DECODE_RF_U1408 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6795, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6699, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6439, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6436);
   DLX_INST_DATA_PATH_DECODE_RF_U1407 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4736, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4190, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4446, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6438);
   DLX_INST_DATA_PATH_DECODE_RF_U1406 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6891, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6667, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6438, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6437);
   DLX_INST_DATA_PATH_DECODE_RF_U1405 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6434, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6435, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6436, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6437, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6432);
   DLX_INST_DATA_PATH_DECODE_RF_U1404 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4640, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6433);
   DLX_INST_DATA_PATH_DECODE_RF_U1403 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6432, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_4_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6433, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6425);
   DLX_INST_DATA_PATH_DECODE_RF_U1402 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4608, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4350, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6431);
   DLX_INST_DATA_PATH_DECODE_RF_U1401 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7051, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7083, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6431, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6426);
   DLX_INST_DATA_PATH_DECODE_RF_U1400 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4672, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4414, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6430);
   DLX_INST_DATA_PATH_DECODE_RF_U1399 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6923, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6987, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6430, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6427);
   DLX_INST_DATA_PATH_DECODE_RF_U1398 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4544, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4286, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6429);
   DLX_INST_DATA_PATH_DECODE_RF_U1397 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7019, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6955, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6429, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6428);
   DLX_INST_DATA_PATH_DECODE_RF_U1396 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6425, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6426, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6427, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6428, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4103);
   DLX_INST_DATA_PATH_DECODE_RF_U1395 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4575, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4317, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6424);
   DLX_INST_DATA_PATH_DECODE_RF_U1394 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6762, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6858, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6424, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6417);
   DLX_INST_DATA_PATH_DECODE_RF_U1393 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4703, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4221, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4477, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6423);
   DLX_INST_DATA_PATH_DECODE_RF_U1392 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6730, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6826, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6423, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6418);
   DLX_INST_DATA_PATH_DECODE_RF_U1391 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4511, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4253, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6422);
   DLX_INST_DATA_PATH_DECODE_RF_U1390 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6794, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6698, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6422, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6419);
   DLX_INST_DATA_PATH_DECODE_RF_U1389 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4735, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4189, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4445, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6421);
   DLX_INST_DATA_PATH_DECODE_RF_U1388 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6890, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6666, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6421, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6420);
   DLX_INST_DATA_PATH_DECODE_RF_U1387 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6417, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6418, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6419, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6420, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6415);
   DLX_INST_DATA_PATH_DECODE_RF_U1386 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4639, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4381, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6416);
   DLX_INST_DATA_PATH_DECODE_RF_U1385 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6415, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_5_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6416, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6408);
   DLX_INST_DATA_PATH_DECODE_RF_U1384 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4607, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4349, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6414);
   DLX_INST_DATA_PATH_DECODE_RF_U1383 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7050, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7082, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6414, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6409);
   DLX_INST_DATA_PATH_DECODE_RF_U1382 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4671, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4413, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6413);
   DLX_INST_DATA_PATH_DECODE_RF_U1381 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6922, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6986, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6413, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6410);
   DLX_INST_DATA_PATH_DECODE_RF_U1380 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4543, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4285, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6412);
   DLX_INST_DATA_PATH_DECODE_RF_U1379 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7018, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6954, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6412, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6411);
   DLX_INST_DATA_PATH_DECODE_RF_U1378 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6408, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6409, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6410, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6411, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4104);
   DLX_INST_DATA_PATH_DECODE_RF_U1377 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4574, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4316, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6407);
   DLX_INST_DATA_PATH_DECODE_RF_U1376 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6761, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6857, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6407, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6400);
   DLX_INST_DATA_PATH_DECODE_RF_U1375 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4702, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4220, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4476, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6406);
   DLX_INST_DATA_PATH_DECODE_RF_U1374 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6729, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6825, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6406, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6401);
   DLX_INST_DATA_PATH_DECODE_RF_U1373 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4510, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4252, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6405);
   DLX_INST_DATA_PATH_DECODE_RF_U1372 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6793, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6697, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6405, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6402);
   DLX_INST_DATA_PATH_DECODE_RF_U1371 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4734, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4188, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4444, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6404);
   DLX_INST_DATA_PATH_DECODE_RF_U1370 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6889, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6665, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6404, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6403);
   DLX_INST_DATA_PATH_DECODE_RF_U1369 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6400, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6401, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6402, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6403, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6398);
   DLX_INST_DATA_PATH_DECODE_RF_U1368 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4638, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4380, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6399);
   DLX_INST_DATA_PATH_DECODE_RF_U1367 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6398, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_6_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6399, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6391);
   DLX_INST_DATA_PATH_DECODE_RF_U1366 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4606, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4348, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6397);
   DLX_INST_DATA_PATH_DECODE_RF_U1365 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7049, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7081, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6397, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6392);
   DLX_INST_DATA_PATH_DECODE_RF_U1364 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4670, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4412, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6396);
   DLX_INST_DATA_PATH_DECODE_RF_U1363 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6921, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6985, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6396, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6393);
   DLX_INST_DATA_PATH_DECODE_RF_U1362 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4284, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6395);
   DLX_INST_DATA_PATH_DECODE_RF_U1361 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7017, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6953, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6395, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6394);
   DLX_INST_DATA_PATH_DECODE_RF_U1360 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6391, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6392, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6393, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6394, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4105);
   DLX_INST_DATA_PATH_DECODE_RF_U1359 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4573, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4315, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6390);
   DLX_INST_DATA_PATH_DECODE_RF_U1358 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6760, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6856, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6390, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6383);
   DLX_INST_DATA_PATH_DECODE_RF_U1357 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4701, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4219, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4475, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6389);
   DLX_INST_DATA_PATH_DECODE_RF_U1356 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6728, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6824, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6389, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6384);
   DLX_INST_DATA_PATH_DECODE_RF_U1355 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4509, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4251, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6388);
   DLX_INST_DATA_PATH_DECODE_RF_U1354 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6792, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6696, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6388, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6385);
   DLX_INST_DATA_PATH_DECODE_RF_U1353 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4733, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4187, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4443, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6387);
   DLX_INST_DATA_PATH_DECODE_RF_U1352 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6888, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6664, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6387, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6386);
   DLX_INST_DATA_PATH_DECODE_RF_U1351 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6383, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6384, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6385, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6386, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6381);
   DLX_INST_DATA_PATH_DECODE_RF_U1350 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4637, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4379, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6382);
   DLX_INST_DATA_PATH_DECODE_RF_U1349 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6381, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_7_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6382, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6374);
   DLX_INST_DATA_PATH_DECODE_RF_U1348 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4605, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6380);
   DLX_INST_DATA_PATH_DECODE_RF_U1347 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7048, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7080, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6380, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6375);
   DLX_INST_DATA_PATH_DECODE_RF_U1346 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4669, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4411, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6379);
   DLX_INST_DATA_PATH_DECODE_RF_U1345 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6920, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6984, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6379, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6376);
   DLX_INST_DATA_PATH_DECODE_RF_U1344 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4541, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4283, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6378);
   DLX_INST_DATA_PATH_DECODE_RF_U1343 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7016, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6952, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6378, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6377);
   DLX_INST_DATA_PATH_DECODE_RF_U1342 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6374, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6375, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6376, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6377, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4106);
   DLX_INST_DATA_PATH_DECODE_RF_U1341 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4572, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4314, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6373);
   DLX_INST_DATA_PATH_DECODE_RF_U1340 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6759, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6855, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6373, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6366);
   DLX_INST_DATA_PATH_DECODE_RF_U1339 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4700, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4218, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4474, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6372);
   DLX_INST_DATA_PATH_DECODE_RF_U1338 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6727, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6823, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6372, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6367);
   DLX_INST_DATA_PATH_DECODE_RF_U1337 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4508, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4250, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6371);
   DLX_INST_DATA_PATH_DECODE_RF_U1336 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6791, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6695, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6371, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6368);
   DLX_INST_DATA_PATH_DECODE_RF_U1335 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4732, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4186, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4442, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6370);
   DLX_INST_DATA_PATH_DECODE_RF_U1334 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6887, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6663, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6370, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6369);
   DLX_INST_DATA_PATH_DECODE_RF_U1333 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6366, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6367, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6368, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6369, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6364);
   DLX_INST_DATA_PATH_DECODE_RF_U1332 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4636, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4378, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6365);
   DLX_INST_DATA_PATH_DECODE_RF_U1331 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6364, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_8_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6365, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6357);
   DLX_INST_DATA_PATH_DECODE_RF_U1330 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4604, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4346, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6363);
   DLX_INST_DATA_PATH_DECODE_RF_U1329 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7047, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7079, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6363, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6358);
   DLX_INST_DATA_PATH_DECODE_RF_U1328 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4668, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4410, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6362);
   DLX_INST_DATA_PATH_DECODE_RF_U1327 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6919, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6983, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6362, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6359);
   DLX_INST_DATA_PATH_DECODE_RF_U1326 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4540, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4282, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6361);
   DLX_INST_DATA_PATH_DECODE_RF_U1325 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7015, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6951, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6361, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6360);
   DLX_INST_DATA_PATH_DECODE_RF_U1324 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6357, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6358, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6359, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6360, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4107);
   DLX_INST_DATA_PATH_DECODE_RF_U1323 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4571, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4313, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6356);
   DLX_INST_DATA_PATH_DECODE_RF_U1322 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6758, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6854, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6356, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6349);
   DLX_INST_DATA_PATH_DECODE_RF_U1321 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4699, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4217, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4473, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6355);
   DLX_INST_DATA_PATH_DECODE_RF_U1320 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6726, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6822, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6355, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6350);
   DLX_INST_DATA_PATH_DECODE_RF_U1319 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4507, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4249, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6354);
   DLX_INST_DATA_PATH_DECODE_RF_U1318 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6790, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6694, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6354, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6351);
   DLX_INST_DATA_PATH_DECODE_RF_U1317 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4731, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4185, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4441, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6353);
   DLX_INST_DATA_PATH_DECODE_RF_U1316 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6886, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6662, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6353, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6352);
   DLX_INST_DATA_PATH_DECODE_RF_U1315 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6349, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6350, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6351, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6352, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6347);
   DLX_INST_DATA_PATH_DECODE_RF_U1314 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4635, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6348);
   DLX_INST_DATA_PATH_DECODE_RF_U1313 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6347, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_9_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6348, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6340);
   DLX_INST_DATA_PATH_DECODE_RF_U1312 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4603, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4345, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6346);
   DLX_INST_DATA_PATH_DECODE_RF_U1311 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7046, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7078, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6346, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6341);
   DLX_INST_DATA_PATH_DECODE_RF_U1310 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4667, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4409, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6345);
   DLX_INST_DATA_PATH_DECODE_RF_U1309 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6918, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6982, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6345, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6342);
   DLX_INST_DATA_PATH_DECODE_RF_U1308 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4539, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4281, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6344);
   DLX_INST_DATA_PATH_DECODE_RF_U1307 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7014, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6950, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6344, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6343);
   DLX_INST_DATA_PATH_DECODE_RF_U1306 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6340, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6341, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6342, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6343, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4108);
   DLX_INST_DATA_PATH_DECODE_RF_U1305 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4570, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4312, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6339);
   DLX_INST_DATA_PATH_DECODE_RF_U1304 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6757, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6853, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6339, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6332);
   DLX_INST_DATA_PATH_DECODE_RF_U1303 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4698, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4216, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4472, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6338);
   DLX_INST_DATA_PATH_DECODE_RF_U1302 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6725, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6821, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6338, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6333);
   DLX_INST_DATA_PATH_DECODE_RF_U1301 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4506, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4248, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6337);
   DLX_INST_DATA_PATH_DECODE_RF_U1300 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6789, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6693, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6337, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6334);
   DLX_INST_DATA_PATH_DECODE_RF_U1299 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4730, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4184, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4440, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6336);
   DLX_INST_DATA_PATH_DECODE_RF_U1298 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6885, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6661, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6336, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6335);
   DLX_INST_DATA_PATH_DECODE_RF_U1297 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6332, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6333, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6334, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6335, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6330);
   DLX_INST_DATA_PATH_DECODE_RF_U1296 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4634, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4376, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6331);
   DLX_INST_DATA_PATH_DECODE_RF_U1295 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6330, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_10_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6331, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6323);
   DLX_INST_DATA_PATH_DECODE_RF_U1294 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4602, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4344, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6329);
   DLX_INST_DATA_PATH_DECODE_RF_U1293 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7045, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7077, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6329, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6324);
   DLX_INST_DATA_PATH_DECODE_RF_U1292 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4666, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4408, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6328);
   DLX_INST_DATA_PATH_DECODE_RF_U1291 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6917, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6981, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6328, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6325);
   DLX_INST_DATA_PATH_DECODE_RF_U1290 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4538, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4280, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6327);
   DLX_INST_DATA_PATH_DECODE_RF_U1289 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7013, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6949, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6327, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6326);
   DLX_INST_DATA_PATH_DECODE_RF_U1288 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6323, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6324, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6325, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6326, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4109);
   DLX_INST_DATA_PATH_DECODE_RF_U1287 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4569, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4311, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6322);
   DLX_INST_DATA_PATH_DECODE_RF_U1286 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6756, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6852, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6322, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6315);
   DLX_INST_DATA_PATH_DECODE_RF_U1285 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4697, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4215, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4471, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6321);
   DLX_INST_DATA_PATH_DECODE_RF_U1284 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6724, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6820, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6321, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6316);
   DLX_INST_DATA_PATH_DECODE_RF_U1283 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4505, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4247, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6320);
   DLX_INST_DATA_PATH_DECODE_RF_U1282 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6788, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6692, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6320, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6317);
   DLX_INST_DATA_PATH_DECODE_RF_U1281 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4729, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4183, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4439, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6319);
   DLX_INST_DATA_PATH_DECODE_RF_U1280 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6884, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6660, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6319, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6318);
   DLX_INST_DATA_PATH_DECODE_RF_U1279 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6315, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6316, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6317, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6318, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6313);
   DLX_INST_DATA_PATH_DECODE_RF_U1278 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4633, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4375, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6314);
   DLX_INST_DATA_PATH_DECODE_RF_U1277 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6313, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_11_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6314, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6306);
   DLX_INST_DATA_PATH_DECODE_RF_U1276 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4601, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4343, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6312);
   DLX_INST_DATA_PATH_DECODE_RF_U1275 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7044, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7076, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6312, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6307);
   DLX_INST_DATA_PATH_DECODE_RF_U1274 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4665, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4407, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6311);
   DLX_INST_DATA_PATH_DECODE_RF_U1273 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6916, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6980, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6311, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6308);
   DLX_INST_DATA_PATH_DECODE_RF_U1272 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4537, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4279, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6310);
   DLX_INST_DATA_PATH_DECODE_RF_U1271 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7012, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6948, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6310, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6309);
   DLX_INST_DATA_PATH_DECODE_RF_U1270 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6306, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6307, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6308, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6309, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4110);
   DLX_INST_DATA_PATH_DECODE_RF_U1269 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4568, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4310, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6305);
   DLX_INST_DATA_PATH_DECODE_RF_U1268 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6755, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6851, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6305, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6298);
   DLX_INST_DATA_PATH_DECODE_RF_U1267 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4696, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4214, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4470, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6304);
   DLX_INST_DATA_PATH_DECODE_RF_U1266 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6723, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6819, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6304, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6299);
   DLX_INST_DATA_PATH_DECODE_RF_U1265 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4504, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4246, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6303);
   DLX_INST_DATA_PATH_DECODE_RF_U1264 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6787, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6691, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6303, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6300);
   DLX_INST_DATA_PATH_DECODE_RF_U1263 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4728, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4182, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4438, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6302);
   DLX_INST_DATA_PATH_DECODE_RF_U1262 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6883, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6659, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6302, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6301);
   DLX_INST_DATA_PATH_DECODE_RF_U1261 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6298, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6299, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6300, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6301, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6296);
   DLX_INST_DATA_PATH_DECODE_RF_U1260 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4632, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4374, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6297);
   DLX_INST_DATA_PATH_DECODE_RF_U1259 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6296, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_12_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6297, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6289);
   DLX_INST_DATA_PATH_DECODE_RF_U1258 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4600, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4342, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6295);
   DLX_INST_DATA_PATH_DECODE_RF_U1257 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7043, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7075, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6295, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6290);
   DLX_INST_DATA_PATH_DECODE_RF_U1256 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4664, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4406, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6294);
   DLX_INST_DATA_PATH_DECODE_RF_U1255 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6915, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6979, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6294, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6291);
   DLX_INST_DATA_PATH_DECODE_RF_U1254 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4536, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4278, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6293);
   DLX_INST_DATA_PATH_DECODE_RF_U1253 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7011, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6947, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6293, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6292);
   DLX_INST_DATA_PATH_DECODE_RF_U1252 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6289, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6290, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6291, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6292, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4111);
   DLX_INST_DATA_PATH_DECODE_RF_U1251 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4567, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4309, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6288);
   DLX_INST_DATA_PATH_DECODE_RF_U1250 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6754, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6850, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6288, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6281);
   DLX_INST_DATA_PATH_DECODE_RF_U1249 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4695, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4213, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4469, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6287);
   DLX_INST_DATA_PATH_DECODE_RF_U1248 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6722, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6818, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6287, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6282);
   DLX_INST_DATA_PATH_DECODE_RF_U1247 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4503, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4245, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6286);
   DLX_INST_DATA_PATH_DECODE_RF_U1246 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6786, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6690, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6286, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6283);
   DLX_INST_DATA_PATH_DECODE_RF_U1245 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4727, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4181, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4437, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6285);
   DLX_INST_DATA_PATH_DECODE_RF_U1244 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6882, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6658, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6285, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6284);
   DLX_INST_DATA_PATH_DECODE_RF_U1243 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6281, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6282, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6283, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6284, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6279);
   DLX_INST_DATA_PATH_DECODE_RF_U1242 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4631, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4373, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6280);
   DLX_INST_DATA_PATH_DECODE_RF_U1241 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6279, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_13_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6280, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6272);
   DLX_INST_DATA_PATH_DECODE_RF_U1240 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4599, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4341, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6278);
   DLX_INST_DATA_PATH_DECODE_RF_U1239 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7042, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7074, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6278, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6273);
   DLX_INST_DATA_PATH_DECODE_RF_U1238 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4663, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4405, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6277);
   DLX_INST_DATA_PATH_DECODE_RF_U1237 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6914, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6978, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6277, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6274);
   DLX_INST_DATA_PATH_DECODE_RF_U1236 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4535, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4277, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6276);
   DLX_INST_DATA_PATH_DECODE_RF_U1235 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7010, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6946, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6276, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6275);
   DLX_INST_DATA_PATH_DECODE_RF_U1234 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6272, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6273, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6274, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6275, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4112);
   DLX_INST_DATA_PATH_DECODE_RF_U1233 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4566, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4308, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6271);
   DLX_INST_DATA_PATH_DECODE_RF_U1232 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6753, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6849, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6271, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6264);
   DLX_INST_DATA_PATH_DECODE_RF_U1231 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4694, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4212, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4468, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6270);
   DLX_INST_DATA_PATH_DECODE_RF_U1230 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6721, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6817, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6270, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6265);
   DLX_INST_DATA_PATH_DECODE_RF_U1229 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4502, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4244, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6269);
   DLX_INST_DATA_PATH_DECODE_RF_U1228 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6785, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6689, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6269, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6266);
   DLX_INST_DATA_PATH_DECODE_RF_U1227 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4726, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4180, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4436, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6268);
   DLX_INST_DATA_PATH_DECODE_RF_U1226 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6881, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6657, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6268, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6267);
   DLX_INST_DATA_PATH_DECODE_RF_U1225 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6264, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6265, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6266, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6267, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6262);
   DLX_INST_DATA_PATH_DECODE_RF_U1224 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4630, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4372, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6263);
   DLX_INST_DATA_PATH_DECODE_RF_U1223 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6262, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_14_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6263, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6255);
   DLX_INST_DATA_PATH_DECODE_RF_U1222 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4598, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4340, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6261);
   DLX_INST_DATA_PATH_DECODE_RF_U1221 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7041, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7073, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6261, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6256);
   DLX_INST_DATA_PATH_DECODE_RF_U1220 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4662, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4404, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6260);
   DLX_INST_DATA_PATH_DECODE_RF_U1219 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6913, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6977, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6260, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6257);
   DLX_INST_DATA_PATH_DECODE_RF_U1218 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4276, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6259);
   DLX_INST_DATA_PATH_DECODE_RF_U1217 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7009, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6945, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6259, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6258);
   DLX_INST_DATA_PATH_DECODE_RF_U1216 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6255, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6256, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6257, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6258, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4113);
   DLX_INST_DATA_PATH_DECODE_RF_U1215 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4565, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4307, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6254);
   DLX_INST_DATA_PATH_DECODE_RF_U1214 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6752, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6848, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6254, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6247);
   DLX_INST_DATA_PATH_DECODE_RF_U1213 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4693, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4211, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4467, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6253);
   DLX_INST_DATA_PATH_DECODE_RF_U1212 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6720, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6816, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6253, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6248);
   DLX_INST_DATA_PATH_DECODE_RF_U1211 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4501, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4243, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6252);
   DLX_INST_DATA_PATH_DECODE_RF_U1210 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6784, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6688, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6252, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6249);
   DLX_INST_DATA_PATH_DECODE_RF_U1209 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4725, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4179, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4435, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6251);
   DLX_INST_DATA_PATH_DECODE_RF_U1208 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6880, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6656, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6251, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6250);
   DLX_INST_DATA_PATH_DECODE_RF_U1207 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6247, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6248, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6249, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6250, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6245);
   DLX_INST_DATA_PATH_DECODE_RF_U1206 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4629, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6246);
   DLX_INST_DATA_PATH_DECODE_RF_U1205 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6245, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_15_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6246, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6238);
   DLX_INST_DATA_PATH_DECODE_RF_U1204 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4597, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4339, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6244);
   DLX_INST_DATA_PATH_DECODE_RF_U1203 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7040, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7072, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6244, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6239);
   DLX_INST_DATA_PATH_DECODE_RF_U1202 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4661, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4403, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6243);
   DLX_INST_DATA_PATH_DECODE_RF_U1201 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6912, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6976, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6243, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6240);
   DLX_INST_DATA_PATH_DECODE_RF_U1200 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4533, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4275, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6242);
   DLX_INST_DATA_PATH_DECODE_RF_U1199 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7008, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6944, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6242, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6241);
   DLX_INST_DATA_PATH_DECODE_RF_U1198 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6238, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6239, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6240, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6241, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4114);
   DLX_INST_DATA_PATH_DECODE_RF_U1197 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4564, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4306, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6237);
   DLX_INST_DATA_PATH_DECODE_RF_U1196 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6751, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6847, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6237, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6230);
   DLX_INST_DATA_PATH_DECODE_RF_U1195 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4692, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4210, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4466, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6236);
   DLX_INST_DATA_PATH_DECODE_RF_U1194 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6719, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6815, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6236, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6231);
   DLX_INST_DATA_PATH_DECODE_RF_U1193 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4500, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4242, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6235);
   DLX_INST_DATA_PATH_DECODE_RF_U1192 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6783, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6687, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6235, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6232);
   DLX_INST_DATA_PATH_DECODE_RF_U1191 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4724, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4178, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4434, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6234);
   DLX_INST_DATA_PATH_DECODE_RF_U1190 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6879, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6655, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6234, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6233);
   DLX_INST_DATA_PATH_DECODE_RF_U1189 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6230, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6231, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6232, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6233, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6228);
   DLX_INST_DATA_PATH_DECODE_RF_U1188 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4628, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4370, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6229);
   DLX_INST_DATA_PATH_DECODE_RF_U1187 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6228, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_16_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6229, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6221);
   DLX_INST_DATA_PATH_DECODE_RF_U1186 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4596, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4338, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6227);
   DLX_INST_DATA_PATH_DECODE_RF_U1185 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7039, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7071, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6227, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6222);
   DLX_INST_DATA_PATH_DECODE_RF_U1184 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4660, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4402, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6226);
   DLX_INST_DATA_PATH_DECODE_RF_U1183 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6911, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6975, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6226, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6223);
   DLX_INST_DATA_PATH_DECODE_RF_U1182 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4532, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4274, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6225);
   DLX_INST_DATA_PATH_DECODE_RF_U1181 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7007, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6943, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6225, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6224);
   DLX_INST_DATA_PATH_DECODE_RF_U1180 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6221, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6222, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6223, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6224, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4115);
   DLX_INST_DATA_PATH_DECODE_RF_U1179 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4563, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4305, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6220);
   DLX_INST_DATA_PATH_DECODE_RF_U1178 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6750, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6846, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6220, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6213);
   DLX_INST_DATA_PATH_DECODE_RF_U1177 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4691, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4209, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4465, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6219);
   DLX_INST_DATA_PATH_DECODE_RF_U1176 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6718, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6814, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6219, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6214);
   DLX_INST_DATA_PATH_DECODE_RF_U1175 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4499, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4241, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6218);
   DLX_INST_DATA_PATH_DECODE_RF_U1174 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6782, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6686, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6218, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6215);
   DLX_INST_DATA_PATH_DECODE_RF_U1173 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4723, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4177, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4433, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6217);
   DLX_INST_DATA_PATH_DECODE_RF_U1172 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6878, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6654, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6217, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6216);
   DLX_INST_DATA_PATH_DECODE_RF_U1171 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6213, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6214, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6215, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6216, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6211);
   DLX_INST_DATA_PATH_DECODE_RF_U1170 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4627, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4369, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6212);
   DLX_INST_DATA_PATH_DECODE_RF_U1169 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6211, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_17_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6212, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6204);
   DLX_INST_DATA_PATH_DECODE_RF_U1168 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4595, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4337, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6210);
   DLX_INST_DATA_PATH_DECODE_RF_U1167 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7038, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7070, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6210, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6205);
   DLX_INST_DATA_PATH_DECODE_RF_U1166 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4659, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4401, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6209);
   DLX_INST_DATA_PATH_DECODE_RF_U1165 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6910, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6974, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6209, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6206);
   DLX_INST_DATA_PATH_DECODE_RF_U1164 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4531, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4273, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6208);
   DLX_INST_DATA_PATH_DECODE_RF_U1163 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7006, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6942, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6208, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6207);
   DLX_INST_DATA_PATH_DECODE_RF_U1162 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6204, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6205, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6206, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6207, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4116);
   DLX_INST_DATA_PATH_DECODE_RF_U1161 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4562, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4304, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6203);
   DLX_INST_DATA_PATH_DECODE_RF_U1160 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6749, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6845, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6203, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6196);
   DLX_INST_DATA_PATH_DECODE_RF_U1159 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4690, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4208, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4464, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6202);
   DLX_INST_DATA_PATH_DECODE_RF_U1158 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6717, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6813, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6202, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6197);
   DLX_INST_DATA_PATH_DECODE_RF_U1157 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4498, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4240, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6201);
   DLX_INST_DATA_PATH_DECODE_RF_U1156 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6781, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6685, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6201, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6198);
   DLX_INST_DATA_PATH_DECODE_RF_U1155 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4722, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4176, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4432, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6200);
   DLX_INST_DATA_PATH_DECODE_RF_U1154 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6877, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6653, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6200, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6199);
   DLX_INST_DATA_PATH_DECODE_RF_U1153 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6196, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6197, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6198, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6199, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6194);
   DLX_INST_DATA_PATH_DECODE_RF_U1152 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4626, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4368, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6195);
   DLX_INST_DATA_PATH_DECODE_RF_U1151 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6194, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_18_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6195, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6187);
   DLX_INST_DATA_PATH_DECODE_RF_U1150 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4594, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4336, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6193);
   DLX_INST_DATA_PATH_DECODE_RF_U1149 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7037, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7069, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6193, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6188);
   DLX_INST_DATA_PATH_DECODE_RF_U1148 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4658, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4400, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6192);
   DLX_INST_DATA_PATH_DECODE_RF_U1147 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6909, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6973, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6192, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6189);
   DLX_INST_DATA_PATH_DECODE_RF_U1146 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4530, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4272, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6191);
   DLX_INST_DATA_PATH_DECODE_RF_U1145 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7005, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6941, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6191, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6190);
   DLX_INST_DATA_PATH_DECODE_RF_U1144 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6187, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6188, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6189, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6190, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4117);
   DLX_INST_DATA_PATH_DECODE_RF_U1143 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4561, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4303, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6186);
   DLX_INST_DATA_PATH_DECODE_RF_U1142 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6748, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6844, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6186, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6179);
   DLX_INST_DATA_PATH_DECODE_RF_U1141 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4689, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4207, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4463, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6185);
   DLX_INST_DATA_PATH_DECODE_RF_U1140 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6716, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6812, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6185, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6180);
   DLX_INST_DATA_PATH_DECODE_RF_U1139 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4497, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4239, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6184);
   DLX_INST_DATA_PATH_DECODE_RF_U1138 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6780, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6684, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6184, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6181);
   DLX_INST_DATA_PATH_DECODE_RF_U1137 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4721, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4175, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4431, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6183);
   DLX_INST_DATA_PATH_DECODE_RF_U1136 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6876, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6652, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6183, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6182);
   DLX_INST_DATA_PATH_DECODE_RF_U1135 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6179, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6180, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6181, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6182, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6177);
   DLX_INST_DATA_PATH_DECODE_RF_U1134 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4625, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4367, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6178);
   DLX_INST_DATA_PATH_DECODE_RF_U1133 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6177, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_19_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6178, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6170);
   DLX_INST_DATA_PATH_DECODE_RF_U1132 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4593, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4335, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6176);
   DLX_INST_DATA_PATH_DECODE_RF_U1131 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7036, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7068, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6176, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6171);
   DLX_INST_DATA_PATH_DECODE_RF_U1130 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4657, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4399, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6175);
   DLX_INST_DATA_PATH_DECODE_RF_U1129 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6908, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6972, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6175, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6172);
   DLX_INST_DATA_PATH_DECODE_RF_U1128 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4529, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4271, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6174);
   DLX_INST_DATA_PATH_DECODE_RF_U1127 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7004, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6940, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6174, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6173);
   DLX_INST_DATA_PATH_DECODE_RF_U1126 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6170, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6171, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6172, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6173, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4118);
   DLX_INST_DATA_PATH_DECODE_RF_U1125 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4560, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4302, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6169);
   DLX_INST_DATA_PATH_DECODE_RF_U1124 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6747, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6843, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6169, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6162);
   DLX_INST_DATA_PATH_DECODE_RF_U1123 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4688, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4206, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4462, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6168);
   DLX_INST_DATA_PATH_DECODE_RF_U1122 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6715, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6811, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6168, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6163);
   DLX_INST_DATA_PATH_DECODE_RF_U1121 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4496, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4238, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6167);
   DLX_INST_DATA_PATH_DECODE_RF_U1120 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6779, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6683, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6167, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6164);
   DLX_INST_DATA_PATH_DECODE_RF_U1119 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4720, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4174, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4430, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6166);
   DLX_INST_DATA_PATH_DECODE_RF_U1118 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6875, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6651, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6166, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6165);
   DLX_INST_DATA_PATH_DECODE_RF_U1117 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6162, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6163, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6164, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6165, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6160);
   DLX_INST_DATA_PATH_DECODE_RF_U1116 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4624, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4366, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6161);
   DLX_INST_DATA_PATH_DECODE_RF_U1115 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6160, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_20_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6161, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6153);
   DLX_INST_DATA_PATH_DECODE_RF_U1114 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4592, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4334, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6159);
   DLX_INST_DATA_PATH_DECODE_RF_U1113 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7035, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7067, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6159, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6154);
   DLX_INST_DATA_PATH_DECODE_RF_U1112 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4656, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4398, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6158);
   DLX_INST_DATA_PATH_DECODE_RF_U1111 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6907, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6971, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6158, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6155);
   DLX_INST_DATA_PATH_DECODE_RF_U1110 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4528, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4270, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6157);
   DLX_INST_DATA_PATH_DECODE_RF_U1109 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7003, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6939, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6157, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6156);
   DLX_INST_DATA_PATH_DECODE_RF_U1108 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6153, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6154, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6155, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6156, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4119);
   DLX_INST_DATA_PATH_DECODE_RF_U1107 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4301, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6152);
   DLX_INST_DATA_PATH_DECODE_RF_U1106 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6746, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6842, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6152, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6145);
   DLX_INST_DATA_PATH_DECODE_RF_U1105 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4687, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4205, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4461, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6151);
   DLX_INST_DATA_PATH_DECODE_RF_U1104 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6714, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6810, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6151, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6146);
   DLX_INST_DATA_PATH_DECODE_RF_U1103 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4495, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4237, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6150);
   DLX_INST_DATA_PATH_DECODE_RF_U1102 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6778, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6682, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6150, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6147);
   DLX_INST_DATA_PATH_DECODE_RF_U1101 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4719, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4173, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4429, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6149);
   DLX_INST_DATA_PATH_DECODE_RF_U1100 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6874, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6650, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6149, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6148);
   DLX_INST_DATA_PATH_DECODE_RF_U1099 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6145, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6146, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6147, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6148, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6143);
   DLX_INST_DATA_PATH_DECODE_RF_U1098 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4623, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4365, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6144);
   DLX_INST_DATA_PATH_DECODE_RF_U1097 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6143, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_21_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6144, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6136);
   DLX_INST_DATA_PATH_DECODE_RF_U1096 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4591, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4333, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6142);
   DLX_INST_DATA_PATH_DECODE_RF_U1095 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7034, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7066, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6142, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6137);
   DLX_INST_DATA_PATH_DECODE_RF_U1094 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4655, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4397, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6141);
   DLX_INST_DATA_PATH_DECODE_RF_U1093 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6906, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6970, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6141, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6138);
   DLX_INST_DATA_PATH_DECODE_RF_U1092 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4527, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4269, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6140);
   DLX_INST_DATA_PATH_DECODE_RF_U1091 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7002, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6938, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6140, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6139);
   DLX_INST_DATA_PATH_DECODE_RF_U1090 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6136, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6137, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6138, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6139, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4120);
   DLX_INST_DATA_PATH_DECODE_RF_U1089 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4558, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4300, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6135);
   DLX_INST_DATA_PATH_DECODE_RF_U1088 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6745, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6841, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6135, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6128);
   DLX_INST_DATA_PATH_DECODE_RF_U1087 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4686, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4204, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4460, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6134);
   DLX_INST_DATA_PATH_DECODE_RF_U1086 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6713, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6809, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6134, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6129);
   DLX_INST_DATA_PATH_DECODE_RF_U1085 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4494, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4236, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6133);
   DLX_INST_DATA_PATH_DECODE_RF_U1084 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6777, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6681, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6133, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6130);
   DLX_INST_DATA_PATH_DECODE_RF_U1083 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4718, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4172, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4428, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6132);
   DLX_INST_DATA_PATH_DECODE_RF_U1082 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6873, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6649, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6132, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6131);
   DLX_INST_DATA_PATH_DECODE_RF_U1081 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6128, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6129, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6130, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6131, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6126);
   DLX_INST_DATA_PATH_DECODE_RF_U1080 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4622, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4364, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6127);
   DLX_INST_DATA_PATH_DECODE_RF_U1079 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6126, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_22_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6127, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6119);
   DLX_INST_DATA_PATH_DECODE_RF_U1078 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4590, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4332, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6125);
   DLX_INST_DATA_PATH_DECODE_RF_U1077 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7033, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7065, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6125, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6120);
   DLX_INST_DATA_PATH_DECODE_RF_U1076 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4654, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4396, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6124);
   DLX_INST_DATA_PATH_DECODE_RF_U1075 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6905, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6969, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6124, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6121);
   DLX_INST_DATA_PATH_DECODE_RF_U1074 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4526, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4268, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6123);
   DLX_INST_DATA_PATH_DECODE_RF_U1073 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7001, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6937, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6123, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6122);
   DLX_INST_DATA_PATH_DECODE_RF_U1072 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6119, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6120, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6121, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6122, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4121);
   DLX_INST_DATA_PATH_DECODE_RF_U1071 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4557, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4299, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6118);
   DLX_INST_DATA_PATH_DECODE_RF_U1070 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6744, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6840, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6118, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6111);
   DLX_INST_DATA_PATH_DECODE_RF_U1069 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4685, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4203, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4459, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6117);
   DLX_INST_DATA_PATH_DECODE_RF_U1068 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6712, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6808, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6117, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6112);
   DLX_INST_DATA_PATH_DECODE_RF_U1067 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4493, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4235, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6116);
   DLX_INST_DATA_PATH_DECODE_RF_U1066 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6776, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6680, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6116, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6113);
   DLX_INST_DATA_PATH_DECODE_RF_U1065 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4717, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4171, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4427, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6115);
   DLX_INST_DATA_PATH_DECODE_RF_U1064 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6872, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6648, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6115, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6114);
   DLX_INST_DATA_PATH_DECODE_RF_U1063 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6111, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6112, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6113, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6114, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6109);
   DLX_INST_DATA_PATH_DECODE_RF_U1062 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4621, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4363, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6110);
   DLX_INST_DATA_PATH_DECODE_RF_U1061 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6109, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_23_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6110, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6102);
   DLX_INST_DATA_PATH_DECODE_RF_U1060 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4589, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4331, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6108);
   DLX_INST_DATA_PATH_DECODE_RF_U1059 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7032, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7064, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6108, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6103);
   DLX_INST_DATA_PATH_DECODE_RF_U1058 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4653, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4395, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6107);
   DLX_INST_DATA_PATH_DECODE_RF_U1057 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6904, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6968, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6107, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6104);
   DLX_INST_DATA_PATH_DECODE_RF_U1056 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4525, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4267, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6106);
   DLX_INST_DATA_PATH_DECODE_RF_U1055 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7000, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6936, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6106, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6105);
   DLX_INST_DATA_PATH_DECODE_RF_U1054 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6102, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6103, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6104, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6105, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4122);
   DLX_INST_DATA_PATH_DECODE_RF_U1053 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4556, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4298, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6101);
   DLX_INST_DATA_PATH_DECODE_RF_U1052 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6743, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6839, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6101, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6094);
   DLX_INST_DATA_PATH_DECODE_RF_U1051 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4684, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4202, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4458, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6100);
   DLX_INST_DATA_PATH_DECODE_RF_U1050 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6711, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6807, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6100, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6095);
   DLX_INST_DATA_PATH_DECODE_RF_U1049 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4492, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4234, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6099);
   DLX_INST_DATA_PATH_DECODE_RF_U1048 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6775, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6679, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6099, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6096);
   DLX_INST_DATA_PATH_DECODE_RF_U1047 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4716, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4170, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4426, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6098);
   DLX_INST_DATA_PATH_DECODE_RF_U1046 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6871, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6647, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6098, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6097);
   DLX_INST_DATA_PATH_DECODE_RF_U1045 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6094, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6095, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6096, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6097, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6092);
   DLX_INST_DATA_PATH_DECODE_RF_U1044 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4620, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6093);
   DLX_INST_DATA_PATH_DECODE_RF_U1043 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6092, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_24_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6093, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6085);
   DLX_INST_DATA_PATH_DECODE_RF_U1042 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4588, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4330, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6091);
   DLX_INST_DATA_PATH_DECODE_RF_U1041 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7031, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7063, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6091, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6086);
   DLX_INST_DATA_PATH_DECODE_RF_U1040 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4652, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4394, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6090);
   DLX_INST_DATA_PATH_DECODE_RF_U1039 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6903, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6967, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6090, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6087);
   DLX_INST_DATA_PATH_DECODE_RF_U1038 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4524, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4266, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6089);
   DLX_INST_DATA_PATH_DECODE_RF_U1037 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6999, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6935, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6089, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6088);
   DLX_INST_DATA_PATH_DECODE_RF_U1036 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6085, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6086, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6087, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6088, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4123);
   DLX_INST_DATA_PATH_DECODE_RF_U1035 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4555, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4297, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6084);
   DLX_INST_DATA_PATH_DECODE_RF_U1034 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6742, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6838, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6084, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6077);
   DLX_INST_DATA_PATH_DECODE_RF_U1033 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4683, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4201, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4457, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6083);
   DLX_INST_DATA_PATH_DECODE_RF_U1032 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6710, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6806, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6083, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6078);
   DLX_INST_DATA_PATH_DECODE_RF_U1031 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4491, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4233, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6082);
   DLX_INST_DATA_PATH_DECODE_RF_U1030 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6774, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6678, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6082, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6079);
   DLX_INST_DATA_PATH_DECODE_RF_U1029 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4715, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4169, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4425, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6081);
   DLX_INST_DATA_PATH_DECODE_RF_U1028 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6870, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6646, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6081, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6080);
   DLX_INST_DATA_PATH_DECODE_RF_U1027 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6077, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6078, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6079, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6080, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6075);
   DLX_INST_DATA_PATH_DECODE_RF_U1026 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4619, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4361, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6076);
   DLX_INST_DATA_PATH_DECODE_RF_U1025 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6075, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_25_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6076, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6068);
   DLX_INST_DATA_PATH_DECODE_RF_U1024 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4587, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4329, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6074);
   DLX_INST_DATA_PATH_DECODE_RF_U1023 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7030, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7062, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6074, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6069);
   DLX_INST_DATA_PATH_DECODE_RF_U1022 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4651, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4393, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6073);
   DLX_INST_DATA_PATH_DECODE_RF_U1021 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6902, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6966, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6073, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6070);
   DLX_INST_DATA_PATH_DECODE_RF_U1020 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4523, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4265, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6072);
   DLX_INST_DATA_PATH_DECODE_RF_U1019 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6998, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6934, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6072, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6071);
   DLX_INST_DATA_PATH_DECODE_RF_U1018 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6068, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6069, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6070, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6071, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4124);
   DLX_INST_DATA_PATH_DECODE_RF_U1017 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4554, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4296, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6067);
   DLX_INST_DATA_PATH_DECODE_RF_U1016 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6741, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6837, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6067, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6060);
   DLX_INST_DATA_PATH_DECODE_RF_U1015 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4682, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4200, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4456, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6066);
   DLX_INST_DATA_PATH_DECODE_RF_U1014 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6709, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6805, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6066, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6061);
   DLX_INST_DATA_PATH_DECODE_RF_U1013 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4490, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4232, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6065);
   DLX_INST_DATA_PATH_DECODE_RF_U1012 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6773, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6677, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6065, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6062);
   DLX_INST_DATA_PATH_DECODE_RF_U1011 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4714, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4168, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4424, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6064);
   DLX_INST_DATA_PATH_DECODE_RF_U1010 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6869, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6645, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6064, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6063);
   DLX_INST_DATA_PATH_DECODE_RF_U1009 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6060, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6061, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6062, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6063, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6058);
   DLX_INST_DATA_PATH_DECODE_RF_U1008 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4618, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4360, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6059);
   DLX_INST_DATA_PATH_DECODE_RF_U1007 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6058, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_26_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6059, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6051);
   DLX_INST_DATA_PATH_DECODE_RF_U1006 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4586, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4328, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6057);
   DLX_INST_DATA_PATH_DECODE_RF_U1005 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7029, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7061, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6057, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6052);
   DLX_INST_DATA_PATH_DECODE_RF_U1004 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4650, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4392, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6056);
   DLX_INST_DATA_PATH_DECODE_RF_U1003 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6901, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6965, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6056, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6053);
   DLX_INST_DATA_PATH_DECODE_RF_U1002 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4522, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4264, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6055);
   DLX_INST_DATA_PATH_DECODE_RF_U1001 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6997, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6933, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6055, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6054);
   DLX_INST_DATA_PATH_DECODE_RF_U1000 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6051, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6052, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6053, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6054, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4125);
   DLX_INST_DATA_PATH_DECODE_RF_U999 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4553, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4295, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6050);
   DLX_INST_DATA_PATH_DECODE_RF_U998 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6740, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6836, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6050, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6043);
   DLX_INST_DATA_PATH_DECODE_RF_U997 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4681, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4199, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4455, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6049);
   DLX_INST_DATA_PATH_DECODE_RF_U996 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6708, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6804, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6049, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6044);
   DLX_INST_DATA_PATH_DECODE_RF_U995 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4489, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4231, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6048);
   DLX_INST_DATA_PATH_DECODE_RF_U994 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6772, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6676, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6048, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6045);
   DLX_INST_DATA_PATH_DECODE_RF_U993 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4713, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4167, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4423, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6047);
   DLX_INST_DATA_PATH_DECODE_RF_U992 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6868, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6644, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6047, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6046);
   DLX_INST_DATA_PATH_DECODE_RF_U991 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6043, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6044, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6045, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6046, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6041);
   DLX_INST_DATA_PATH_DECODE_RF_U990 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4617, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4359, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6042);
   DLX_INST_DATA_PATH_DECODE_RF_U989 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6041, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_27_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6042, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6034);
   DLX_INST_DATA_PATH_DECODE_RF_U988 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4585, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4327, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6040);
   DLX_INST_DATA_PATH_DECODE_RF_U987 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7028, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7060, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6040, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6035);
   DLX_INST_DATA_PATH_DECODE_RF_U986 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4649, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4391, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6039);
   DLX_INST_DATA_PATH_DECODE_RF_U985 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6900, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6964, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6039, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6036);
   DLX_INST_DATA_PATH_DECODE_RF_U984 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4521, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4263, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6038);
   DLX_INST_DATA_PATH_DECODE_RF_U983 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6996, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6932, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6038, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6037);
   DLX_INST_DATA_PATH_DECODE_RF_U982 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6034, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6035, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6036, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6037, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4126);
   DLX_INST_DATA_PATH_DECODE_RF_U981 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4552, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4294, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6033);
   DLX_INST_DATA_PATH_DECODE_RF_U980 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6739, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6835, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6033, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6026);
   DLX_INST_DATA_PATH_DECODE_RF_U979 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4680, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4198, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4454, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6032);
   DLX_INST_DATA_PATH_DECODE_RF_U978 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6707, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6803, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6032, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6027);
   DLX_INST_DATA_PATH_DECODE_RF_U977 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4488, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4230, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6031);
   DLX_INST_DATA_PATH_DECODE_RF_U976 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6771, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6675, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6031, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6028);
   DLX_INST_DATA_PATH_DECODE_RF_U975 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4712, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4166, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4422, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6030);
   DLX_INST_DATA_PATH_DECODE_RF_U974 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6867, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6643, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6030, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6029);
   DLX_INST_DATA_PATH_DECODE_RF_U973 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6026, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6027, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6028, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6029, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6024);
   DLX_INST_DATA_PATH_DECODE_RF_U972 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4616, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6025);
   DLX_INST_DATA_PATH_DECODE_RF_U971 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6024, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_28_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6025, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6017);
   DLX_INST_DATA_PATH_DECODE_RF_U970 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4584, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4326, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6023);
   DLX_INST_DATA_PATH_DECODE_RF_U969 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7027, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7059, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6023, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6018);
   DLX_INST_DATA_PATH_DECODE_RF_U968 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4648, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4390, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6022);
   DLX_INST_DATA_PATH_DECODE_RF_U967 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6899, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6963, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6022, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6019);
   DLX_INST_DATA_PATH_DECODE_RF_U966 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4520, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4262, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6021);
   DLX_INST_DATA_PATH_DECODE_RF_U965 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6995, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6931, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6021, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6020);
   DLX_INST_DATA_PATH_DECODE_RF_U964 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6017, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6018, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6019, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6020, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4127);
   DLX_INST_DATA_PATH_DECODE_RF_U963 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4293, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6016);
   DLX_INST_DATA_PATH_DECODE_RF_U962 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6738, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6834, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6016, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6009);
   DLX_INST_DATA_PATH_DECODE_RF_U961 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4679, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4197, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4453, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6015);
   DLX_INST_DATA_PATH_DECODE_RF_U960 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6706, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6802, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6015, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6010);
   DLX_INST_DATA_PATH_DECODE_RF_U959 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4487, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4229, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6014);
   DLX_INST_DATA_PATH_DECODE_RF_U958 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6770, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6674, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6014, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6011);
   DLX_INST_DATA_PATH_DECODE_RF_U957 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4711, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4165, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4421, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6013);
   DLX_INST_DATA_PATH_DECODE_RF_U956 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6866, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6642, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6013, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6012);
   DLX_INST_DATA_PATH_DECODE_RF_U955 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6009, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6010, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6011, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6012, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6007);
   DLX_INST_DATA_PATH_DECODE_RF_U954 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4615, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6008);
   DLX_INST_DATA_PATH_DECODE_RF_U953 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6007, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_29_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6008, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6000);
   DLX_INST_DATA_PATH_DECODE_RF_U952 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4583, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4325, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6006);
   DLX_INST_DATA_PATH_DECODE_RF_U951 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7026, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7058, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6006, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6001);
   DLX_INST_DATA_PATH_DECODE_RF_U950 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4647, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4389, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6005);
   DLX_INST_DATA_PATH_DECODE_RF_U949 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6898, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6962, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6005, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6002);
   DLX_INST_DATA_PATH_DECODE_RF_U948 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4519, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4261, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6004);
   DLX_INST_DATA_PATH_DECODE_RF_U947 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6994, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6930, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6004, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6003);
   DLX_INST_DATA_PATH_DECODE_RF_U946 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6000, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6001, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6002, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6003, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4128);
   DLX_INST_DATA_PATH_DECODE_RF_U945 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4550, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4292, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5999);
   DLX_INST_DATA_PATH_DECODE_RF_U944 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6737, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6833, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5999, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5992);
   DLX_INST_DATA_PATH_DECODE_RF_U943 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4678, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4196, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4452, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5998);
   DLX_INST_DATA_PATH_DECODE_RF_U942 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6705, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6801, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5998, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5993);
   DLX_INST_DATA_PATH_DECODE_RF_U941 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4486, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4228, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5997);
   DLX_INST_DATA_PATH_DECODE_RF_U940 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6769, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6673, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5997, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5994);
   DLX_INST_DATA_PATH_DECODE_RF_U939 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4710, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4164, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4420, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5996);
   DLX_INST_DATA_PATH_DECODE_RF_U938 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6865, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6641, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5996, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5995);
   DLX_INST_DATA_PATH_DECODE_RF_U937 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5992, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5993, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5994, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5995, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5990);
   DLX_INST_DATA_PATH_DECODE_RF_U936 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4614, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4356, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5991);
   DLX_INST_DATA_PATH_DECODE_RF_U935 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5990, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_30_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5991, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5983);
   DLX_INST_DATA_PATH_DECODE_RF_U934 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4582, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4324, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5989);
   DLX_INST_DATA_PATH_DECODE_RF_U933 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7025, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7057, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5989, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5984);
   DLX_INST_DATA_PATH_DECODE_RF_U932 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4646, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5988);
   DLX_INST_DATA_PATH_DECODE_RF_U931 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6897, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6961, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5988, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5985);
   DLX_INST_DATA_PATH_DECODE_RF_U930 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4518, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4260, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5987);
   DLX_INST_DATA_PATH_DECODE_RF_U929 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6993, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6929, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5987, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5986);
   DLX_INST_DATA_PATH_DECODE_RF_U928 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5983, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5984, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5985, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5986, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4129);
   DLX_INST_DATA_PATH_DECODE_RF_U927 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4549, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4291, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5980);
   DLX_INST_DATA_PATH_DECODE_RF_U926 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6736, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6832, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5980, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5957);
   DLX_INST_DATA_PATH_DECODE_RF_U925 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4677, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4195, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4451, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5974);
   DLX_INST_DATA_PATH_DECODE_RF_U924 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6704, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6800, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5974, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5958);
   DLX_INST_DATA_PATH_DECODE_RF_U923 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4485, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4227, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5969);
   DLX_INST_DATA_PATH_DECODE_RF_U922 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6768, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6672, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5969, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5959);
   DLX_INST_DATA_PATH_DECODE_RF_U921 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4709, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4163, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4419, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5963);
   DLX_INST_DATA_PATH_DECODE_RF_U920 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6864, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6640, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5963, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5960);
   DLX_INST_DATA_PATH_DECODE_RF_U919 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5957, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5958, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5959, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5960, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5953);
   DLX_INST_DATA_PATH_DECODE_RF_U918 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4613, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4355, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5954);
   DLX_INST_DATA_PATH_DECODE_RF_U917 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5953, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190, C2 => 
                           DLX_INST_DATA_PATH_B_outs_31_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5954, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5933);
   DLX_INST_DATA_PATH_DECODE_RF_U916 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4581, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4323, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5949);
   DLX_INST_DATA_PATH_DECODE_RF_U915 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7024, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7056, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5949, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5934);
   DLX_INST_DATA_PATH_DECODE_RF_U914 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4645, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4387, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5944);
   DLX_INST_DATA_PATH_DECODE_RF_U913 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6896, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6960, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5944, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5935);
   DLX_INST_DATA_PATH_DECODE_RF_U912 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4517, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4259, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5939);
   DLX_INST_DATA_PATH_DECODE_RF_U911 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6992, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6928, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5939, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5936);
   DLX_INST_DATA_PATH_DECODE_RF_U910 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5933, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5934, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5935, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5936, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4130);
   DLX_INST_DATA_PATH_DECODE_RF_U909 : NOR2_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_25_port, A2 => 
                           DLX_INST_IR_OUT_signal_24_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5924);
   DLX_INST_DATA_PATH_DECODE_RF_U908 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_23_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5930);
   DLX_INST_DATA_PATH_DECODE_RF_U907 : NOR3_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_21_port, A2 => 
                           DLX_INST_IR_OUT_signal_22_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5930, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5904);
   DLX_INST_DATA_PATH_DECODE_RF_U906 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_24_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5932);
   DLX_INST_DATA_PATH_DECODE_RF_U905 : NOR2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5932, A2 => 
                           DLX_INST_IR_OUT_signal_25_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5925);
   DLX_INST_DATA_PATH_DECODE_RF_U904 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_22_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5929);
   DLX_INST_DATA_PATH_DECODE_RF_U903 : INV_X1 port map( A => 
                           DLX_INST_IR_OUT_signal_21_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5927);
   DLX_INST_DATA_PATH_DECODE_RF_U902 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5930, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5929, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5927, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5912);
   DLX_INST_DATA_PATH_DECODE_RF_U901 : AND2_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_25_port, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5932, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5915);
   DLX_INST_DATA_PATH_DECODE_RF_U900 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5930, A2 => 
                           DLX_INST_IR_OUT_signal_22_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5927, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5910);
   DLX_INST_DATA_PATH_DECODE_RF_U899 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4580, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4322, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5931);
   DLX_INST_DATA_PATH_DECODE_RF_U898 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6767, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6863, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5931, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5919);
   DLX_INST_DATA_PATH_DECODE_RF_U897 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5929, A2 => 
                           DLX_INST_IR_OUT_signal_23_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5927, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5914);
   DLX_INST_DATA_PATH_DECODE_RF_U896 : NOR3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5929, A2 => 
                           DLX_INST_IR_OUT_signal_21_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5930, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5908);
   DLX_INST_DATA_PATH_DECODE_RF_U895 : NOR3_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_21_port, A2 => 
                           DLX_INST_IR_OUT_signal_23_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5929, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5913);
   DLX_INST_DATA_PATH_DECODE_RF_U894 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4708, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4226, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4482, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5928);
   DLX_INST_DATA_PATH_DECODE_RF_U893 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6735, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6831, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5928, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5920);
   DLX_INST_DATA_PATH_DECODE_RF_U892 : NOR3_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_22_port, A2 => 
                           DLX_INST_IR_OUT_signal_23_port, A3 => 
                           DLX_INST_IR_OUT_signal_21_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5907);
   DLX_INST_DATA_PATH_DECODE_RF_U891 : NOR3_X1 port map( A1 => 
                           DLX_INST_IR_OUT_signal_22_port, A2 => 
                           DLX_INST_IR_OUT_signal_23_port, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5927, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5906);
   DLX_INST_DATA_PATH_DECODE_RF_U890 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4516, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4258, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5926);
   DLX_INST_DATA_PATH_DECODE_RF_U889 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6799, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6703, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5926, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5921);
   DLX_INST_DATA_PATH_DECODE_RF_U888 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4740, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4194, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4450, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5923);
   DLX_INST_DATA_PATH_DECODE_RF_U887 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6895, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6671, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5923, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5922);
   DLX_INST_DATA_PATH_DECODE_RF_U886 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5919, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5920, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5921, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5922, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5917);
   DLX_INST_DATA_PATH_DECODE_RF_U885 : AND3_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, A2 => 
                           DLX_INST_IR_OUT_signal_25_port, A3 => 
                           DLX_INST_IR_OUT_signal_24_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5911);
   DLX_INST_DATA_PATH_DECODE_RF_U884 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4644, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4386, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5918);
   DLX_INST_DATA_PATH_DECODE_RF_U883 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5917, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_0_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5918, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5899);
   DLX_INST_DATA_PATH_DECODE_RF_U882 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4612, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4354, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5916);
   DLX_INST_DATA_PATH_DECODE_RF_U881 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7055, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7087, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5916, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5900);
   DLX_INST_DATA_PATH_DECODE_RF_U880 : AND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5915, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5905);
   DLX_INST_DATA_PATH_DECODE_RF_U879 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4676, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4418, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5909);
   DLX_INST_DATA_PATH_DECODE_RF_U878 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6927, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6991, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5909, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5901);
   DLX_INST_DATA_PATH_DECODE_RF_U877 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4548, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4290, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5903);
   DLX_INST_DATA_PATH_DECODE_RF_U876 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7023, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6959, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5903, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5902);
   DLX_INST_DATA_PATH_DECODE_RF_U875 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5899, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5900, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5901, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5902, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4131);
   DLX_INST_DATA_PATH_DECODE_RF_U874 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4579, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4321, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5898);
   DLX_INST_DATA_PATH_DECODE_RF_U873 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6766, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6862, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5898, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5891);
   DLX_INST_DATA_PATH_DECODE_RF_U872 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4707, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4225, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4481, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5897);
   DLX_INST_DATA_PATH_DECODE_RF_U871 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6734, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6830, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5897, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5892);
   DLX_INST_DATA_PATH_DECODE_RF_U870 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4515, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4257, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5896);
   DLX_INST_DATA_PATH_DECODE_RF_U869 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6798, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6702, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5896, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5893);
   DLX_INST_DATA_PATH_DECODE_RF_U868 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4739, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4193, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4449, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5895);
   DLX_INST_DATA_PATH_DECODE_RF_U867 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6894, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6670, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5895, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5894);
   DLX_INST_DATA_PATH_DECODE_RF_U866 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5891, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5892, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5893, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5894, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5889);
   DLX_INST_DATA_PATH_DECODE_RF_U865 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4643, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4385, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5890);
   DLX_INST_DATA_PATH_DECODE_RF_U864 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5889, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_1_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5890, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5882);
   DLX_INST_DATA_PATH_DECODE_RF_U863 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4611, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4353, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5888);
   DLX_INST_DATA_PATH_DECODE_RF_U862 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7054, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7086, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5888, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5883);
   DLX_INST_DATA_PATH_DECODE_RF_U861 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4675, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4417, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5887);
   DLX_INST_DATA_PATH_DECODE_RF_U860 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6926, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6990, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5887, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5884);
   DLX_INST_DATA_PATH_DECODE_RF_U859 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4547, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4289, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5886);
   DLX_INST_DATA_PATH_DECODE_RF_U858 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7022, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6958, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5886, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5885);
   DLX_INST_DATA_PATH_DECODE_RF_U857 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5882, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5883, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5884, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5885, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4132);
   DLX_INST_DATA_PATH_DECODE_RF_U856 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4578, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4320, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5881);
   DLX_INST_DATA_PATH_DECODE_RF_U855 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6765, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6861, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5881, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5874);
   DLX_INST_DATA_PATH_DECODE_RF_U854 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4706, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4224, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4480, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5880);
   DLX_INST_DATA_PATH_DECODE_RF_U853 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6733, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6829, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5880, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5875);
   DLX_INST_DATA_PATH_DECODE_RF_U852 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4514, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4256, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5879);
   DLX_INST_DATA_PATH_DECODE_RF_U851 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6797, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6701, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5879, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5876);
   DLX_INST_DATA_PATH_DECODE_RF_U850 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4738, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4192, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4448, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5878);
   DLX_INST_DATA_PATH_DECODE_RF_U849 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6893, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6669, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5878, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5877);
   DLX_INST_DATA_PATH_DECODE_RF_U848 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5874, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5875, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5876, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5877, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5872);
   DLX_INST_DATA_PATH_DECODE_RF_U847 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4642, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4384, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5873);
   DLX_INST_DATA_PATH_DECODE_RF_U846 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5872, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_2_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5873, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5865);
   DLX_INST_DATA_PATH_DECODE_RF_U845 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4610, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4352, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5871);
   DLX_INST_DATA_PATH_DECODE_RF_U844 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7053, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7085, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5871, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5866);
   DLX_INST_DATA_PATH_DECODE_RF_U843 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4674, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4416, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5870);
   DLX_INST_DATA_PATH_DECODE_RF_U842 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6925, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6989, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5870, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5867);
   DLX_INST_DATA_PATH_DECODE_RF_U841 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4546, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4288, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5869);
   DLX_INST_DATA_PATH_DECODE_RF_U840 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7021, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6957, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5869, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5868);
   DLX_INST_DATA_PATH_DECODE_RF_U839 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5865, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5866, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5867, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5868, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4133);
   DLX_INST_DATA_PATH_DECODE_RF_U838 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4577, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4319, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5864);
   DLX_INST_DATA_PATH_DECODE_RF_U837 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6764, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6860, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5864, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5857);
   DLX_INST_DATA_PATH_DECODE_RF_U836 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4705, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4223, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4479, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5863);
   DLX_INST_DATA_PATH_DECODE_RF_U835 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6732, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6828, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5863, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5858);
   DLX_INST_DATA_PATH_DECODE_RF_U834 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4513, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4255, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5862);
   DLX_INST_DATA_PATH_DECODE_RF_U833 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6796, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6700, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5862, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5859);
   DLX_INST_DATA_PATH_DECODE_RF_U832 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4737, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4191, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4447, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5861);
   DLX_INST_DATA_PATH_DECODE_RF_U831 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6892, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6668, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5861, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5860);
   DLX_INST_DATA_PATH_DECODE_RF_U830 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5857, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5858, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5859, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5860, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5855);
   DLX_INST_DATA_PATH_DECODE_RF_U829 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4641, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4383, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5856);
   DLX_INST_DATA_PATH_DECODE_RF_U828 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5855, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_3_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5856, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5848);
   DLX_INST_DATA_PATH_DECODE_RF_U827 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4609, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4351, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5854);
   DLX_INST_DATA_PATH_DECODE_RF_U826 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7052, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7084, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5854, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5849);
   DLX_INST_DATA_PATH_DECODE_RF_U825 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4673, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4415, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5853);
   DLX_INST_DATA_PATH_DECODE_RF_U824 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6924, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6988, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5853, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5850);
   DLX_INST_DATA_PATH_DECODE_RF_U823 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4545, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4287, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5852);
   DLX_INST_DATA_PATH_DECODE_RF_U822 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7020, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6956, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5852, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5851);
   DLX_INST_DATA_PATH_DECODE_RF_U821 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5848, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5849, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5850, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5851, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4134);
   DLX_INST_DATA_PATH_DECODE_RF_U820 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4576, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4318, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5847);
   DLX_INST_DATA_PATH_DECODE_RF_U819 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6763, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6859, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5847, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5840);
   DLX_INST_DATA_PATH_DECODE_RF_U818 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4704, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4222, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4478, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5846);
   DLX_INST_DATA_PATH_DECODE_RF_U817 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6731, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6827, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5846, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5841);
   DLX_INST_DATA_PATH_DECODE_RF_U816 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4512, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4254, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5845);
   DLX_INST_DATA_PATH_DECODE_RF_U815 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6795, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6699, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5845, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5842);
   DLX_INST_DATA_PATH_DECODE_RF_U814 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4736, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4190, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4446, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5844);
   DLX_INST_DATA_PATH_DECODE_RF_U813 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6891, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6667, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5844, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5843);
   DLX_INST_DATA_PATH_DECODE_RF_U812 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5840, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5841, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5842, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5843, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5838);
   DLX_INST_DATA_PATH_DECODE_RF_U811 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4640, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4382, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5839);
   DLX_INST_DATA_PATH_DECODE_RF_U810 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5838, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_4_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5839, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5831);
   DLX_INST_DATA_PATH_DECODE_RF_U809 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4608, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4350, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5837);
   DLX_INST_DATA_PATH_DECODE_RF_U808 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7051, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7083, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5837, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5832);
   DLX_INST_DATA_PATH_DECODE_RF_U807 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4672, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4414, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5836);
   DLX_INST_DATA_PATH_DECODE_RF_U806 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6923, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6987, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5836, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5833);
   DLX_INST_DATA_PATH_DECODE_RF_U805 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4544, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4286, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5835);
   DLX_INST_DATA_PATH_DECODE_RF_U804 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7019, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6955, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5835, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5834);
   DLX_INST_DATA_PATH_DECODE_RF_U803 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5831, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5832, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5833, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5834, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4135);
   DLX_INST_DATA_PATH_DECODE_RF_U802 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4575, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4317, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5830);
   DLX_INST_DATA_PATH_DECODE_RF_U801 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6762, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6858, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5830, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5823);
   DLX_INST_DATA_PATH_DECODE_RF_U800 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4703, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4221, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4477, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5829);
   DLX_INST_DATA_PATH_DECODE_RF_U799 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6730, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6826, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5829, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5824);
   DLX_INST_DATA_PATH_DECODE_RF_U798 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4511, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4253, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5828);
   DLX_INST_DATA_PATH_DECODE_RF_U797 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6794, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6698, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5828, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5825);
   DLX_INST_DATA_PATH_DECODE_RF_U796 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4735, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4189, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4445, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5827);
   DLX_INST_DATA_PATH_DECODE_RF_U795 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6890, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6666, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5827, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5826);
   DLX_INST_DATA_PATH_DECODE_RF_U794 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5823, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5824, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5825, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5826, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5821);
   DLX_INST_DATA_PATH_DECODE_RF_U793 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4639, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4381, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5822);
   DLX_INST_DATA_PATH_DECODE_RF_U792 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5821, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_5_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5822, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5814);
   DLX_INST_DATA_PATH_DECODE_RF_U791 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4607, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4349, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5820);
   DLX_INST_DATA_PATH_DECODE_RF_U790 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7050, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7082, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5820, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5815);
   DLX_INST_DATA_PATH_DECODE_RF_U789 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4671, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4413, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5819);
   DLX_INST_DATA_PATH_DECODE_RF_U788 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6922, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6986, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5819, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5816);
   DLX_INST_DATA_PATH_DECODE_RF_U787 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4543, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4285, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5818);
   DLX_INST_DATA_PATH_DECODE_RF_U786 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7018, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6954, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5818, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5817);
   DLX_INST_DATA_PATH_DECODE_RF_U785 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5814, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5815, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5816, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5817, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4136);
   DLX_INST_DATA_PATH_DECODE_RF_U784 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4574, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4316, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5813);
   DLX_INST_DATA_PATH_DECODE_RF_U783 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6761, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6857, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5813, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5806);
   DLX_INST_DATA_PATH_DECODE_RF_U782 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4702, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4220, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4476, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5812);
   DLX_INST_DATA_PATH_DECODE_RF_U781 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6729, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6825, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5812, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5807);
   DLX_INST_DATA_PATH_DECODE_RF_U780 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4510, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4252, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5811);
   DLX_INST_DATA_PATH_DECODE_RF_U779 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6793, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6697, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5811, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5808);
   DLX_INST_DATA_PATH_DECODE_RF_U778 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4734, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4188, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4444, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5810);
   DLX_INST_DATA_PATH_DECODE_RF_U777 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6889, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6665, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5810, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5809);
   DLX_INST_DATA_PATH_DECODE_RF_U776 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5806, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5807, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5808, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5809, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5804);
   DLX_INST_DATA_PATH_DECODE_RF_U775 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4638, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4380, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5805);
   DLX_INST_DATA_PATH_DECODE_RF_U774 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5804, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_6_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5805, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5797);
   DLX_INST_DATA_PATH_DECODE_RF_U773 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4606, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4348, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5803);
   DLX_INST_DATA_PATH_DECODE_RF_U772 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7049, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7081, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5803, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5798);
   DLX_INST_DATA_PATH_DECODE_RF_U771 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4670, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4412, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5802);
   DLX_INST_DATA_PATH_DECODE_RF_U770 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6921, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6985, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5802, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5799);
   DLX_INST_DATA_PATH_DECODE_RF_U769 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4542, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4284, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5801);
   DLX_INST_DATA_PATH_DECODE_RF_U768 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7017, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6953, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5801, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5800);
   DLX_INST_DATA_PATH_DECODE_RF_U767 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5797, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5798, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5799, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5800, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4137);
   DLX_INST_DATA_PATH_DECODE_RF_U766 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4573, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4315, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5796);
   DLX_INST_DATA_PATH_DECODE_RF_U765 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6760, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6856, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5796, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5789);
   DLX_INST_DATA_PATH_DECODE_RF_U764 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4701, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4219, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4475, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5795);
   DLX_INST_DATA_PATH_DECODE_RF_U763 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6728, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6824, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5795, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5790);
   DLX_INST_DATA_PATH_DECODE_RF_U762 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4509, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4251, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5794);
   DLX_INST_DATA_PATH_DECODE_RF_U761 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6792, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6696, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5794, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5791);
   DLX_INST_DATA_PATH_DECODE_RF_U760 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4733, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4187, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4443, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5793);
   DLX_INST_DATA_PATH_DECODE_RF_U759 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6888, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6664, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5793, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5792);
   DLX_INST_DATA_PATH_DECODE_RF_U758 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5789, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5790, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5791, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5792, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5787);
   DLX_INST_DATA_PATH_DECODE_RF_U757 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4637, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4379, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5788);
   DLX_INST_DATA_PATH_DECODE_RF_U756 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5787, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_7_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5788, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5780);
   DLX_INST_DATA_PATH_DECODE_RF_U755 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4605, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4347, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5786);
   DLX_INST_DATA_PATH_DECODE_RF_U754 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7048, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7080, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5786, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5781);
   DLX_INST_DATA_PATH_DECODE_RF_U753 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4669, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4411, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5785);
   DLX_INST_DATA_PATH_DECODE_RF_U752 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6920, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6984, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5785, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5782);
   DLX_INST_DATA_PATH_DECODE_RF_U751 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4541, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4283, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5784);
   DLX_INST_DATA_PATH_DECODE_RF_U750 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7016, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6952, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5784, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5783);
   DLX_INST_DATA_PATH_DECODE_RF_U749 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5780, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5781, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5782, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5783, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4138);
   DLX_INST_DATA_PATH_DECODE_RF_U748 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4572, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4314, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5779);
   DLX_INST_DATA_PATH_DECODE_RF_U747 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6759, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6855, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5779, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5772);
   DLX_INST_DATA_PATH_DECODE_RF_U746 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4700, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4218, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4474, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5778);
   DLX_INST_DATA_PATH_DECODE_RF_U745 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6727, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6823, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5778, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5773);
   DLX_INST_DATA_PATH_DECODE_RF_U744 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4508, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4250, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5777);
   DLX_INST_DATA_PATH_DECODE_RF_U743 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6791, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6695, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5777, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5774);
   DLX_INST_DATA_PATH_DECODE_RF_U742 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4732, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4186, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4442, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5776);
   DLX_INST_DATA_PATH_DECODE_RF_U741 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6887, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6663, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5776, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5775);
   DLX_INST_DATA_PATH_DECODE_RF_U740 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5772, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5773, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5774, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5775, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5770);
   DLX_INST_DATA_PATH_DECODE_RF_U739 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4636, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4378, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5771);
   DLX_INST_DATA_PATH_DECODE_RF_U738 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5770, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_8_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5771, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5763);
   DLX_INST_DATA_PATH_DECODE_RF_U737 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4604, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4346, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5769);
   DLX_INST_DATA_PATH_DECODE_RF_U736 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7047, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7079, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5769, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5764);
   DLX_INST_DATA_PATH_DECODE_RF_U735 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4668, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4410, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5768);
   DLX_INST_DATA_PATH_DECODE_RF_U734 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6919, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6983, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5768, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5765);
   DLX_INST_DATA_PATH_DECODE_RF_U733 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4540, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4282, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5767);
   DLX_INST_DATA_PATH_DECODE_RF_U732 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7015, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6951, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5767, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5766);
   DLX_INST_DATA_PATH_DECODE_RF_U731 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5763, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5764, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5765, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5766, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4139);
   DLX_INST_DATA_PATH_DECODE_RF_U730 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4571, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4313, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5762);
   DLX_INST_DATA_PATH_DECODE_RF_U729 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6758, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6854, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5762, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5755);
   DLX_INST_DATA_PATH_DECODE_RF_U728 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4699, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4217, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4473, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5761);
   DLX_INST_DATA_PATH_DECODE_RF_U727 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6726, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6822, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5761, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5756);
   DLX_INST_DATA_PATH_DECODE_RF_U726 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4507, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4249, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5760);
   DLX_INST_DATA_PATH_DECODE_RF_U725 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6790, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6694, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5760, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5757);
   DLX_INST_DATA_PATH_DECODE_RF_U724 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4731, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4185, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4441, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5759);
   DLX_INST_DATA_PATH_DECODE_RF_U723 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6886, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6662, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5759, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5758);
   DLX_INST_DATA_PATH_DECODE_RF_U722 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5755, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5756, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5757, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5758, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5753);
   DLX_INST_DATA_PATH_DECODE_RF_U721 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4635, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4377, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5754);
   DLX_INST_DATA_PATH_DECODE_RF_U720 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5753, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_9_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5754, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5746);
   DLX_INST_DATA_PATH_DECODE_RF_U719 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4603, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4345, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5752);
   DLX_INST_DATA_PATH_DECODE_RF_U718 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7046, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7078, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5752, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5747);
   DLX_INST_DATA_PATH_DECODE_RF_U717 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4667, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4409, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5751);
   DLX_INST_DATA_PATH_DECODE_RF_U716 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6918, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6982, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5751, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5748);
   DLX_INST_DATA_PATH_DECODE_RF_U715 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4539, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4281, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5750);
   DLX_INST_DATA_PATH_DECODE_RF_U714 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7014, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6950, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5750, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5749);
   DLX_INST_DATA_PATH_DECODE_RF_U713 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5746, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5747, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5748, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5749, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4140);
   DLX_INST_DATA_PATH_DECODE_RF_U712 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4570, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4312, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5745);
   DLX_INST_DATA_PATH_DECODE_RF_U711 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6757, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6853, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5745, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5738);
   DLX_INST_DATA_PATH_DECODE_RF_U710 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4698, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4216, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4472, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5744);
   DLX_INST_DATA_PATH_DECODE_RF_U709 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6725, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6821, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5744, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5739);
   DLX_INST_DATA_PATH_DECODE_RF_U708 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4506, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4248, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5743);
   DLX_INST_DATA_PATH_DECODE_RF_U707 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6789, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6693, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5743, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5740);
   DLX_INST_DATA_PATH_DECODE_RF_U706 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4730, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4184, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4440, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5742);
   DLX_INST_DATA_PATH_DECODE_RF_U705 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6885, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6661, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5742, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5741);
   DLX_INST_DATA_PATH_DECODE_RF_U704 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5738, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5739, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5740, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5741, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5736);
   DLX_INST_DATA_PATH_DECODE_RF_U703 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4634, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4376, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5737);
   DLX_INST_DATA_PATH_DECODE_RF_U702 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5736, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_10_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5737, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5729);
   DLX_INST_DATA_PATH_DECODE_RF_U701 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4602, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4344, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5735);
   DLX_INST_DATA_PATH_DECODE_RF_U700 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7045, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7077, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5735, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5730);
   DLX_INST_DATA_PATH_DECODE_RF_U699 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4666, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4408, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5734);
   DLX_INST_DATA_PATH_DECODE_RF_U698 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6917, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6981, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5734, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5731);
   DLX_INST_DATA_PATH_DECODE_RF_U697 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4538, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4280, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5733);
   DLX_INST_DATA_PATH_DECODE_RF_U696 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7013, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6949, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5733, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5732);
   DLX_INST_DATA_PATH_DECODE_RF_U695 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5729, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5730, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5731, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5732, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4141);
   DLX_INST_DATA_PATH_DECODE_RF_U694 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4569, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4311, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5728);
   DLX_INST_DATA_PATH_DECODE_RF_U693 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6756, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6852, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5728, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5721);
   DLX_INST_DATA_PATH_DECODE_RF_U692 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4697, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4215, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4471, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5727);
   DLX_INST_DATA_PATH_DECODE_RF_U691 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6724, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6820, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5727, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5722);
   DLX_INST_DATA_PATH_DECODE_RF_U690 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4505, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4247, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5726);
   DLX_INST_DATA_PATH_DECODE_RF_U689 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6788, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6692, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5726, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5723);
   DLX_INST_DATA_PATH_DECODE_RF_U688 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4729, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4183, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4439, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5725);
   DLX_INST_DATA_PATH_DECODE_RF_U687 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6884, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6660, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5725, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5724);
   DLX_INST_DATA_PATH_DECODE_RF_U686 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5721, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5722, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5723, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5724, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5719);
   DLX_INST_DATA_PATH_DECODE_RF_U685 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4633, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4375, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5720);
   DLX_INST_DATA_PATH_DECODE_RF_U684 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5719, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_11_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5720, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5712);
   DLX_INST_DATA_PATH_DECODE_RF_U683 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4601, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4343, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5718);
   DLX_INST_DATA_PATH_DECODE_RF_U682 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7044, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7076, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5718, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5713);
   DLX_INST_DATA_PATH_DECODE_RF_U681 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4665, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4407, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5717);
   DLX_INST_DATA_PATH_DECODE_RF_U680 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6916, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6980, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5717, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5714);
   DLX_INST_DATA_PATH_DECODE_RF_U679 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4537, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4279, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5716);
   DLX_INST_DATA_PATH_DECODE_RF_U678 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7012, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6948, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5716, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5715);
   DLX_INST_DATA_PATH_DECODE_RF_U677 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5712, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5713, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5714, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5715, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4142);
   DLX_INST_DATA_PATH_DECODE_RF_U676 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4568, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4310, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5711);
   DLX_INST_DATA_PATH_DECODE_RF_U675 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6755, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6851, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5711, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5704);
   DLX_INST_DATA_PATH_DECODE_RF_U674 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4696, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4214, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4470, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5710);
   DLX_INST_DATA_PATH_DECODE_RF_U673 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6723, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6819, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5710, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5705);
   DLX_INST_DATA_PATH_DECODE_RF_U672 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4504, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4246, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5709);
   DLX_INST_DATA_PATH_DECODE_RF_U671 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6787, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6691, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5709, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5706);
   DLX_INST_DATA_PATH_DECODE_RF_U670 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4728, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4182, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4438, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5708);
   DLX_INST_DATA_PATH_DECODE_RF_U669 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6883, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6659, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5708, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5707);
   DLX_INST_DATA_PATH_DECODE_RF_U668 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5704, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5705, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5706, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5707, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5702);
   DLX_INST_DATA_PATH_DECODE_RF_U667 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4632, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4374, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5703);
   DLX_INST_DATA_PATH_DECODE_RF_U666 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5702, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_12_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5703, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5695);
   DLX_INST_DATA_PATH_DECODE_RF_U665 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4600, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4342, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5701);
   DLX_INST_DATA_PATH_DECODE_RF_U664 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7043, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7075, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5701, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5696);
   DLX_INST_DATA_PATH_DECODE_RF_U663 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4664, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4406, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5700);
   DLX_INST_DATA_PATH_DECODE_RF_U662 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6915, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6979, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5700, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5697);
   DLX_INST_DATA_PATH_DECODE_RF_U661 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4536, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4278, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5699);
   DLX_INST_DATA_PATH_DECODE_RF_U660 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7011, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6947, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5699, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5698);
   DLX_INST_DATA_PATH_DECODE_RF_U659 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5695, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5696, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5697, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5698, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4143);
   DLX_INST_DATA_PATH_DECODE_RF_U658 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4567, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4309, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5694);
   DLX_INST_DATA_PATH_DECODE_RF_U657 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6754, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6850, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5694, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5687);
   DLX_INST_DATA_PATH_DECODE_RF_U656 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4695, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4213, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4469, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5693);
   DLX_INST_DATA_PATH_DECODE_RF_U655 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6722, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6818, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5693, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5688);
   DLX_INST_DATA_PATH_DECODE_RF_U654 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4503, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4245, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5692);
   DLX_INST_DATA_PATH_DECODE_RF_U653 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6786, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6690, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5692, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5689);
   DLX_INST_DATA_PATH_DECODE_RF_U652 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4727, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4181, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4437, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5691);
   DLX_INST_DATA_PATH_DECODE_RF_U651 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6882, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6658, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5691, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5690);
   DLX_INST_DATA_PATH_DECODE_RF_U650 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5687, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5688, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5689, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5690, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5685);
   DLX_INST_DATA_PATH_DECODE_RF_U649 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4631, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4373, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5686);
   DLX_INST_DATA_PATH_DECODE_RF_U648 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5685, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_13_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5686, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5678);
   DLX_INST_DATA_PATH_DECODE_RF_U647 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4599, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4341, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5684);
   DLX_INST_DATA_PATH_DECODE_RF_U646 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7042, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7074, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5684, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5679);
   DLX_INST_DATA_PATH_DECODE_RF_U645 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4663, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4405, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5683);
   DLX_INST_DATA_PATH_DECODE_RF_U644 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6914, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6978, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5683, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5680);
   DLX_INST_DATA_PATH_DECODE_RF_U643 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4535, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4277, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5682);
   DLX_INST_DATA_PATH_DECODE_RF_U642 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7010, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6946, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5682, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5681);
   DLX_INST_DATA_PATH_DECODE_RF_U641 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5678, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5679, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5680, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5681, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4144);
   DLX_INST_DATA_PATH_DECODE_RF_U640 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4566, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4308, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5677);
   DLX_INST_DATA_PATH_DECODE_RF_U639 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6753, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6849, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5677, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5670);
   DLX_INST_DATA_PATH_DECODE_RF_U638 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4694, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4212, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4468, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5676);
   DLX_INST_DATA_PATH_DECODE_RF_U637 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6721, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6817, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5676, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5671);
   DLX_INST_DATA_PATH_DECODE_RF_U636 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4502, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4244, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5675);
   DLX_INST_DATA_PATH_DECODE_RF_U635 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6785, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6689, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5675, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5672);
   DLX_INST_DATA_PATH_DECODE_RF_U634 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4726, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4180, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4436, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5674);
   DLX_INST_DATA_PATH_DECODE_RF_U633 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6881, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6657, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5674, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5673);
   DLX_INST_DATA_PATH_DECODE_RF_U632 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5670, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5671, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5672, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5673, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5668);
   DLX_INST_DATA_PATH_DECODE_RF_U631 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4630, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4372, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5669);
   DLX_INST_DATA_PATH_DECODE_RF_U630 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5668, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_14_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5669, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5661);
   DLX_INST_DATA_PATH_DECODE_RF_U629 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4598, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4340, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5667);
   DLX_INST_DATA_PATH_DECODE_RF_U628 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7041, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7073, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5667, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5662);
   DLX_INST_DATA_PATH_DECODE_RF_U627 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4662, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4404, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5666);
   DLX_INST_DATA_PATH_DECODE_RF_U626 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6913, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6977, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5666, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5663);
   DLX_INST_DATA_PATH_DECODE_RF_U625 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4534, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4276, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5665);
   DLX_INST_DATA_PATH_DECODE_RF_U624 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7009, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6945, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5665, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5664);
   DLX_INST_DATA_PATH_DECODE_RF_U623 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5661, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5662, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5663, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5664, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4145);
   DLX_INST_DATA_PATH_DECODE_RF_U622 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4565, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4307, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5660);
   DLX_INST_DATA_PATH_DECODE_RF_U621 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6752, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6848, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5660, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5653);
   DLX_INST_DATA_PATH_DECODE_RF_U620 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4693, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4211, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4467, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5659);
   DLX_INST_DATA_PATH_DECODE_RF_U619 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6720, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6816, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5659, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5654);
   DLX_INST_DATA_PATH_DECODE_RF_U618 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4501, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4243, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5658);
   DLX_INST_DATA_PATH_DECODE_RF_U617 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6784, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6688, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5658, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5655);
   DLX_INST_DATA_PATH_DECODE_RF_U616 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4725, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4179, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4435, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5657);
   DLX_INST_DATA_PATH_DECODE_RF_U615 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6880, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6656, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5657, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5656);
   DLX_INST_DATA_PATH_DECODE_RF_U614 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5653, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5654, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5655, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5656, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5651);
   DLX_INST_DATA_PATH_DECODE_RF_U613 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4629, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4371, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5652);
   DLX_INST_DATA_PATH_DECODE_RF_U612 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5651, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_15_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5652, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5644);
   DLX_INST_DATA_PATH_DECODE_RF_U611 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4597, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4339, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5650);
   DLX_INST_DATA_PATH_DECODE_RF_U610 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7040, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7072, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5650, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5645);
   DLX_INST_DATA_PATH_DECODE_RF_U609 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4661, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4403, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5649);
   DLX_INST_DATA_PATH_DECODE_RF_U608 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6912, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6976, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5649, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5646);
   DLX_INST_DATA_PATH_DECODE_RF_U607 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4533, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4275, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5648);
   DLX_INST_DATA_PATH_DECODE_RF_U606 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7008, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6944, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5648, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5647);
   DLX_INST_DATA_PATH_DECODE_RF_U605 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5644, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5645, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5646, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5647, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4146);
   DLX_INST_DATA_PATH_DECODE_RF_U604 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4564, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4306, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5643);
   DLX_INST_DATA_PATH_DECODE_RF_U603 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6751, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6847, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5643, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5636);
   DLX_INST_DATA_PATH_DECODE_RF_U602 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4692, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4210, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4466, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5642);
   DLX_INST_DATA_PATH_DECODE_RF_U601 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6719, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6815, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5642, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5637);
   DLX_INST_DATA_PATH_DECODE_RF_U600 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4500, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4242, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5641);
   DLX_INST_DATA_PATH_DECODE_RF_U599 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6783, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6687, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5641, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5638);
   DLX_INST_DATA_PATH_DECODE_RF_U598 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4724, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4178, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4434, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5640);
   DLX_INST_DATA_PATH_DECODE_RF_U597 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6879, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6655, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5640, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5639);
   DLX_INST_DATA_PATH_DECODE_RF_U596 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5636, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5637, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5638, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5639, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5634);
   DLX_INST_DATA_PATH_DECODE_RF_U595 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4628, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4370, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5635);
   DLX_INST_DATA_PATH_DECODE_RF_U594 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5634, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_16_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5635, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5627);
   DLX_INST_DATA_PATH_DECODE_RF_U593 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4596, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4338, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5633);
   DLX_INST_DATA_PATH_DECODE_RF_U592 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7039, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7071, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5633, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5628);
   DLX_INST_DATA_PATH_DECODE_RF_U591 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4660, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4402, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5632);
   DLX_INST_DATA_PATH_DECODE_RF_U590 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6911, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6975, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5632, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5629);
   DLX_INST_DATA_PATH_DECODE_RF_U589 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4532, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4274, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5631);
   DLX_INST_DATA_PATH_DECODE_RF_U588 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7007, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6943, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5631, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5630);
   DLX_INST_DATA_PATH_DECODE_RF_U587 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5627, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5628, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5629, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5630, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4147);
   DLX_INST_DATA_PATH_DECODE_RF_U586 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4563, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4305, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5626);
   DLX_INST_DATA_PATH_DECODE_RF_U585 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6750, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6846, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5626, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5619);
   DLX_INST_DATA_PATH_DECODE_RF_U584 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4691, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4209, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4465, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5625);
   DLX_INST_DATA_PATH_DECODE_RF_U583 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6718, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6814, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5625, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5620);
   DLX_INST_DATA_PATH_DECODE_RF_U582 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4499, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4241, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5624);
   DLX_INST_DATA_PATH_DECODE_RF_U581 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6782, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6686, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5624, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5621);
   DLX_INST_DATA_PATH_DECODE_RF_U580 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4723, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4177, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4433, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5623);
   DLX_INST_DATA_PATH_DECODE_RF_U579 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6878, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6654, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5623, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5622);
   DLX_INST_DATA_PATH_DECODE_RF_U578 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5619, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5620, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5621, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5622, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5617);
   DLX_INST_DATA_PATH_DECODE_RF_U577 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4627, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4369, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5618);
   DLX_INST_DATA_PATH_DECODE_RF_U576 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5617, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_17_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5618, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5610);
   DLX_INST_DATA_PATH_DECODE_RF_U575 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4595, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4337, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5616);
   DLX_INST_DATA_PATH_DECODE_RF_U574 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7038, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7070, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5616, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5611);
   DLX_INST_DATA_PATH_DECODE_RF_U573 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4659, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4401, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5615);
   DLX_INST_DATA_PATH_DECODE_RF_U572 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6910, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6974, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5615, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5612);
   DLX_INST_DATA_PATH_DECODE_RF_U571 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4531, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4273, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5614);
   DLX_INST_DATA_PATH_DECODE_RF_U570 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7006, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6942, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5614, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5613);
   DLX_INST_DATA_PATH_DECODE_RF_U569 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5610, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5611, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5612, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5613, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4148);
   DLX_INST_DATA_PATH_DECODE_RF_U568 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4562, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4304, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5609);
   DLX_INST_DATA_PATH_DECODE_RF_U567 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6749, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6845, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5609, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5602);
   DLX_INST_DATA_PATH_DECODE_RF_U566 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4690, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4208, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4464, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5608);
   DLX_INST_DATA_PATH_DECODE_RF_U565 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6717, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6813, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5608, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5603);
   DLX_INST_DATA_PATH_DECODE_RF_U564 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4498, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4240, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5607);
   DLX_INST_DATA_PATH_DECODE_RF_U563 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6781, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6685, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5607, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5604);
   DLX_INST_DATA_PATH_DECODE_RF_U562 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4722, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4176, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4432, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5606);
   DLX_INST_DATA_PATH_DECODE_RF_U561 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6877, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6653, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5606, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5605);
   DLX_INST_DATA_PATH_DECODE_RF_U560 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5602, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5603, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5604, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5605, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5600);
   DLX_INST_DATA_PATH_DECODE_RF_U559 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4626, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4368, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5601);
   DLX_INST_DATA_PATH_DECODE_RF_U558 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5600, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_18_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5601, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5593);
   DLX_INST_DATA_PATH_DECODE_RF_U557 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4594, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4336, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5599);
   DLX_INST_DATA_PATH_DECODE_RF_U556 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7037, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7069, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5599, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5594);
   DLX_INST_DATA_PATH_DECODE_RF_U555 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4658, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4400, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5598);
   DLX_INST_DATA_PATH_DECODE_RF_U554 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6909, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6973, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5598, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5595);
   DLX_INST_DATA_PATH_DECODE_RF_U553 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4530, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4272, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5597);
   DLX_INST_DATA_PATH_DECODE_RF_U552 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7005, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6941, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5597, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5596);
   DLX_INST_DATA_PATH_DECODE_RF_U551 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5593, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5594, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5595, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5596, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4149);
   DLX_INST_DATA_PATH_DECODE_RF_U550 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4561, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4303, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5592);
   DLX_INST_DATA_PATH_DECODE_RF_U549 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6748, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6844, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5592, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5585);
   DLX_INST_DATA_PATH_DECODE_RF_U548 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4689, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4207, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4463, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5591);
   DLX_INST_DATA_PATH_DECODE_RF_U547 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6716, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6812, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5591, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5586);
   DLX_INST_DATA_PATH_DECODE_RF_U546 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4497, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4239, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5590);
   DLX_INST_DATA_PATH_DECODE_RF_U545 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6780, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6684, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5590, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5587);
   DLX_INST_DATA_PATH_DECODE_RF_U544 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4721, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4175, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4431, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5589);
   DLX_INST_DATA_PATH_DECODE_RF_U543 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6876, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6652, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5589, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5588);
   DLX_INST_DATA_PATH_DECODE_RF_U542 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5585, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5586, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5587, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5588, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5583);
   DLX_INST_DATA_PATH_DECODE_RF_U541 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4625, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4367, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5584);
   DLX_INST_DATA_PATH_DECODE_RF_U540 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5583, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_19_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5584, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5576);
   DLX_INST_DATA_PATH_DECODE_RF_U539 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4593, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4335, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5582);
   DLX_INST_DATA_PATH_DECODE_RF_U538 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7036, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7068, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5582, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5577);
   DLX_INST_DATA_PATH_DECODE_RF_U537 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4657, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4399, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5581);
   DLX_INST_DATA_PATH_DECODE_RF_U536 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6908, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6972, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5581, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5578);
   DLX_INST_DATA_PATH_DECODE_RF_U535 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4529, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4271, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5580);
   DLX_INST_DATA_PATH_DECODE_RF_U534 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7004, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6940, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5580, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5579);
   DLX_INST_DATA_PATH_DECODE_RF_U533 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5576, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5577, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5578, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5579, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4150);
   DLX_INST_DATA_PATH_DECODE_RF_U532 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4560, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4302, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5575);
   DLX_INST_DATA_PATH_DECODE_RF_U531 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6747, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6843, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5575, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5568);
   DLX_INST_DATA_PATH_DECODE_RF_U530 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4688, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4206, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4462, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5574);
   DLX_INST_DATA_PATH_DECODE_RF_U529 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6715, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6811, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5574, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5569);
   DLX_INST_DATA_PATH_DECODE_RF_U528 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4496, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4238, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5573);
   DLX_INST_DATA_PATH_DECODE_RF_U527 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6779, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6683, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5573, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5570);
   DLX_INST_DATA_PATH_DECODE_RF_U526 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4720, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4174, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4430, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5572);
   DLX_INST_DATA_PATH_DECODE_RF_U525 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6875, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6651, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5572, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5571);
   DLX_INST_DATA_PATH_DECODE_RF_U524 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5568, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5569, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5570, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5571, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5566);
   DLX_INST_DATA_PATH_DECODE_RF_U523 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4624, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4366, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5567);
   DLX_INST_DATA_PATH_DECODE_RF_U522 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5566, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_20_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5567, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5559);
   DLX_INST_DATA_PATH_DECODE_RF_U521 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4592, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4334, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5565);
   DLX_INST_DATA_PATH_DECODE_RF_U520 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7035, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7067, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5565, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5560);
   DLX_INST_DATA_PATH_DECODE_RF_U519 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4656, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4398, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5564);
   DLX_INST_DATA_PATH_DECODE_RF_U518 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6907, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6971, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5564, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5561);
   DLX_INST_DATA_PATH_DECODE_RF_U517 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4528, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4270, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5563);
   DLX_INST_DATA_PATH_DECODE_RF_U516 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7003, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6939, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5563, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5562);
   DLX_INST_DATA_PATH_DECODE_RF_U515 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5559, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5560, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5561, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5562, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4151);
   DLX_INST_DATA_PATH_DECODE_RF_U514 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4559, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4301, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5558);
   DLX_INST_DATA_PATH_DECODE_RF_U513 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6746, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6842, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5558, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5551);
   DLX_INST_DATA_PATH_DECODE_RF_U512 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4687, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4205, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4461, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5557);
   DLX_INST_DATA_PATH_DECODE_RF_U511 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6714, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6810, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5557, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5552);
   DLX_INST_DATA_PATH_DECODE_RF_U510 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4495, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4237, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5556);
   DLX_INST_DATA_PATH_DECODE_RF_U509 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6778, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6682, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5556, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5553);
   DLX_INST_DATA_PATH_DECODE_RF_U508 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4719, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4173, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4429, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5555);
   DLX_INST_DATA_PATH_DECODE_RF_U507 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6874, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6650, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5555, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5554);
   DLX_INST_DATA_PATH_DECODE_RF_U506 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5551, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5552, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5553, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5554, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5549);
   DLX_INST_DATA_PATH_DECODE_RF_U505 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4623, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4365, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5550);
   DLX_INST_DATA_PATH_DECODE_RF_U504 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5549, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_21_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5550, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5542);
   DLX_INST_DATA_PATH_DECODE_RF_U503 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4591, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4333, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5548);
   DLX_INST_DATA_PATH_DECODE_RF_U502 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7034, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7066, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5548, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5543);
   DLX_INST_DATA_PATH_DECODE_RF_U501 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4655, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4397, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5547);
   DLX_INST_DATA_PATH_DECODE_RF_U500 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6906, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6970, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5547, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5544);
   DLX_INST_DATA_PATH_DECODE_RF_U499 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4527, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4269, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5546);
   DLX_INST_DATA_PATH_DECODE_RF_U498 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7002, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6938, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5546, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5545);
   DLX_INST_DATA_PATH_DECODE_RF_U497 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5542, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5543, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5544, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5545, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4152);
   DLX_INST_DATA_PATH_DECODE_RF_U496 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4558, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4300, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5541);
   DLX_INST_DATA_PATH_DECODE_RF_U495 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6745, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6841, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5541, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5534);
   DLX_INST_DATA_PATH_DECODE_RF_U494 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4686, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4204, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4460, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5540);
   DLX_INST_DATA_PATH_DECODE_RF_U493 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6713, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6809, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5540, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5535);
   DLX_INST_DATA_PATH_DECODE_RF_U492 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4494, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4236, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5539);
   DLX_INST_DATA_PATH_DECODE_RF_U491 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6777, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6681, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5539, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5536);
   DLX_INST_DATA_PATH_DECODE_RF_U490 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4718, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4172, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4428, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5538);
   DLX_INST_DATA_PATH_DECODE_RF_U489 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6873, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6649, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5538, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5537);
   DLX_INST_DATA_PATH_DECODE_RF_U488 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5534, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5535, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5536, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5537, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5532);
   DLX_INST_DATA_PATH_DECODE_RF_U487 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4622, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4364, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5533);
   DLX_INST_DATA_PATH_DECODE_RF_U486 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5532, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_22_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5533, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5525);
   DLX_INST_DATA_PATH_DECODE_RF_U485 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4590, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4332, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5531);
   DLX_INST_DATA_PATH_DECODE_RF_U484 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7033, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7065, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5531, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5526);
   DLX_INST_DATA_PATH_DECODE_RF_U483 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4654, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4396, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5530);
   DLX_INST_DATA_PATH_DECODE_RF_U482 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6905, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6969, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5530, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5527);
   DLX_INST_DATA_PATH_DECODE_RF_U481 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4526, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4268, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5529);
   DLX_INST_DATA_PATH_DECODE_RF_U480 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7001, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6937, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5529, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5528);
   DLX_INST_DATA_PATH_DECODE_RF_U479 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5525, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5526, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5527, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5528, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4153);
   DLX_INST_DATA_PATH_DECODE_RF_U478 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4557, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4299, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5524);
   DLX_INST_DATA_PATH_DECODE_RF_U477 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6744, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6840, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5524, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5517);
   DLX_INST_DATA_PATH_DECODE_RF_U476 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4685, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4203, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4459, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5523);
   DLX_INST_DATA_PATH_DECODE_RF_U475 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6712, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6808, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5523, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5518);
   DLX_INST_DATA_PATH_DECODE_RF_U474 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4493, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4235, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5522);
   DLX_INST_DATA_PATH_DECODE_RF_U473 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6776, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6680, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5522, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5519);
   DLX_INST_DATA_PATH_DECODE_RF_U472 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4717, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4171, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4427, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5521);
   DLX_INST_DATA_PATH_DECODE_RF_U471 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6872, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6648, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5521, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5520);
   DLX_INST_DATA_PATH_DECODE_RF_U470 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5517, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5518, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5519, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5520, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5515);
   DLX_INST_DATA_PATH_DECODE_RF_U469 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4621, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4363, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5516);
   DLX_INST_DATA_PATH_DECODE_RF_U468 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5515, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_23_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5516, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5508);
   DLX_INST_DATA_PATH_DECODE_RF_U467 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4589, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4331, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5514);
   DLX_INST_DATA_PATH_DECODE_RF_U466 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7032, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7064, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5514, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5509);
   DLX_INST_DATA_PATH_DECODE_RF_U465 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4653, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4395, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5513);
   DLX_INST_DATA_PATH_DECODE_RF_U464 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6904, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6968, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5513, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5510);
   DLX_INST_DATA_PATH_DECODE_RF_U463 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4525, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4267, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5512);
   DLX_INST_DATA_PATH_DECODE_RF_U462 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7000, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6936, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5512, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5511);
   DLX_INST_DATA_PATH_DECODE_RF_U461 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5508, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5509, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5510, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5511, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4154);
   DLX_INST_DATA_PATH_DECODE_RF_U460 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4556, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4298, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5507);
   DLX_INST_DATA_PATH_DECODE_RF_U459 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6743, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6839, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5507, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5500);
   DLX_INST_DATA_PATH_DECODE_RF_U458 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4684, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4202, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4458, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5506);
   DLX_INST_DATA_PATH_DECODE_RF_U457 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6711, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6807, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5506, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5501);
   DLX_INST_DATA_PATH_DECODE_RF_U456 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4492, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4234, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5505);
   DLX_INST_DATA_PATH_DECODE_RF_U455 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6775, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6679, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5505, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5502);
   DLX_INST_DATA_PATH_DECODE_RF_U454 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4716, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4170, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4426, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5504);
   DLX_INST_DATA_PATH_DECODE_RF_U453 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6871, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6647, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5504, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5503);
   DLX_INST_DATA_PATH_DECODE_RF_U452 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5500, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5501, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5502, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5503, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5498);
   DLX_INST_DATA_PATH_DECODE_RF_U451 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4620, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4362, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5499);
   DLX_INST_DATA_PATH_DECODE_RF_U450 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5498, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_24_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5499, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5491);
   DLX_INST_DATA_PATH_DECODE_RF_U449 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4588, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4330, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5497);
   DLX_INST_DATA_PATH_DECODE_RF_U448 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7031, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7063, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5497, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5492);
   DLX_INST_DATA_PATH_DECODE_RF_U447 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4652, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4394, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5496);
   DLX_INST_DATA_PATH_DECODE_RF_U446 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6903, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6967, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5496, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5493);
   DLX_INST_DATA_PATH_DECODE_RF_U445 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4524, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4266, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5495);
   DLX_INST_DATA_PATH_DECODE_RF_U444 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6999, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6935, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5495, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5494);
   DLX_INST_DATA_PATH_DECODE_RF_U443 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5491, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5492, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5493, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5494, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4155);
   DLX_INST_DATA_PATH_DECODE_RF_U442 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4555, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4297, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5490);
   DLX_INST_DATA_PATH_DECODE_RF_U441 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6742, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6838, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5490, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5483);
   DLX_INST_DATA_PATH_DECODE_RF_U440 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4683, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4201, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4457, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5489);
   DLX_INST_DATA_PATH_DECODE_RF_U439 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6710, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6806, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5489, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5484);
   DLX_INST_DATA_PATH_DECODE_RF_U438 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4491, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4233, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5488);
   DLX_INST_DATA_PATH_DECODE_RF_U437 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6774, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6678, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5488, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5485);
   DLX_INST_DATA_PATH_DECODE_RF_U436 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4715, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4169, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4425, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5487);
   DLX_INST_DATA_PATH_DECODE_RF_U435 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6870, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6646, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5487, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5486);
   DLX_INST_DATA_PATH_DECODE_RF_U434 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5483, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5484, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5485, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5486, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5481);
   DLX_INST_DATA_PATH_DECODE_RF_U433 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4619, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4361, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5482);
   DLX_INST_DATA_PATH_DECODE_RF_U432 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5481, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_25_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5482, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5474);
   DLX_INST_DATA_PATH_DECODE_RF_U431 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4587, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4329, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5480);
   DLX_INST_DATA_PATH_DECODE_RF_U430 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7030, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7062, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5480, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5475);
   DLX_INST_DATA_PATH_DECODE_RF_U429 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4651, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4393, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5479);
   DLX_INST_DATA_PATH_DECODE_RF_U428 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6902, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6966, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5479, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5476);
   DLX_INST_DATA_PATH_DECODE_RF_U427 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4523, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4265, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5478);
   DLX_INST_DATA_PATH_DECODE_RF_U426 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6998, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6934, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5478, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5477);
   DLX_INST_DATA_PATH_DECODE_RF_U425 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5474, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5475, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5476, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5477, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4156);
   DLX_INST_DATA_PATH_DECODE_RF_U424 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4554, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4296, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5473);
   DLX_INST_DATA_PATH_DECODE_RF_U423 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6741, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6837, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5473, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5466);
   DLX_INST_DATA_PATH_DECODE_RF_U422 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4682, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4200, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4456, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5472);
   DLX_INST_DATA_PATH_DECODE_RF_U421 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6709, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6805, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5472, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5467);
   DLX_INST_DATA_PATH_DECODE_RF_U420 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4490, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4232, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5471);
   DLX_INST_DATA_PATH_DECODE_RF_U419 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6773, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6677, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5471, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5468);
   DLX_INST_DATA_PATH_DECODE_RF_U418 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4714, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4168, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4424, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5470);
   DLX_INST_DATA_PATH_DECODE_RF_U417 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6869, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6645, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5470, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5469);
   DLX_INST_DATA_PATH_DECODE_RF_U416 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5466, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5467, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5468, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5469, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5464);
   DLX_INST_DATA_PATH_DECODE_RF_U415 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4618, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4360, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5465);
   DLX_INST_DATA_PATH_DECODE_RF_U414 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5464, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_26_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5465, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5457);
   DLX_INST_DATA_PATH_DECODE_RF_U413 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4586, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4328, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5463);
   DLX_INST_DATA_PATH_DECODE_RF_U412 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7029, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7061, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5463, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5458);
   DLX_INST_DATA_PATH_DECODE_RF_U411 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4650, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4392, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5462);
   DLX_INST_DATA_PATH_DECODE_RF_U410 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6901, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6965, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5462, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5459);
   DLX_INST_DATA_PATH_DECODE_RF_U409 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4522, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4264, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5461);
   DLX_INST_DATA_PATH_DECODE_RF_U408 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6997, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6933, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5461, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5460);
   DLX_INST_DATA_PATH_DECODE_RF_U407 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5457, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5458, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5459, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5460, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4157);
   DLX_INST_DATA_PATH_DECODE_RF_U406 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4553, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4295, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5456);
   DLX_INST_DATA_PATH_DECODE_RF_U405 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6740, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6836, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5456, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5449);
   DLX_INST_DATA_PATH_DECODE_RF_U404 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4681, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4199, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4455, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5455);
   DLX_INST_DATA_PATH_DECODE_RF_U403 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6708, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6804, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5455, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5450);
   DLX_INST_DATA_PATH_DECODE_RF_U402 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4489, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4231, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5454);
   DLX_INST_DATA_PATH_DECODE_RF_U401 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6772, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6676, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5454, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5451);
   DLX_INST_DATA_PATH_DECODE_RF_U400 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4713, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4167, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4423, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5453);
   DLX_INST_DATA_PATH_DECODE_RF_U399 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6868, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6644, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5453, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5452);
   DLX_INST_DATA_PATH_DECODE_RF_U398 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5449, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5450, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5451, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5452, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5447);
   DLX_INST_DATA_PATH_DECODE_RF_U397 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4617, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4359, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5448);
   DLX_INST_DATA_PATH_DECODE_RF_U396 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5447, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_27_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5448, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5440);
   DLX_INST_DATA_PATH_DECODE_RF_U395 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4585, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4327, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5446);
   DLX_INST_DATA_PATH_DECODE_RF_U394 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7028, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7060, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5446, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5441);
   DLX_INST_DATA_PATH_DECODE_RF_U393 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4649, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4391, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5445);
   DLX_INST_DATA_PATH_DECODE_RF_U392 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6900, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6964, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5445, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5442);
   DLX_INST_DATA_PATH_DECODE_RF_U391 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4521, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4263, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5444);
   DLX_INST_DATA_PATH_DECODE_RF_U390 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6996, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6932, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5444, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5443);
   DLX_INST_DATA_PATH_DECODE_RF_U389 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5440, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5441, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5442, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5443, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4158);
   DLX_INST_DATA_PATH_DECODE_RF_U388 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4552, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4294, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5439);
   DLX_INST_DATA_PATH_DECODE_RF_U387 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6739, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6835, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5439, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5432);
   DLX_INST_DATA_PATH_DECODE_RF_U386 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4680, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4198, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4454, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5438);
   DLX_INST_DATA_PATH_DECODE_RF_U385 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6707, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6803, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5438, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5433);
   DLX_INST_DATA_PATH_DECODE_RF_U384 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4488, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4230, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5437);
   DLX_INST_DATA_PATH_DECODE_RF_U383 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6771, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6675, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5437, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5434);
   DLX_INST_DATA_PATH_DECODE_RF_U382 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4712, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4166, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4422, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5436);
   DLX_INST_DATA_PATH_DECODE_RF_U381 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6867, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6643, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5436, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5435);
   DLX_INST_DATA_PATH_DECODE_RF_U380 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5432, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5433, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5434, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5435, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5430);
   DLX_INST_DATA_PATH_DECODE_RF_U379 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4616, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4358, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5431);
   DLX_INST_DATA_PATH_DECODE_RF_U378 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5430, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_28_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5431, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5423);
   DLX_INST_DATA_PATH_DECODE_RF_U377 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4584, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4326, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5429);
   DLX_INST_DATA_PATH_DECODE_RF_U376 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7027, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7059, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5429, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5424);
   DLX_INST_DATA_PATH_DECODE_RF_U375 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4648, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4390, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5428);
   DLX_INST_DATA_PATH_DECODE_RF_U374 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6899, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6963, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5428, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5425);
   DLX_INST_DATA_PATH_DECODE_RF_U373 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4520, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4262, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5427);
   DLX_INST_DATA_PATH_DECODE_RF_U372 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6995, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6931, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5427, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5426);
   DLX_INST_DATA_PATH_DECODE_RF_U371 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5423, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5424, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5425, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5426, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4159);
   DLX_INST_DATA_PATH_DECODE_RF_U370 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4551, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4293, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5422);
   DLX_INST_DATA_PATH_DECODE_RF_U369 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6738, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6834, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5422, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5415);
   DLX_INST_DATA_PATH_DECODE_RF_U368 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4679, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4197, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4453, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5421);
   DLX_INST_DATA_PATH_DECODE_RF_U367 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6706, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6802, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5421, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5416);
   DLX_INST_DATA_PATH_DECODE_RF_U366 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4487, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4229, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5420);
   DLX_INST_DATA_PATH_DECODE_RF_U365 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6770, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6674, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5420, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5417);
   DLX_INST_DATA_PATH_DECODE_RF_U364 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4711, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4165, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4421, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5419);
   DLX_INST_DATA_PATH_DECODE_RF_U363 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6866, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6642, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5419, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5418);
   DLX_INST_DATA_PATH_DECODE_RF_U362 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5415, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5416, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5417, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5418, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5413);
   DLX_INST_DATA_PATH_DECODE_RF_U361 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4615, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4357, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5414);
   DLX_INST_DATA_PATH_DECODE_RF_U360 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5413, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_29_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5414, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5406);
   DLX_INST_DATA_PATH_DECODE_RF_U359 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4583, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4325, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5412);
   DLX_INST_DATA_PATH_DECODE_RF_U358 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7026, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7058, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5412, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5407);
   DLX_INST_DATA_PATH_DECODE_RF_U357 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4647, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4389, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5411);
   DLX_INST_DATA_PATH_DECODE_RF_U356 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6898, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6962, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5411, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5408);
   DLX_INST_DATA_PATH_DECODE_RF_U355 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4519, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4261, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5410);
   DLX_INST_DATA_PATH_DECODE_RF_U354 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6994, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6930, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5410, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5409);
   DLX_INST_DATA_PATH_DECODE_RF_U353 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5406, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5407, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5408, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5409, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4160);
   DLX_INST_DATA_PATH_DECODE_RF_U352 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4550, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4292, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5405);
   DLX_INST_DATA_PATH_DECODE_RF_U351 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6737, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6833, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5405, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5398);
   DLX_INST_DATA_PATH_DECODE_RF_U350 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4678, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4196, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4452, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5404);
   DLX_INST_DATA_PATH_DECODE_RF_U349 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6705, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6801, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5404, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5399);
   DLX_INST_DATA_PATH_DECODE_RF_U348 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4486, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4228, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5403);
   DLX_INST_DATA_PATH_DECODE_RF_U347 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6769, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6673, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5403, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5400);
   DLX_INST_DATA_PATH_DECODE_RF_U346 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4710, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4164, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4420, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5402);
   DLX_INST_DATA_PATH_DECODE_RF_U345 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6865, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6641, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5402, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5401);
   DLX_INST_DATA_PATH_DECODE_RF_U344 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5398, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5399, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5400, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5401, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5396);
   DLX_INST_DATA_PATH_DECODE_RF_U343 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4614, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4356, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5397);
   DLX_INST_DATA_PATH_DECODE_RF_U342 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5396, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_30_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5397, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5389);
   DLX_INST_DATA_PATH_DECODE_RF_U341 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4582, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4324, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5395);
   DLX_INST_DATA_PATH_DECODE_RF_U340 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7025, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7057, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5395, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5390);
   DLX_INST_DATA_PATH_DECODE_RF_U339 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4646, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4388, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5394);
   DLX_INST_DATA_PATH_DECODE_RF_U338 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6897, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6961, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5394, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5391);
   DLX_INST_DATA_PATH_DECODE_RF_U337 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4518, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4260, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5393);
   DLX_INST_DATA_PATH_DECODE_RF_U336 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6993, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6929, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5393, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5392);
   DLX_INST_DATA_PATH_DECODE_RF_U335 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5389, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5390, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5391, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5392, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4161);
   DLX_INST_DATA_PATH_DECODE_RF_U334 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4549, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4291, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5386);
   DLX_INST_DATA_PATH_DECODE_RF_U333 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6736, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6832, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5386, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5363);
   DLX_INST_DATA_PATH_DECODE_RF_U332 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4677, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4195, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4451, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5380);
   DLX_INST_DATA_PATH_DECODE_RF_U331 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6704, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6800, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5380, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5364);
   DLX_INST_DATA_PATH_DECODE_RF_U330 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4485, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4227, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5375);
   DLX_INST_DATA_PATH_DECODE_RF_U329 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6768, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6672, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5375, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5365);
   DLX_INST_DATA_PATH_DECODE_RF_U328 : OAI222_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4709, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4163, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4419, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5369);
   DLX_INST_DATA_PATH_DECODE_RF_U327 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6864, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6640, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5369, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5366);
   DLX_INST_DATA_PATH_DECODE_RF_U326 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5363, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5364, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5365, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5366, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5359);
   DLX_INST_DATA_PATH_DECODE_RF_U325 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4613, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4355, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5360);
   DLX_INST_DATA_PATH_DECODE_RF_U324 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5359, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189, C2 => 
                           DLX_INST_DATA_PATH_A_outs_31_port, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5360, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5339);
   DLX_INST_DATA_PATH_DECODE_RF_U323 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4581, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4323, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5355);
   DLX_INST_DATA_PATH_DECODE_RF_U322 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7024, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7056, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5355, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5340);
   DLX_INST_DATA_PATH_DECODE_RF_U321 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4645, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4387, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5350);
   DLX_INST_DATA_PATH_DECODE_RF_U320 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6896, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6960, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5350, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5341);
   DLX_INST_DATA_PATH_DECODE_RF_U319 : OAI22_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4517, B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4259, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5345);
   DLX_INST_DATA_PATH_DECODE_RF_U318 : AOI221_X1 port map( B1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6992, B2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343, C1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6928, C2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344, A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5345, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5342);
   DLX_INST_DATA_PATH_DECODE_RF_U317 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5339, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5340, A3 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5341, A4 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5342, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4162);
   DLX_INST_DATA_PATH_DECODE_RF_U316 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n10, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5191);
   DLX_INST_DATA_PATH_DECODE_RF_U315 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5338, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5337);
   DLX_INST_DATA_PATH_DECODE_RF_U314 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5191, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5195);
   DLX_INST_DATA_PATH_DECODE_RF_U313 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5335, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5334);
   DLX_INST_DATA_PATH_DECODE_RF_U312 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5328, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5327);
   DLX_INST_DATA_PATH_DECODE_RF_U311 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5328, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5326);
   DLX_INST_DATA_PATH_DECODE_RF_U310 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5328, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5325);
   DLX_INST_DATA_PATH_DECODE_RF_U309 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5328, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5324);
   DLX_INST_DATA_PATH_DECODE_RF_U308 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5328, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5323);
   DLX_INST_DATA_PATH_DECODE_RF_U307 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5194, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193);
   DLX_INST_DATA_PATH_DECODE_RF_U306 : INV_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5194, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192);
   DLX_INST_DATA_PATH_DECODE_RF_U305 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5327, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196);
   DLX_INST_DATA_PATH_DECODE_RF_U304 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5327, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197);
   DLX_INST_DATA_PATH_DECODE_RF_U303 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5327, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198);
   DLX_INST_DATA_PATH_DECODE_RF_U302 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5326, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199);
   DLX_INST_DATA_PATH_DECODE_RF_U301 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5326, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200);
   DLX_INST_DATA_PATH_DECODE_RF_U300 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5326, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201);
   DLX_INST_DATA_PATH_DECODE_RF_U299 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5325, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202);
   DLX_INST_DATA_PATH_DECODE_RF_U298 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5325, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203);
   DLX_INST_DATA_PATH_DECODE_RF_U297 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5325, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204);
   DLX_INST_DATA_PATH_DECODE_RF_U296 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5324, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205);
   DLX_INST_DATA_PATH_DECODE_RF_U295 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5324, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206);
   DLX_INST_DATA_PATH_DECODE_RF_U294 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5324, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207);
   DLX_INST_DATA_PATH_DECODE_RF_U293 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5323, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208);
   DLX_INST_DATA_PATH_DECODE_RF_U292 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5323, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209);
   DLX_INST_DATA_PATH_DECODE_RF_U291 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5323, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210);
   DLX_INST_DATA_PATH_DECODE_RF_U290 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5334, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5295);
   DLX_INST_DATA_PATH_DECODE_RF_U289 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5334, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5297);
   DLX_INST_DATA_PATH_DECODE_RF_U288 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5334, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5296);
   DLX_INST_DATA_PATH_DECODE_RF_U287 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5333, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5298);
   DLX_INST_DATA_PATH_DECODE_RF_U286 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5329, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5322);
   DLX_INST_DATA_PATH_DECODE_RF_U285 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5329, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5321);
   DLX_INST_DATA_PATH_DECODE_RF_U284 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5333, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5302);
   DLX_INST_DATA_PATH_DECODE_RF_U283 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5333, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5301);
   DLX_INST_DATA_PATH_DECODE_RF_U282 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5329, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5318);
   DLX_INST_DATA_PATH_DECODE_RF_U281 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5330, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5317);
   DLX_INST_DATA_PATH_DECODE_RF_U280 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5330, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5314);
   DLX_INST_DATA_PATH_DECODE_RF_U279 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5330, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5313);
   DLX_INST_DATA_PATH_DECODE_RF_U278 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5332, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5306);
   DLX_INST_DATA_PATH_DECODE_RF_U277 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5332, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5305);
   DLX_INST_DATA_PATH_DECODE_RF_U276 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5331, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5310);
   DLX_INST_DATA_PATH_DECODE_RF_U275 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5331, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5309);
   DLX_INST_DATA_PATH_DECODE_RF_U274 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5329, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5320);
   DLX_INST_DATA_PATH_DECODE_RF_U273 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5333, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5300);
   DLX_INST_DATA_PATH_DECODE_RF_U272 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5330, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5316);
   DLX_INST_DATA_PATH_DECODE_RF_U271 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5331, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5312);
   DLX_INST_DATA_PATH_DECODE_RF_U270 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5332, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5304);
   DLX_INST_DATA_PATH_DECODE_RF_U269 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5331, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5308);
   DLX_INST_DATA_PATH_DECODE_RF_U268 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5329, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5319);
   DLX_INST_DATA_PATH_DECODE_RF_U267 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5333, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5299);
   DLX_INST_DATA_PATH_DECODE_RF_U266 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5330, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5315);
   DLX_INST_DATA_PATH_DECODE_RF_U265 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5331, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5311);
   DLX_INST_DATA_PATH_DECODE_RF_U264 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5332, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5303);
   DLX_INST_DATA_PATH_DECODE_RF_U263 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5332, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5307);
   DLX_INST_DATA_PATH_DECODE_RF_U262 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5295, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5294);
   DLX_INST_DATA_PATH_DECODE_RF_U261 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5298, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283);
   DLX_INST_DATA_PATH_DECODE_RF_U260 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5298, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284);
   DLX_INST_DATA_PATH_DECODE_RF_U259 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5298, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285);
   DLX_INST_DATA_PATH_DECODE_RF_U258 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5322, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213);
   DLX_INST_DATA_PATH_DECODE_RF_U257 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5321, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214);
   DLX_INST_DATA_PATH_DECODE_RF_U256 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5321, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215);
   DLX_INST_DATA_PATH_DECODE_RF_U255 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5321, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216);
   DLX_INST_DATA_PATH_DECODE_RF_U254 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5302, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271);
   DLX_INST_DATA_PATH_DECODE_RF_U253 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5302, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272);
   DLX_INST_DATA_PATH_DECODE_RF_U252 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5302, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273);
   DLX_INST_DATA_PATH_DECODE_RF_U251 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5301, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274);
   DLX_INST_DATA_PATH_DECODE_RF_U250 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5318, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225);
   DLX_INST_DATA_PATH_DECODE_RF_U249 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5317, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226);
   DLX_INST_DATA_PATH_DECODE_RF_U248 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5317, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227);
   DLX_INST_DATA_PATH_DECODE_RF_U247 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5314, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236);
   DLX_INST_DATA_PATH_DECODE_RF_U246 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5314, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237);
   DLX_INST_DATA_PATH_DECODE_RF_U245 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5313, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238);
   DLX_INST_DATA_PATH_DECODE_RF_U244 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5313, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239);
   DLX_INST_DATA_PATH_DECODE_RF_U243 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5306, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259);
   DLX_INST_DATA_PATH_DECODE_RF_U242 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5306, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260);
   DLX_INST_DATA_PATH_DECODE_RF_U241 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5306, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261);
   DLX_INST_DATA_PATH_DECODE_RF_U240 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5305, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262);
   DLX_INST_DATA_PATH_DECODE_RF_U239 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5310, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248);
   DLX_INST_DATA_PATH_DECODE_RF_U238 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5310, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249);
   DLX_INST_DATA_PATH_DECODE_RF_U237 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5309, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250);
   DLX_INST_DATA_PATH_DECODE_RF_U236 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5309, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251);
   DLX_INST_DATA_PATH_DECODE_RF_U235 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5297, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286);
   DLX_INST_DATA_PATH_DECODE_RF_U234 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5297, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287);
   DLX_INST_DATA_PATH_DECODE_RF_U233 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5297, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288);
   DLX_INST_DATA_PATH_DECODE_RF_U232 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5320, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217);
   DLX_INST_DATA_PATH_DECODE_RF_U231 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5320, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218);
   DLX_INST_DATA_PATH_DECODE_RF_U230 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5320, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219);
   DLX_INST_DATA_PATH_DECODE_RF_U229 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5301, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275);
   DLX_INST_DATA_PATH_DECODE_RF_U228 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5301, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276);
   DLX_INST_DATA_PATH_DECODE_RF_U227 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5300, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277);
   DLX_INST_DATA_PATH_DECODE_RF_U226 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5317, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228);
   DLX_INST_DATA_PATH_DECODE_RF_U225 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5316, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229);
   DLX_INST_DATA_PATH_DECODE_RF_U224 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5316, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230);
   DLX_INST_DATA_PATH_DECODE_RF_U223 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5313, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240);
   DLX_INST_DATA_PATH_DECODE_RF_U222 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5312, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241);
   DLX_INST_DATA_PATH_DECODE_RF_U221 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5312, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242);
   DLX_INST_DATA_PATH_DECODE_RF_U220 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5305, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263);
   DLX_INST_DATA_PATH_DECODE_RF_U219 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5305, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264);
   DLX_INST_DATA_PATH_DECODE_RF_U218 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5304, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265);
   DLX_INST_DATA_PATH_DECODE_RF_U217 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5309, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252);
   DLX_INST_DATA_PATH_DECODE_RF_U216 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5308, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253);
   DLX_INST_DATA_PATH_DECODE_RF_U215 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5308, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254);
   DLX_INST_DATA_PATH_DECODE_RF_U214 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5296, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289);
   DLX_INST_DATA_PATH_DECODE_RF_U213 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5296, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290);
   DLX_INST_DATA_PATH_DECODE_RF_U212 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5296, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291);
   DLX_INST_DATA_PATH_DECODE_RF_U211 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5319, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220);
   DLX_INST_DATA_PATH_DECODE_RF_U210 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5319, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221);
   DLX_INST_DATA_PATH_DECODE_RF_U209 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5319, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222);
   DLX_INST_DATA_PATH_DECODE_RF_U208 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5300, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278);
   DLX_INST_DATA_PATH_DECODE_RF_U207 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5300, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279);
   DLX_INST_DATA_PATH_DECODE_RF_U206 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5299, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280);
   DLX_INST_DATA_PATH_DECODE_RF_U205 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5316, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231);
   DLX_INST_DATA_PATH_DECODE_RF_U204 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5315, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232);
   DLX_INST_DATA_PATH_DECODE_RF_U203 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5315, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233);
   DLX_INST_DATA_PATH_DECODE_RF_U202 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5312, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243);
   DLX_INST_DATA_PATH_DECODE_RF_U201 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5311, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244);
   DLX_INST_DATA_PATH_DECODE_RF_U200 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5311, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245);
   DLX_INST_DATA_PATH_DECODE_RF_U199 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5304, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266);
   DLX_INST_DATA_PATH_DECODE_RF_U198 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5304, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267);
   DLX_INST_DATA_PATH_DECODE_RF_U197 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5303, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268);
   DLX_INST_DATA_PATH_DECODE_RF_U196 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5308, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255);
   DLX_INST_DATA_PATH_DECODE_RF_U195 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5307, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256);
   DLX_INST_DATA_PATH_DECODE_RF_U194 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5295, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292);
   DLX_INST_DATA_PATH_DECODE_RF_U193 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5295, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293);
   DLX_INST_DATA_PATH_DECODE_RF_U192 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5318, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223);
   DLX_INST_DATA_PATH_DECODE_RF_U191 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5318, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224);
   DLX_INST_DATA_PATH_DECODE_RF_U190 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5299, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281);
   DLX_INST_DATA_PATH_DECODE_RF_U189 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5299, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282);
   DLX_INST_DATA_PATH_DECODE_RF_U188 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5315, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234);
   DLX_INST_DATA_PATH_DECODE_RF_U187 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5314, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235);
   DLX_INST_DATA_PATH_DECODE_RF_U186 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5311, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246);
   DLX_INST_DATA_PATH_DECODE_RF_U185 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5310, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247);
   DLX_INST_DATA_PATH_DECODE_RF_U184 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5303, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269);
   DLX_INST_DATA_PATH_DECODE_RF_U183 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5303, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270);
   DLX_INST_DATA_PATH_DECODE_RF_U182 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5307, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257);
   DLX_INST_DATA_PATH_DECODE_RF_U181 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5307, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258);
   DLX_INST_DATA_PATH_DECODE_RF_U180 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5322, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211);
   DLX_INST_DATA_PATH_DECODE_RF_U179 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5322, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212);
   DLX_INST_DATA_PATH_DECODE_RF_U178 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_n11, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5338);
   DLX_INST_DATA_PATH_DECODE_RF_U177 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5338, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5335);
   DLX_INST_DATA_PATH_DECODE_RF_U176 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5338, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5336);
   DLX_INST_DATA_PATH_DECODE_RF_U175 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5337, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5328);
   DLX_INST_DATA_PATH_DECODE_RF_U174 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5191, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5194);
   DLX_INST_DATA_PATH_DECODE_RF_U173 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5335, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5333);
   DLX_INST_DATA_PATH_DECODE_RF_U172 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5336, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5329);
   DLX_INST_DATA_PATH_DECODE_RF_U171 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5336, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5330);
   DLX_INST_DATA_PATH_DECODE_RF_U170 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5335, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5332);
   DLX_INST_DATA_PATH_DECODE_RF_U169 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5336, Z => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5331);
   DLX_INST_DATA_PATH_DECODE_RF_U168 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358);
   DLX_INST_DATA_PATH_DECODE_RF_U167 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, A2 => 
                           DLX_INST_DATA_PATH_DECODE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952);
   DLX_INST_DATA_PATH_DECODE_RF_U166 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6561, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6562, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527);
   DLX_INST_DATA_PATH_DECODE_RF_U165 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6623, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6580, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636);
   DLX_INST_DATA_PATH_DECODE_RF_U164 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6606, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6571, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611);
   DLX_INST_DATA_PATH_DECODE_RF_U163 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6589, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6583, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602);
   DLX_INST_DATA_PATH_DECODE_RF_U162 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5924, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5907, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5376);
   DLX_INST_DATA_PATH_DECODE_RF_U161 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5912, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5915, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5387);
   DLX_INST_DATA_PATH_DECODE_RF_U160 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5906, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5905, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5346);
   DLX_INST_DATA_PATH_DECODE_RF_U159 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5911, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5904, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5361);
   DLX_INST_DATA_PATH_DECODE_RF_U158 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5925, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5914, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5379);
   DLX_INST_DATA_PATH_DECODE_RF_U157 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_0_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6560);
   DLX_INST_DATA_PATH_DECODE_RF_U156 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_1_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6559);
   DLX_INST_DATA_PATH_DECODE_RF_U155 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_2_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6558);
   DLX_INST_DATA_PATH_DECODE_RF_U154 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_3_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6557);
   DLX_INST_DATA_PATH_DECODE_RF_U153 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_4_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6556);
   DLX_INST_DATA_PATH_DECODE_RF_U152 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_5_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6555);
   DLX_INST_DATA_PATH_DECODE_RF_U151 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_6_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6554);
   DLX_INST_DATA_PATH_DECODE_RF_U150 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_7_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6553);
   DLX_INST_DATA_PATH_DECODE_RF_U149 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_8_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6552);
   DLX_INST_DATA_PATH_DECODE_RF_U148 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_9_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6551);
   DLX_INST_DATA_PATH_DECODE_RF_U147 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_10_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6550);
   DLX_INST_DATA_PATH_DECODE_RF_U146 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_11_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6549);
   DLX_INST_DATA_PATH_DECODE_RF_U145 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_12_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6548);
   DLX_INST_DATA_PATH_DECODE_RF_U144 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_13_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6547);
   DLX_INST_DATA_PATH_DECODE_RF_U143 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_14_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6546);
   DLX_INST_DATA_PATH_DECODE_RF_U142 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_15_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6545);
   DLX_INST_DATA_PATH_DECODE_RF_U141 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_16_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6544);
   DLX_INST_DATA_PATH_DECODE_RF_U140 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_17_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6543);
   DLX_INST_DATA_PATH_DECODE_RF_U139 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_18_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6542);
   DLX_INST_DATA_PATH_DECODE_RF_U138 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_19_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6541);
   DLX_INST_DATA_PATH_DECODE_RF_U137 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_20_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6540);
   DLX_INST_DATA_PATH_DECODE_RF_U136 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_21_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6539);
   DLX_INST_DATA_PATH_DECODE_RF_U135 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_22_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6538);
   DLX_INST_DATA_PATH_DECODE_RF_U134 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_23_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6537);
   DLX_INST_DATA_PATH_DECODE_RF_U133 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_24_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6536);
   DLX_INST_DATA_PATH_DECODE_RF_U132 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_25_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6535);
   DLX_INST_DATA_PATH_DECODE_RF_U131 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_26_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6534);
   DLX_INST_DATA_PATH_DECODE_RF_U130 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_27_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6533);
   DLX_INST_DATA_PATH_DECODE_RF_U129 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_28_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6532);
   DLX_INST_DATA_PATH_DECODE_RF_U128 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_29_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6531);
   DLX_INST_DATA_PATH_DECODE_RF_U127 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_30_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6530);
   DLX_INST_DATA_PATH_DECODE_RF_U126 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_31_port, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6528);
   DLX_INST_DATA_PATH_DECODE_RF_U125 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6519, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6507, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5976);
   DLX_INST_DATA_PATH_DECODE_RF_U124 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6518, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6504, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5965);
   DLX_INST_DATA_PATH_DECODE_RF_U123 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6636, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6637);
   DLX_INST_DATA_PATH_DECODE_RF_U122 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6611, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6612);
   DLX_INST_DATA_PATH_DECODE_RF_U121 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6505, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6500, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5951);
   DLX_INST_DATA_PATH_DECODE_RF_U120 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6498, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6499, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5941);
   DLX_INST_DATA_PATH_DECODE_RF_U119 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6527, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6529);
   DLX_INST_DATA_PATH_DECODE_RF_U118 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6506, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6509, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5981);
   DLX_INST_DATA_PATH_DECODE_RF_U117 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6623, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6568, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627);
   DLX_INST_DATA_PATH_DECODE_RF_U116 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6606, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6580, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617);
   DLX_INST_DATA_PATH_DECODE_RF_U115 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6589, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6574, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596);
   DLX_INST_DATA_PATH_DECODE_RF_U114 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6571, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6562, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569);
   DLX_INST_DATA_PATH_DECODE_RF_U113 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5912, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5911, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5351);
   DLX_INST_DATA_PATH_DECODE_RF_U112 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5924, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5913, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5374);
   DLX_INST_DATA_PATH_DECODE_RF_U111 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5925, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5904, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5385);
   DLX_INST_DATA_PATH_DECODE_RF_U110 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5907, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5905, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5344);
   DLX_INST_DATA_PATH_DECODE_RF_U109 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5910, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5915, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5388);
   DLX_INST_DATA_PATH_DECODE_RF_U108 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6627, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6628);
   DLX_INST_DATA_PATH_DECODE_RF_U107 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6602, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6603);
   DLX_INST_DATA_PATH_DECODE_RF_U106 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6569, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6570);
   DLX_INST_DATA_PATH_DECODE_RF_U105 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6519, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6500, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5971);
   DLX_INST_DATA_PATH_DECODE_RF_U104 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6504, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6509, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5982);
   DLX_INST_DATA_PATH_DECODE_RF_U103 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6505, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6508, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5956);
   DLX_INST_DATA_PATH_DECODE_RF_U102 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6518, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6502, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5975);
   DLX_INST_DATA_PATH_DECODE_RF_U101 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6501, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6499, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5938);
   DLX_INST_DATA_PATH_DECODE_RF_U100 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6606, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6568, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609);
   DLX_INST_DATA_PATH_DECODE_RF_U99 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6589, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6571, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594);
   DLX_INST_DATA_PATH_DECODE_RF_U98 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6574, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6562, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572);
   DLX_INST_DATA_PATH_DECODE_RF_U97 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6623, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6583, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638);
   DLX_INST_DATA_PATH_DECODE_RF_U96 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5911, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5907, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5356);
   DLX_INST_DATA_PATH_DECODE_RF_U95 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5913, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5905, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5349);
   DLX_INST_DATA_PATH_DECODE_RF_U94 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5924, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5906, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5368);
   DLX_INST_DATA_PATH_DECODE_RF_U93 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6617, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6618);
   DLX_INST_DATA_PATH_DECODE_RF_U92 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6609, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6610);
   DLX_INST_DATA_PATH_DECODE_RF_U91 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6504, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6505, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5946);
   DLX_INST_DATA_PATH_DECODE_RF_U90 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5925, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5908, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5383);
   DLX_INST_DATA_PATH_DECODE_RF_U89 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6519, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6508, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5973);
   DLX_INST_DATA_PATH_DECODE_RF_U88 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6518, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6500, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5962);
   DLX_INST_DATA_PATH_DECODE_RF_U87 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6507, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6499, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5943);
   DLX_INST_DATA_PATH_DECODE_RF_U86 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6606, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6561, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604);
   DLX_INST_DATA_PATH_DECODE_RF_U85 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6568, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6562, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566);
   DLX_INST_DATA_PATH_DECODE_RF_U84 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6623, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6577, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634);
   DLX_INST_DATA_PATH_DECODE_RF_U83 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6589, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6580, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600);
   DLX_INST_DATA_PATH_DECODE_RF_U82 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5911, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5908, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5354);
   DLX_INST_DATA_PATH_DECODE_RF_U81 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5925, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5906, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5377);
   DLX_INST_DATA_PATH_DECODE_RF_U80 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5904, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5905, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5347);
   DLX_INST_DATA_PATH_DECODE_RF_U79 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5924, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5910, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5371);
   DLX_INST_DATA_PATH_DECODE_RF_U78 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6604, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6605);
   DLX_INST_DATA_PATH_DECODE_RF_U77 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6638, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6639);
   DLX_INST_DATA_PATH_DECODE_RF_U76 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6519, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6504, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5964);
   DLX_INST_DATA_PATH_DECODE_RF_U75 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6505, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6502, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5948);
   DLX_INST_DATA_PATH_DECODE_RF_U74 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6518, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6507, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5968);
   DLX_INST_DATA_PATH_DECODE_RF_U73 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6500, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6499, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5940);
   DLX_INST_DATA_PATH_DECODE_RF_U72 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6589, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6561, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587);
   DLX_INST_DATA_PATH_DECODE_RF_U71 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6565, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6562, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563);
   DLX_INST_DATA_PATH_DECODE_RF_U70 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6623, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6574, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632);
   DLX_INST_DATA_PATH_DECODE_RF_U69 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6606, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6583, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619);
   DLX_INST_DATA_PATH_DECODE_RF_U68 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5910, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5911, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5352);
   DLX_INST_DATA_PATH_DECODE_RF_U67 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5925, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5913, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5382);
   DLX_INST_DATA_PATH_DECODE_RF_U66 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6596, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6597);
   DLX_INST_DATA_PATH_DECODE_RF_U65 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6634, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6635);
   DLX_INST_DATA_PATH_DECODE_RF_U64 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5924, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5912, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5372);
   DLX_INST_DATA_PATH_DECODE_RF_U63 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6519, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6498, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5979);
   DLX_INST_DATA_PATH_DECODE_RF_U62 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5914, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5905, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5348);
   DLX_INST_DATA_PATH_DECODE_RF_U61 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6518, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6501, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5970);
   DLX_INST_DATA_PATH_DECODE_RF_U60 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6506, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6505, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5945);
   DLX_INST_DATA_PATH_DECODE_RF_U59 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6502, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6499, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5937);
   DLX_INST_DATA_PATH_DECODE_RF_U58 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6623, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6571, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630);
   DLX_INST_DATA_PATH_DECODE_RF_U57 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6606, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6577, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615);
   DLX_INST_DATA_PATH_DECODE_RF_U56 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6589, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6568, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592);
   DLX_INST_DATA_PATH_DECODE_RF_U55 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6583, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6562, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581);
   DLX_INST_DATA_PATH_DECODE_RF_U54 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5911, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5906, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5357);
   DLX_INST_DATA_PATH_DECODE_RF_U53 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6594, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6595);
   DLX_INST_DATA_PATH_DECODE_RF_U52 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6632, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6633);
   DLX_INST_DATA_PATH_DECODE_RF_U51 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5925, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5907, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5373);
   DLX_INST_DATA_PATH_DECODE_RF_U50 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5924, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5914, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5378);
   DLX_INST_DATA_PATH_DECODE_RF_U49 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5908, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5905, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5343);
   DLX_INST_DATA_PATH_DECODE_RF_U48 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6505, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6501, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5950);
   DLX_INST_DATA_PATH_DECODE_RF_U47 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6519, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6502, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5977);
   DLX_INST_DATA_PATH_DECODE_RF_U46 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6518, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6506, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5966);
   DLX_INST_DATA_PATH_DECODE_RF_U45 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6508, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6499, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5942);
   DLX_INST_DATA_PATH_DECODE_RF_U44 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6623, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6565, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624);
   DLX_INST_DATA_PATH_DECODE_RF_U43 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6606, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6574, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613);
   DLX_INST_DATA_PATH_DECODE_RF_U42 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6589, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6577, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598);
   DLX_INST_DATA_PATH_DECODE_RF_U41 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6580, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6562, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578);
   DLX_INST_DATA_PATH_DECODE_RF_U40 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5911, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5914, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5362);
   DLX_INST_DATA_PATH_DECODE_RF_U39 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6587, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6588);
   DLX_INST_DATA_PATH_DECODE_RF_U38 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6630, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6631);
   DLX_INST_DATA_PATH_DECODE_RF_U37 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5924, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5904, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5384);
   DLX_INST_DATA_PATH_DECODE_RF_U36 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5925, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5912, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5367);
   DLX_INST_DATA_PATH_DECODE_RF_U35 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6505, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6498, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5955);
   DLX_INST_DATA_PATH_DECODE_RF_U34 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6518, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6508, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5972);
   DLX_INST_DATA_PATH_DECODE_RF_U33 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6519, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6506, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5961);
   DLX_INST_DATA_PATH_DECODE_RF_U32 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6623, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6561, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621);
   DLX_INST_DATA_PATH_DECODE_RF_U31 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6606, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6565, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607);
   DLX_INST_DATA_PATH_DECODE_RF_U30 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6577, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6562, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575);
   DLX_INST_DATA_PATH_DECODE_RF_U29 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6624, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6625);
   DLX_INST_DATA_PATH_DECODE_RF_U28 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6607, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6608);
   DLX_INST_DATA_PATH_DECODE_RF_U27 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5911, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5913, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5353);
   DLX_INST_DATA_PATH_DECODE_RF_U26 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5925, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5910, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5370);
   DLX_INST_DATA_PATH_DECODE_RF_U25 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5924, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5908, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5381);
   DLX_INST_DATA_PATH_DECODE_RF_U24 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6518, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6498, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5978);
   DLX_INST_DATA_PATH_DECODE_RF_U23 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6505, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6507, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5947);
   DLX_INST_DATA_PATH_DECODE_RF_U22 : AND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6519, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6501, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5967);
   DLX_INST_DATA_PATH_DECODE_RF_U21 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6589, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6565, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590);
   DLX_INST_DATA_PATH_DECODE_RF_U20 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6621, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6622);
   DLX_INST_DATA_PATH_DECODE_RF_U19 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6600, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6601);
   DLX_INST_DATA_PATH_DECODE_RF_U18 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4484, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5190);
   DLX_INST_DATA_PATH_DECODE_RF_U17 : INV_X2 port map( A => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4483, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5189);
   DLX_INST_DATA_PATH_DECODE_RF_U16 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6619, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6620);
   DLX_INST_DATA_PATH_DECODE_RF_U15 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6615, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6616);
   DLX_INST_DATA_PATH_DECODE_RF_U14 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6613, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6614);
   DLX_INST_DATA_PATH_DECODE_RF_U13 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6598, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6599);
   DLX_INST_DATA_PATH_DECODE_RF_U12 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6592, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6593);
   DLX_INST_DATA_PATH_DECODE_RF_U11 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6590, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6591);
   DLX_INST_DATA_PATH_DECODE_RF_U10 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6581, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6582);
   DLX_INST_DATA_PATH_DECODE_RF_U9 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6578, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6579);
   DLX_INST_DATA_PATH_DECODE_RF_U8 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6575, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6576);
   DLX_INST_DATA_PATH_DECODE_RF_U7 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6572, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6573);
   DLX_INST_DATA_PATH_DECODE_RF_U6 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5193, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6566, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6567);
   DLX_INST_DATA_PATH_DECODE_RF_U5 : NAND2_X2 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5192, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6563, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6564);
   DLX_INST_DATA_PATH_DECODE_RF_U4 : OR2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5195, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5952, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4484);
   DLX_INST_DATA_PATH_DECODE_RF_U3 : OR2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5195, A2 => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5358, ZN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4483);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4131, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5294, Q => 
                           DLX_INST_DATA_PATH_A_outs_0_port, QN => n_1196);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4132, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204, Q => 
                           DLX_INST_DATA_PATH_A_outs_1_port, QN => n_1197);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4133, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203, Q => 
                           DLX_INST_DATA_PATH_A_outs_2_port, QN => n_1198);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4134, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203, Q => 
                           DLX_INST_DATA_PATH_A_outs_3_port, QN => n_1199);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4135, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203, Q => 
                           DLX_INST_DATA_PATH_A_outs_4_port, QN => n_1200);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4136, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203, Q => 
                           DLX_INST_DATA_PATH_A_outs_5_port, QN => n_1201);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4137, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202, Q => 
                           DLX_INST_DATA_PATH_A_outs_6_port, QN => n_1202);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4138, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202, Q => 
                           DLX_INST_DATA_PATH_A_outs_7_port, QN => n_1203);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4139, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202, Q => 
                           DLX_INST_DATA_PATH_A_outs_8_port, QN => n_1204);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4140, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202, Q => 
                           DLX_INST_DATA_PATH_A_outs_9_port, QN => n_1205);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_10_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4141, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201, Q => 
                           DLX_INST_DATA_PATH_A_outs_10_port, QN => n_1206);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_11_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4142, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201, Q => 
                           DLX_INST_DATA_PATH_A_outs_11_port, QN => n_1207);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_12_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4143, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201, Q => 
                           DLX_INST_DATA_PATH_A_outs_12_port, QN => n_1208);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_13_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4144, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200, Q => 
                           DLX_INST_DATA_PATH_A_outs_13_port, QN => n_1209);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_14_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4145, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200, Q => 
                           DLX_INST_DATA_PATH_A_outs_14_port, QN => n_1210);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_15_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4146, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200, Q => 
                           DLX_INST_DATA_PATH_A_outs_15_port, QN => n_1211);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_16_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4147, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200, Q => 
                           DLX_INST_DATA_PATH_A_outs_16_port, QN => n_1212);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_17_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4148, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199, Q => 
                           DLX_INST_DATA_PATH_A_outs_17_port, QN => n_1213);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_18_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4149, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199, Q => 
                           DLX_INST_DATA_PATH_A_outs_18_port, QN => n_1214);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_19_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4150, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199, Q => 
                           DLX_INST_DATA_PATH_A_outs_19_port, QN => n_1215);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_20_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4151, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199, Q => 
                           DLX_INST_DATA_PATH_A_outs_20_port, QN => n_1216);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_21_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4152, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198, Q => 
                           DLX_INST_DATA_PATH_A_outs_21_port, QN => n_1217);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_22_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4153, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198, Q => 
                           DLX_INST_DATA_PATH_A_outs_22_port, QN => n_1218);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_23_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4154, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198, Q => 
                           DLX_INST_DATA_PATH_A_outs_23_port, QN => n_1219);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_24_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4155, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197, Q => 
                           DLX_INST_DATA_PATH_A_outs_24_port, QN => n_1220);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_25_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4156, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197, Q => 
                           DLX_INST_DATA_PATH_A_outs_25_port, QN => n_1221);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_26_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4157, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197, Q => 
                           DLX_INST_DATA_PATH_A_outs_26_port, QN => n_1222);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_27_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4158, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197, Q => 
                           DLX_INST_DATA_PATH_A_outs_27_port, QN => n_1223);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_28_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4159, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196, Q => 
                           DLX_INST_DATA_PATH_A_outs_28_port, QN => n_1224);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_29_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4160, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196, Q => 
                           DLX_INST_DATA_PATH_A_outs_29_port, QN => n_1225);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_30_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4161, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196, Q => 
                           DLX_INST_DATA_PATH_A_outs_30_port, QN => n_1226);
   DLX_INST_DATA_PATH_DECODE_RF_OUT1_reg_31_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4162, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196, Q => 
                           DLX_INST_DATA_PATH_A_outs_31_port, QN => n_1227);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1303, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213, Q => n_1228, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4676);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1304, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213, Q => n_1229, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4675);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1305, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213, Q => n_1230, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4674);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1306, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213, Q => n_1231, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4673);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1307, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212, Q => n_1232, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4672);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1308, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212, Q => n_1233, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4671);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1309, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212, Q => n_1234, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4670);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1310, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212, Q => n_1235, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4669);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1311, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212, Q => n_1236, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4668);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1312, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212, Q => n_1237, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4667);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1313, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212, Q => n_1238, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4666);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1314, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212, Q => n_1239, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4665);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1315, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212, Q => n_1240, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4664);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1316, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212, Q => n_1241, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4663);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1317, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5212, Q => n_1242, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4662);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1318, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211, Q => n_1243, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4661);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1319, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211, Q => n_1244, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4660);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1320, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211, Q => n_1245, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4659);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1321, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211, Q => n_1246, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4658);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1322, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211, Q => n_1247, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4657);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1323, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211, Q => n_1248, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4656);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1324, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211, Q => n_1249, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4655);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1325, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211, Q => n_1250, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4654);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1326, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211, Q => n_1251, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4653);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1327, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211, Q => n_1252, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4652);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1328, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5211, Q => n_1253, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4651);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1329, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210, Q => n_1254, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4650);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1330, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210, Q => n_1255, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4649);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1331, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210, Q => n_1256, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4648);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1332, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210, Q => n_1257, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4647);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1333, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210, Q => n_1258, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4646);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_31_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1334, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210, Q => n_1259, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4645);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1335, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7087, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5188);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1336, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7086, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5187);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1337, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7085, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5186);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1338, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7084, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5185);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1339, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7083, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5184);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1340, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7082, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5183);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1341, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7081, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5182);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1342, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7080, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5181);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1343, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7079, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5180);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1344, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7078, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5179);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1345, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7077, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5178);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1346, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7076, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5177);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1347, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7075, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5176);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1348, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7074, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5175);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1349, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7073, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5174);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1350, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7072, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5173);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1351, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7071, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5172);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1352, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7070, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5171);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1353, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7069, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5170);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1354, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7068, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5169);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1355, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5258, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7067, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5168);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1356, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7066, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5167);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1357, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7065, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5166);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1358, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7064, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5165);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1359, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7063, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5164);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1360, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7062, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5163);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1361, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7061, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5162);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1362, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7060, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5161);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1363, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7059, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5160);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1364, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7058, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5159);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1365, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7057, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5158);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_30_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1366, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5257, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7056, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5157);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1367, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271, Q => n_1260, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4418);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1368, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271, Q => n_1261, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4417);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1369, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271, Q => n_1262, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4416);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1370, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271, Q => n_1263, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4415);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1371, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271, Q => n_1264, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4414);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1372, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271, Q => n_1265, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4413);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1373, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270, Q => n_1266, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4412);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1374, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270, Q => n_1267, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4411);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1375, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270, Q => n_1268, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4410);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1376, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270, Q => n_1269, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4409);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1377, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270, Q => n_1270, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4408);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1378, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270, Q => n_1271, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4407);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1379, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270, Q => n_1272, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4406);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1380, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270, Q => n_1273, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4405);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1381, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270, Q => n_1274, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4404);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1382, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270, Q => n_1275, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4403);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1383, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5270, Q => n_1276, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4402);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1384, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269, Q => n_1277, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4401);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1385, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269, Q => n_1278, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4400);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1386, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269, Q => n_1279, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4399);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1387, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269, Q => n_1280, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4398);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1388, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269, Q => n_1281, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4397);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1389, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269, Q => n_1282, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4396);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1390, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269, Q => n_1283, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4395);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1391, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269, Q => n_1284, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4394);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1392, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269, Q => n_1285, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4393);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1393, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269, Q => n_1286, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4392);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1394, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5269, Q => n_1287, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4391);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1395, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268, Q => n_1288, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4390);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1396, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268, Q => n_1289, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4389);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1397, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268, Q => n_1290, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4388);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_29_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1398, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268, Q => n_1291, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4387);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1399, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248, Q => n_1292, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4644);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1400, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248, Q => n_1293, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4643);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1401, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248, Q => n_1294, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4642);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1402, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247, Q => n_1295, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4641);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1403, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247, Q => n_1296, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4640);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1404, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247, Q => n_1297, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4639);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1405, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247, Q => n_1298, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4638);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1406, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247, Q => n_1299, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4637);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1407, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247, Q => n_1300, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4636);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1408, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247, Q => n_1301, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4635);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1409, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247, Q => n_1302, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4634);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1410, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247, Q => n_1303, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4633);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1411, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247, Q => n_1304, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4632);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1412, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5247, Q => n_1305, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4631);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1413, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246, Q => n_1306, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4630);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1414, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246, Q => n_1307, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4629);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1415, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246, Q => n_1308, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4628);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1416, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246, Q => n_1309, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4627);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1417, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246, Q => n_1310, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4626);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1418, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246, Q => n_1311, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4625);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1419, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246, Q => n_1312, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4624);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1420, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246, Q => n_1313, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4623);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1421, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246, Q => n_1314, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4622);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1422, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246, Q => n_1315, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4621);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1423, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5246, Q => n_1316, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4620);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1424, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245, Q => n_1317, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4619);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1425, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245, Q => n_1318, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4618);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1426, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245, Q => n_1319, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4617);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1427, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245, Q => n_1320, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4616);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1428, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245, Q => n_1321, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4615);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1429, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245, Q => n_1322, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4614);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_28_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1430, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245, Q => n_1323, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4613);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1431, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236, Q => n_1324, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4386);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1432, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236, Q => n_1325, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4385);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1433, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236, Q => n_1326, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4384);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1434, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236, Q => n_1327, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4383);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1435, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236, Q => n_1328, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4382);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1436, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236, Q => n_1329, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4381);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1437, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236, Q => n_1330, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4380);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1438, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235, Q => n_1331, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4379);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1439, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235, Q => n_1332, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4378);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1440, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235, Q => n_1333, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4377);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1441, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235, Q => n_1334, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4376);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1442, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235, Q => n_1335, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4375);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1443, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235, Q => n_1336, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4374);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1444, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235, Q => n_1337, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4373);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1445, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235, Q => n_1338, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4372);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1446, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235, Q => n_1339, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4371);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1447, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235, Q => n_1340, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4370);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1448, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5235, Q => n_1341, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4369);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1449, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234, Q => n_1342, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4368);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1450, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234, Q => n_1343, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4367);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1451, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234, Q => n_1344, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4366);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1452, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234, Q => n_1345, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4365);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1453, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234, Q => n_1346, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4364);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1454, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234, Q => n_1347, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4363);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1455, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234, Q => n_1348, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4362);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1456, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234, Q => n_1349, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4361);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1457, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234, Q => n_1350, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4360);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1458, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234, Q => n_1351, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4359);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1459, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5234, Q => n_1352, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4358);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1460, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233, Q => n_1353, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4357);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1461, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233, Q => n_1354, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4356);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_27_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1462, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233, Q => n_1355, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4355);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1463, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7055, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4964);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1464, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7054, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4963);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1465, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7053, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4962);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1466, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7052, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4961);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1467, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7051, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4960);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1468, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7050, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4959);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1469, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7049, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4958);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1470, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7048, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4957);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1471, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7047, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4956);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1472, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7046, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4955);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1473, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7045, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4954);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1474, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7044, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4953);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1475, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5282, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7043, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4952);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1476, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7042, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4951);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1477, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7041, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4950);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1478, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7040, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4949);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1479, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7039, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4948);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1480, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7038, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4947);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1481, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7037, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4946);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1482, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7036, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4945);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1483, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7035, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4944);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1484, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7034, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4943);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1485, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7033, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4942);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1486, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5281, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7032, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4941);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1487, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7031, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4940);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1488, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7030, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4939);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1489, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7029, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4938);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1490, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7028, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4937);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1491, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7027, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4936);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1492, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7026, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4935);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1493, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7025, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4934);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_26_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1494, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7024, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4933);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1495, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224, Q => n_1356, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4354);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1496, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224, Q => n_1357, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4353);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1497, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224, Q => n_1358, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4352);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1498, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224, Q => n_1359, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4351);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1499, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224, Q => n_1360, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4350);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1500, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224, Q => n_1361, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4349);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1501, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224, Q => n_1362, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4348);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1502, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224, Q => n_1363, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4347);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1503, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224, Q => n_1364, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4346);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1504, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224, Q => n_1365, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4345);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1505, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5224, Q => n_1366, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4344);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1506, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223, Q => n_1367, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4343);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1507, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223, Q => n_1368, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4342);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1508, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223, Q => n_1369, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4341);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1509, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223, Q => n_1370, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4340);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1510, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223, Q => n_1371, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4339);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1511, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223, Q => n_1372, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4338);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1512, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223, Q => n_1373, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4337);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1513, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223, Q => n_1374, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4336);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1514, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223, Q => n_1375, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4335);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1515, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223, Q => n_1376, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4334);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1516, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5223, Q => n_1377, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4333);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1517, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222, Q => n_1378, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4332);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1518, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222, Q => n_1379, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4331);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1519, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222, Q => n_1380, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4330);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1520, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222, Q => n_1381, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4329);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1521, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222, Q => n_1382, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4328);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1522, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222, Q => n_1383, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4327);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1523, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222, Q => n_1384, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4326);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1524, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222, Q => n_1385, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4325);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1525, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222, Q => n_1386, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4324);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_25_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1526, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222, Q => n_1387, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4323);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1527, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5294, Q => n_1388, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4612);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1528, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5294, Q => n_1389, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4611);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1529, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5294, Q => n_1390, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4610);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1530, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5294, Q => n_1391, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4609);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1531, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5294, Q => n_1392, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4608);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1532, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5294, Q => n_1393, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4607);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1533, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5294, Q => n_1394, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4606);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1534, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5294, Q => n_1395, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4605);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1535, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293, Q => n_1396, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4604);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1536, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293, Q => n_1397, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4603);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1537, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293, Q => n_1398, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4602);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1538, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293, Q => n_1399, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4601);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1539, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293, Q => n_1400, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4600);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1540, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293, Q => n_1401, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4599);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1541, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293, Q => n_1402, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4598);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1542, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293, Q => n_1403, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4597);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1543, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293, Q => n_1404, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4596);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1544, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293, Q => n_1405, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4595);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1545, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5293, Q => n_1406, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4594);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1546, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292, Q => n_1407, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4593);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1547, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292, Q => n_1408, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4592);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1548, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292, Q => n_1409, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4591);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1549, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292, Q => n_1410, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4590);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1550, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292, Q => n_1411, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4589);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1551, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292, Q => n_1412, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4588);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1552, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292, Q => n_1413, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4587);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1553, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292, Q => n_1414, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4586);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1554, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292, Q => n_1415, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4585);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1555, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292, Q => n_1416, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4584);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1556, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5292, Q => n_1417, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4583);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1557, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291, Q => n_1418, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4582);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_24_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1558, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291, Q => n_1419, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4581);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1559, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210, Q => n_1420, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4580);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1560, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210, Q => n_1421, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4579);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1561, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210, Q => n_1422, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4578);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1562, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210, Q => n_1423, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4577);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1563, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5210, Q => n_1424, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4576);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1564, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209, Q => n_1425, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4575);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1565, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209, Q => n_1426, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4574);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1566, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209, Q => n_1427, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4573);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1567, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209, Q => n_1428, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4572);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1568, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209, Q => n_1429, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4571);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1569, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209, Q => n_1430, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4570);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1570, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209, Q => n_1431, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4569);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1571, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209, Q => n_1432, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4568);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1572, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209, Q => n_1433, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4567);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1573, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209, Q => n_1434, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4566);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1574, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5209, Q => n_1435, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4565);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1575, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208, Q => n_1436, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4564);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1576, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208, Q => n_1437, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4563);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1577, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208, Q => n_1438, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4562);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1578, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208, Q => n_1439, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4561);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1579, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208, Q => n_1440, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4560);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1580, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208, Q => n_1441, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4559);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1581, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208, Q => n_1442, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4558);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1582, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208, Q => n_1443, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4557);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1583, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208, Q => n_1444, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4556);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1584, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208, Q => n_1445, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4555);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1585, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5208, Q => n_1446, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4554);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1586, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207, Q => n_1447, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4553);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1587, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207, Q => n_1448, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4552);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1588, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207, Q => n_1449, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4551);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1589, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207, Q => n_1450, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4550);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_23_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1590, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207, Q => n_1451, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4549);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1591, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7023, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4932);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1592, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7022, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4931);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1593, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7021, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4930);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1594, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7020, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4929);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1595, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7019, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4928);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1596, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7018, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4927);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1597, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7017, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4926);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1598, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7016, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4925);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1599, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7015, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4924);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1600, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7014, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4923);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1601, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5256, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7013, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4922);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1602, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7012, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4921);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1603, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7011, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4920);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1604, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7010, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4919);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1605, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7009, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4918);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1606, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7008, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4917);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1607, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7007, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4916);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1608, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7006, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4915);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1609, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7005, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4914);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1610, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7004, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4913);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1611, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7003, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4912);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1612, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5255, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7002, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4911);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1613, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7001, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4910);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1614, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n7000, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4909);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1615, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6999, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4908);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1616, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6998, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4907);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1617, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6997, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4906);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1618, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6996, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4905);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1619, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6995, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4904);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1620, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6994, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4903);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1621, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6993, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4902);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_22_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1622, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6992, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4901);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1623, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268, Q => n_1452, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4322);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1624, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268, Q => n_1453, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4321);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1625, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268, Q => n_1454, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4320);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1626, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268, Q => n_1455, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4319);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1627, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268, Q => n_1456, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4318);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1628, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268, Q => n_1457, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4317);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1629, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5268, Q => n_1458, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4316);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1630, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267, Q => n_1459, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4315);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1631, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267, Q => n_1460, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4314);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1632, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267, Q => n_1461, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4313);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1633, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267, Q => n_1462, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4312);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1634, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267, Q => n_1463, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4311);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1635, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267, Q => n_1464, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4310);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1636, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267, Q => n_1465, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4309);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1637, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267, Q => n_1466, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4308);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1638, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267, Q => n_1467, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4307);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1639, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267, Q => n_1468, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4306);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1640, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5267, Q => n_1469, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4305);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1641, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266, Q => n_1470, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4304);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1642, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266, Q => n_1471, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4303);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1643, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266, Q => n_1472, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4302);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1644, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266, Q => n_1473, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4301);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1645, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266, Q => n_1474, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4300);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1646, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266, Q => n_1475, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4299);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1647, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266, Q => n_1476, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4298);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1648, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266, Q => n_1477, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4297);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1649, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266, Q => n_1478, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4296);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1650, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266, Q => n_1479, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4295);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1651, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5266, Q => n_1480, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4294);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1652, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265, Q => n_1481, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4293);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1653, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265, Q => n_1482, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4292);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_21_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1654, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265, Q => n_1483, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4291);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1655, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245, Q => n_1484, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4290);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1656, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245, Q => n_1485, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4289);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1657, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245, Q => n_1486, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4288);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1658, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5245, Q => n_1487, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4287);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1659, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244, Q => n_1488, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4286);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1660, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244, Q => n_1489, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4285);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1661, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244, Q => n_1490, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4284);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1662, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244, Q => n_1491, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4283);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1663, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244, Q => n_1492, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4282);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1664, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244, Q => n_1493, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4281);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1665, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244, Q => n_1494, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4280);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1666, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244, Q => n_1495, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4279);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1667, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244, Q => n_1496, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4278);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1668, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244, Q => n_1497, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4277);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1669, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5244, Q => n_1498, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4276);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1670, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243, Q => n_1499, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4275);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1671, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243, Q => n_1500, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4274);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1672, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243, Q => n_1501, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4273);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1673, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243, Q => n_1502, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4272);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1674, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243, Q => n_1503, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4271);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1675, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243, Q => n_1504, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4270);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1676, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243, Q => n_1505, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4269);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1677, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243, Q => n_1506, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4268);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1678, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243, Q => n_1507, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4267);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1679, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243, Q => n_1508, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4266);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1680, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5243, Q => n_1509, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4265);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1681, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242, Q => n_1510, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4264);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1682, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242, Q => n_1511, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4263);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1683, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242, Q => n_1512, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4262);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1684, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242, Q => n_1513, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4261);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1685, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242, Q => n_1514, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4260);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_20_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1686, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242, Q => n_1515, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4259);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1687, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6927, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4900);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1688, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6926, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4899);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1689, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6925, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4898);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1690, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6924, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4897);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1691, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6923, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4896);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1692, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6922, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4895);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1693, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6921, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4894);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1694, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5233, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6920, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4893);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1695, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6919, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4892);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1696, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6918, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4891);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1697, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6917, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4890);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1698, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6916, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4889);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1699, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6915, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4888);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1700, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6914, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4887);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1701, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6913, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4886);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1702, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6912, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4885);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1703, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6911, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4884);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1704, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6910, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4883);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1705, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5232, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6909, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4882);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1706, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6908, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4881);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1707, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6907, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4880);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1708, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6906, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4879);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1709, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6905, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4878);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1710, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6904, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4877);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1711, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6903, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4876);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1712, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6902, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4875);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1713, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6901, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4874);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1714, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6900, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4873);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1715, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6899, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4872);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1716, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5231, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6898, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4871);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1717, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6897, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4870);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_19_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1718, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6896, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4869);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1719, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6991, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5156);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1720, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6990, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5155);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1721, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5280, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6989, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5154);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1722, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6988, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5153);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1723, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6987, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5152);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1724, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6986, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5151);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1725, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6985, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5150);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1726, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6984, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5149);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1727, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6983, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5148);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1728, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6982, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5147);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1729, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6981, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5146);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1730, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6980, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5145);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1731, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6979, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5144);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1732, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5279, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6978, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5143);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1733, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6977, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5142);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1734, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6976, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5141);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1735, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6975, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5140);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1736, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6974, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5139);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1737, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6973, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5138);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1738, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6972, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5137);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1739, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6971, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5136);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1740, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6970, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5135);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1741, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6969, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5134);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1742, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6968, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5133);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1743, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5278, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6967, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5132);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1744, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6966, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5131);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1745, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6965, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5130);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1746, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6964, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5129);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1747, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6963, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5128);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1748, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6962, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5127);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1749, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6961, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5126);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_18_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1750, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6960, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5125);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1751, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5222, Q => n_1516, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4548);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1752, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221, Q => n_1517, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4547);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1753, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221, Q => n_1518, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4546);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1754, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221, Q => n_1519, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4545);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1755, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221, Q => n_1520, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4544);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1756, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221, Q => n_1521, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4543);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1757, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221, Q => n_1522, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4542);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1758, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221, Q => n_1523, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4541);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1759, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221, Q => n_1524, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4540);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1760, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221, Q => n_1525, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4539);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1761, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221, Q => n_1526, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4538);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1762, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5221, Q => n_1527, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4537);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1763, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220, Q => n_1528, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4536);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1764, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220, Q => n_1529, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4535);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1765, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220, Q => n_1530, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4534);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1766, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220, Q => n_1531, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4533);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1767, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220, Q => n_1532, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4532);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1768, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220, Q => n_1533, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4531);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1769, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220, Q => n_1534, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4530);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1770, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220, Q => n_1535, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4529);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1771, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220, Q => n_1536, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4528);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1772, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220, Q => n_1537, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4527);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1773, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5220, Q => n_1538, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4526);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1774, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219, Q => n_1539, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4525);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1775, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219, Q => n_1540, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4524);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1776, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219, Q => n_1541, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4523);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1777, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219, Q => n_1542, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4522);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1778, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219, Q => n_1543, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4521);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1779, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219, Q => n_1544, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4520);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1780, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219, Q => n_1545, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4519);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1781, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219, Q => n_1546, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4518);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_17_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1782, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219, Q => n_1547, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4517);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1783, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6959, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5124);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1784, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6958, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5123);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1785, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6957, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5122);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1786, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6956, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5121);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1787, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6955, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5120);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1788, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6954, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5119);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1789, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6953, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5118);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1790, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6952, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5117);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1791, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5291, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6951, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5116);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1792, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6950, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5115);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1793, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6949, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5114);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1794, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6948, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5113);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1795, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6947, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5112);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1796, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6946, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5111);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1797, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6945, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5110);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1798, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6944, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5109);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1799, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6943, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5108);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1800, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6942, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5107);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1801, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6941, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5106);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1802, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5290, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6940, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5105);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1803, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6939, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5104);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1804, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6938, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5103);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1805, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6937, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5102);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1806, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6936, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5101);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1807, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6935, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5100);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1808, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6934, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5099);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1809, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6933, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5098);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1810, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6932, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5097);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1811, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6931, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5096);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1812, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6930, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5095);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1813, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5289, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6929, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5094);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_16_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1814, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6928, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5093);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1815, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6895, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4868);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1816, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6894, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4867);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1817, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6893, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4866);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1818, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6892, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4865);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1819, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6891, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4864);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1820, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5207, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6890, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4863);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1821, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6889, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4862);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1822, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6888, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4861);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1823, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6887, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4860);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1824, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6886, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4859);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1825, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6885, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4858);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1826, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6884, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4857);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1827, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6883, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4856);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1828, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6882, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4855);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1829, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6881, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4854);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1830, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6880, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4853);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1831, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5206, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6879, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4852);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1832, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6878, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4851);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1833, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6877, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4850);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1834, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6876, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4849);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1835, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6875, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4848);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1836, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6874, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4847);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1837, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6873, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4846);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1838, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6872, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4845);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1839, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6871, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4844);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1840, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6870, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4843);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1841, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6869, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4842);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1842, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5205, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6868, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4841);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1843, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6867, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4840);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1844, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6866, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4839);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1845, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6865, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4838);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_15_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1846, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6864, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4837);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1847, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5254, Q => n_1548, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4482);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1848, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253, Q => n_1549, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4481);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1849, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253, Q => n_1550, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4480);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1850, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253, Q => n_1551, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4479);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1851, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253, Q => n_1552, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4478);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1852, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253, Q => n_1553, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4477);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1853, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253, Q => n_1554, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4476);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1854, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253, Q => n_1555, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4475);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1855, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253, Q => n_1556, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4474);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1856, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253, Q => n_1557, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4473);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1857, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253, Q => n_1558, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4472);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1858, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5253, Q => n_1559, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4471);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1859, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252, Q => n_1560, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4470);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1860, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252, Q => n_1561, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4469);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1861, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252, Q => n_1562, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4468);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1862, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252, Q => n_1563, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4467);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1863, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252, Q => n_1564, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4466);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1864, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252, Q => n_1565, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4465);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1865, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252, Q => n_1566, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4464);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1866, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252, Q => n_1567, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4463);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1867, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252, Q => n_1568, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4462);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1868, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252, Q => n_1569, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4461);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1869, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5252, Q => n_1570, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4460);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1870, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251, Q => n_1571, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4459);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1871, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251, Q => n_1572, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4458);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1872, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251, Q => n_1573, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4457);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1873, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251, Q => n_1574, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4456);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1874, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251, Q => n_1575, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4455);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1875, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251, Q => n_1576, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4454);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1876, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251, Q => n_1577, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4453);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1877, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251, Q => n_1578, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4452);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_14_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1878, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251, Q => n_1579, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4451);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1879, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265, Q => n_1580, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4740);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1880, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265, Q => n_1581, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4739);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1881, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265, Q => n_1582, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4738);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1882, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265, Q => n_1583, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4737);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1883, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265, Q => n_1584, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4736);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1884, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265, Q => n_1585, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4735);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1885, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265, Q => n_1586, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4734);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1886, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5265, Q => n_1587, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4733);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1887, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264, Q => n_1588, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4732);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1888, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264, Q => n_1589, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4731);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1889, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264, Q => n_1590, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4730);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1890, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264, Q => n_1591, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4729);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1891, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264, Q => n_1592, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4728);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1892, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264, Q => n_1593, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4727);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1893, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264, Q => n_1594, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4726);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1894, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264, Q => n_1595, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4725);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1895, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264, Q => n_1596, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4724);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1896, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264, Q => n_1597, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4723);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1897, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5264, Q => n_1598, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4722);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1898, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263, Q => n_1599, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4721);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1899, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263, Q => n_1600, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4720);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1900, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263, Q => n_1601, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4719);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1901, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263, Q => n_1602, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4718);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1902, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263, Q => n_1603, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4717);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1903, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263, Q => n_1604, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4716);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1904, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263, Q => n_1605, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4715);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1905, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263, Q => n_1606, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4714);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1906, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263, Q => n_1607, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4713);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1907, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263, Q => n_1608, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4712);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1908, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5263, Q => n_1609, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4711);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1909, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262, Q => n_1610, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4710);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_13_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1910, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262, Q => n_1611, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4709);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1911, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6863, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5092);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1912, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6862, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5091);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1913, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6861, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5090);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1914, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6860, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5089);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1915, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5242, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6859, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5088);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1916, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6858, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5087);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1917, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6857, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5086);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1918, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6856, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5085);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1919, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6855, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5084);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1920, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6854, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5083);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1921, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6853, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5082);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1922, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6852, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5081);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1923, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6851, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5080);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1924, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6850, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5079);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1925, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6849, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5078);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1926, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5241, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6848, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5077);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1927, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6847, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5076);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1928, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6846, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5075);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1929, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6845, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5074);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1930, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6844, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5073);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1931, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6843, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5072);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1932, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6842, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5071);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1933, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6841, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5070);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1934, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6840, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5069);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1935, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6839, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5068);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1936, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6838, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5067);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1937, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5240, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6837, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5066);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1938, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6836, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5065);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1939, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6835, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5064);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1940, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6834, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5063);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1941, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6833, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5062);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_12_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1942, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6832, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5061);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1943, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6831, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5060);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1944, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6830, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5059);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1945, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6829, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5058);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1946, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6828, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5057);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1947, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6827, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5056);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1948, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6826, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5055);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1949, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6825, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5054);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1950, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6824, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5053);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1951, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5230, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6823, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5052);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1952, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6822, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5051);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1953, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6821, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5050);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1954, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6820, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5049);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1955, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6819, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5048);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1956, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6818, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5047);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1957, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6817, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5046);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1958, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6816, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5045);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1959, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6815, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5044);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1960, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6814, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5043);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1961, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6813, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5042);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1962, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5229, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6812, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5041);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1963, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6811, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5040);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1964, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6810, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5039);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1965, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6809, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5038);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1966, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6808, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5037);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1967, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6807, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5036);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1968, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6806, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5035);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1969, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6805, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5034);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1970, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6804, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5033);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1971, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6803, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5032);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1972, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6802, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5031);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1973, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5228, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6801, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5030);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_11_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1974, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6800, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5029);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_0_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1975, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277, Q => n_1612, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4226);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_1_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1976, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277, Q => n_1613, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4225);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_2_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1977, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277, Q => n_1614, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4224);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_3_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1978, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5277, Q => n_1615, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4223);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_4_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1979, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276, Q => n_1616, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4222);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_5_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1980, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276, Q => n_1617, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4221);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_6_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1981, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276, Q => n_1618, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4220);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_7_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1982, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276, Q => n_1619, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4219);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_8_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1983, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276, Q => n_1620, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4218);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_9_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n1984, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276, Q => n_1621, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4217);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_10_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1985, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276, Q => n_1622, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4216);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_11_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1986, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276, Q => n_1623, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4215);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_12_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1987, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276, Q => n_1624, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4214);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_13_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1988, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276, Q => n_1625, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4213);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_14_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1989, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5276, Q => n_1626, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4212);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_15_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1990, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275, Q => n_1627, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4211);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_16_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1991, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275, Q => n_1628, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4210);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_17_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1992, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275, Q => n_1629, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4209);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_18_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1993, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275, Q => n_1630, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4208);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_19_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1994, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275, Q => n_1631, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4207);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_20_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1995, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275, Q => n_1632, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4206);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_21_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1996, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275, Q => n_1633, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4205);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_22_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1997, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275, Q => n_1634, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4204);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_23_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1998, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275, Q => n_1635, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4203);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_24_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n1999, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275, Q => n_1636, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4202);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_25_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n2000, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5275, Q => n_1637, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4201);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_26_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n2001, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274, Q => n_1638, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4200);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_27_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n2002, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274, Q => n_1639, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4199);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_28_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n2003, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274, Q => n_1640, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4198);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_29_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n2004, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274, Q => n_1641, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4197);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_30_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n2005, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274, Q => n_1642, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4196);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_10_31_inst : DFF_X1 port map( D 
                           => DLX_INST_DATA_PATH_DECODE_RF_n2006, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274, Q => n_1643, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4195);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2007, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219, Q => n_1644, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4258);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2008, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5219, Q => n_1645, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4257);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2009, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218, Q => n_1646, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4256);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2010, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218, Q => n_1647, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4255);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2011, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218, Q => n_1648, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4254);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2012, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218, Q => n_1649, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4253);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2013, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218, Q => n_1650, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4252);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2014, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218, Q => n_1651, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4251);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2015, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218, Q => n_1652, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4250);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2016, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218, Q => n_1653, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4249);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_10_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2017, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218, Q => n_1654, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4248);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_11_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2018, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218, Q => n_1655, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4247);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_12_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2019, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5218, Q => n_1656, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4246);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_13_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2020, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217, Q => n_1657, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4245);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_14_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2021, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217, Q => n_1658, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4244);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_15_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2022, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217, Q => n_1659, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4243);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_16_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2023, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217, Q => n_1660, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4242);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_17_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2024, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217, Q => n_1661, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4241);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_18_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2025, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217, Q => n_1662, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4240);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_19_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2026, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217, Q => n_1663, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4239);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_20_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2027, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217, Q => n_1664, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4238);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_21_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2028, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217, Q => n_1665, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4237);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_22_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2029, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217, Q => n_1666, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4236);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_23_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2030, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5217, Q => n_1667, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4235);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_24_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2031, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216, Q => n_1668, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4234);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_25_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2032, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216, Q => n_1669, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4233);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_26_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2033, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216, Q => n_1670, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4232);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_27_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2034, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216, Q => n_1671, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4231);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_28_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2035, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216, Q => n_1672, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4230);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_29_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2036, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216, Q => n_1673, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4229);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_30_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2037, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216, Q => n_1674, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4228);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_9_31_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2038, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216, Q => n_1675, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4227);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2039, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6799, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4836);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2040, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6798, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4835);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2041, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6797, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4834);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2042, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6796, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4833);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2043, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6795, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4832);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2044, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6794, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4831);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2045, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6793, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4830);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2046, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6792, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4829);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2047, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6791, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4828);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2048, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5288, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6790, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4827);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_10_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2049, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6789, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4826);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_11_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2050, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6788, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4825);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_12_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2051, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6787, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4824);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_13_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2052, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6786, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4823);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_14_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2053, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6785, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4822);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_15_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2054, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6784, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4821);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_16_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2055, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6783, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4820);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_17_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2056, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6782, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4819);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_18_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2057, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6781, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4818);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_19_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2058, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6780, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4817);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_20_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2059, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5287, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6779, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4816);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_21_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2060, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6778, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4815);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_22_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2061, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6777, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4814);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_23_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2062, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6776, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4813);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_24_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2063, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6775, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4812);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_25_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2064, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6774, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4811);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_26_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2065, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6773, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4810);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_27_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2066, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6772, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4809);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_28_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2067, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6771, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4808);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_29_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2068, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6770, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4807);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_30_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2069, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6769, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4806);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_8_31_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2070, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5286, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6768, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4805);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2071, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204, Q => n_1676, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4450);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2072, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204, Q => n_1677, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4449);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2073, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204, Q => n_1678, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4448);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2074, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203, Q => n_1679, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4447);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2075, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203, Q => n_1680, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4446);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2076, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203, Q => n_1681, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4445);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2077, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203, Q => n_1682, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4444);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2078, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202, Q => n_1683, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4443);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2079, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202, Q => n_1684, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4442);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2080, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202, Q => n_1685, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4441);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_10_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2081, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201, Q => n_1686, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4440);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_11_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2082, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201, Q => n_1687, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4439);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_12_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2083, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201, Q => n_1688, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4438);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_13_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2084, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201, Q => n_1689, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4437);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_14_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2085, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200, Q => n_1690, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4436);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_15_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2086, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200, Q => n_1691, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4435);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_16_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2087, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200, Q => n_1692, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4434);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_17_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2088, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200, Q => n_1693, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4433);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_18_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2089, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199, Q => n_1694, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4432);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_19_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2090, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199, Q => n_1695, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4431);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_20_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2091, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199, Q => n_1696, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4430);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_21_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2092, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198, Q => n_1697, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4429);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_22_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2093, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198, Q => n_1698, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4428);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_23_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2094, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198, Q => n_1699, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4427);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_24_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2095, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198, Q => n_1700, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4426);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_25_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2096, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197, Q => n_1701, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4425);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_26_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2097, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197, Q => n_1702, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4424);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_27_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2098, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197, Q => n_1703, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4423);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_28_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2099, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197, Q => n_1704, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4422);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_29_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2100, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196, Q => n_1705, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4421);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_30_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2101, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196, Q => n_1706, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4420);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_7_31_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2102, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196, Q => n_1707, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4419);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2103, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251, Q => n_1708, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4708);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2104, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5251, Q => n_1709, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4707);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2105, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250, Q => n_1710, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4706);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2106, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250, Q => n_1711, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4705);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2107, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250, Q => n_1712, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4704);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2108, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250, Q => n_1713, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4703);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2109, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250, Q => n_1714, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4702);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2110, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250, Q => n_1715, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4701);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2111, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250, Q => n_1716, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4700);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2112, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250, Q => n_1717, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4699);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_10_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2113, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250, Q => n_1718, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4698);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_11_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2114, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250, Q => n_1719, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4697);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_12_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2115, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5250, Q => n_1720, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4696);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_13_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2116, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249, Q => n_1721, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4695);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_14_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2117, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249, Q => n_1722, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4694);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_15_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2118, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249, Q => n_1723, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4693);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_16_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2119, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249, Q => n_1724, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4692);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_17_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2120, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249, Q => n_1725, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4691);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_18_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2121, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249, Q => n_1726, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4690);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_19_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2122, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249, Q => n_1727, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4689);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_20_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2123, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249, Q => n_1728, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4688);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_21_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2124, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249, Q => n_1729, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4687);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_22_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2125, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249, Q => n_1730, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4686);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_23_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2126, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5249, Q => n_1731, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4685);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_24_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2127, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248, Q => n_1732, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4684);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_25_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2128, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248, Q => n_1733, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4683);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_26_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2129, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248, Q => n_1734, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4682);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_27_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2130, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248, Q => n_1735, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4681);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_28_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2131, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248, Q => n_1736, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4680);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_29_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2132, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248, Q => n_1737, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4679);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_30_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2133, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248, Q => n_1738, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4678);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_6_31_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2134, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5248, Q => n_1739, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4677);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2135, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262, Q => n_1740, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4194);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2136, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262, Q => n_1741, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4193);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2137, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262, Q => n_1742, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4192);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2138, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262, Q => n_1743, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4191);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2139, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262, Q => n_1744, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4190);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2140, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262, Q => n_1745, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4189);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2141, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262, Q => n_1746, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4188);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2142, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262, Q => n_1747, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4187);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2143, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5262, Q => n_1748, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4186);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2144, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261, Q => n_1749, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4185);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_10_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2145, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261, Q => n_1750, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4184);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_11_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2146, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261, Q => n_1751, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4183);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_12_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2147, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261, Q => n_1752, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4182);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_13_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2148, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261, Q => n_1753, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4181);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_14_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2149, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261, Q => n_1754, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4180);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_15_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2150, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261, Q => n_1755, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4179);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_16_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2151, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261, Q => n_1756, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4178);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_17_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2152, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261, Q => n_1757, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4177);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_18_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2153, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261, Q => n_1758, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4176);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_19_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2154, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5261, Q => n_1759, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4175);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_20_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2155, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260, Q => n_1760, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4174);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_21_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2156, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260, Q => n_1761, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4173);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_22_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2157, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260, Q => n_1762, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4172);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_23_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2158, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260, Q => n_1763, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4171);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_24_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2159, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260, Q => n_1764, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4170);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_25_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2160, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260, Q => n_1765, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4169);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_26_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2161, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260, Q => n_1766, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4168);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_27_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2162, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260, Q => n_1767, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4167);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_28_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2163, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260, Q => n_1768, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4166);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_29_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2164, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260, Q => n_1769, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4165);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_30_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2165, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5260, Q => n_1770, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4164);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_5_31_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2166, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5259, Q => n_1771, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4163);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2167, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6767, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4804);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2168, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6766, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4803);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2169, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6765, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4802);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2170, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6764, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4801);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2171, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6763, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4800);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2172, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5239, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6762, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4799);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2173, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6761, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4798);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2174, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6760, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4797);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2175, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6759, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4796);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2176, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6758, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4795);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_10_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2177, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6757, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4794);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_11_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2178, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6756, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4793);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_12_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2179, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6755, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4792);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_13_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2180, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6754, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4791);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_14_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2181, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6753, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4790);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_15_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2182, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6752, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4789);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_16_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2183, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5238, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6751, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4788);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_17_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2184, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6750, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4787);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_18_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2185, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6749, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4786);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_19_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2186, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6748, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4785);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_20_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2187, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6747, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4784);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_21_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2188, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6746, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4783);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_22_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2189, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6745, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4782);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_23_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2190, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6744, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4781);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_24_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2191, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6743, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4780);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_25_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2192, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6742, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4779);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_26_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2193, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6741, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4778);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_27_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2194, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5237, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6740, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4777);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_28_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2195, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6739, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4776);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_29_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2196, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6738, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4775);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_30_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2197, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6737, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4774);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_4_31_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2198, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5236, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6736, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4773);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2199, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6735, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4772);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2200, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6734, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4771);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2201, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6733, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4770);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2202, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6732, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4769);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2203, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6731, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4768);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2204, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6730, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4767);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2205, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6729, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4766);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2206, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6728, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4765);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2207, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6727, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4764);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2208, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5227, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6726, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4763);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_10_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2209, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6725, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4762);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_11_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2210, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6724, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4761);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_12_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2211, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6723, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4760);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_13_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2212, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6722, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4759);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_14_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2213, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6721, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4758);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_15_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2214, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6720, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4757);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_16_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2215, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6719, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4756);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_17_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2216, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6718, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4755);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_18_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2217, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6717, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4754);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_19_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2218, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6716, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4753);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_20_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2219, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5226, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6715, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4752);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_21_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2220, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6714, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4751);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_22_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2221, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6713, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4750);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_23_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2222, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6712, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4749);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_24_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2223, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6711, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4748);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_25_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2224, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6710, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4747);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_26_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2225, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6709, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4746);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_27_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2226, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6708, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4745);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_28_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2227, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6707, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4744);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_29_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2228, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6706, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4743);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_30_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2229, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6705, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4742);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_3_31_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2230, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5225, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6704, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4741);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2231, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6703, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5028);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2232, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6702, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5027);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2233, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6701, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5026);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2234, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6700, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5025);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2235, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5274, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6699, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5024);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2236, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6698, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5023);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2237, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6697, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5022);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2238, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6696, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5021);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2239, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6695, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5020);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2240, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6694, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5019);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_10_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2241, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6693, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5018);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_11_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2242, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6692, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5017);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_12_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2243, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6691, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5016);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_13_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2244, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6690, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5015);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_14_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2245, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6689, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5014);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_15_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2246, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5273, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6688, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5013);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_16_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2247, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6687, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5012);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_17_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2248, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6686, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5011);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_18_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2249, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6685, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5010);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_19_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2250, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6684, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5009);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_20_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2251, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6683, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5008);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_21_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2252, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6682, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5007);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_22_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2253, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6681, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5006);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_23_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2254, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6680, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5005);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_24_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2255, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6679, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5004);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_25_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2256, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6678, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5003);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_26_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2257, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5272, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6677, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5002);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_27_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2258, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6676, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5001);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_28_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2259, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6675, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5000);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_29_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2260, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6674, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4999);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_30_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2261, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6673, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4998);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_2_31_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2262, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5271, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6672, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4997);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2263, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6671, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4996);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2264, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6670, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4995);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2265, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5216, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6669, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4994);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2266, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6668, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4993);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2267, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6667, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4992);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2268, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6666, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4991);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2269, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6665, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4990);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2270, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6664, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4989);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2271, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6663, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4988);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2272, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6662, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4987);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_10_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2273, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6661, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4986);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_11_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2274, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6660, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4985);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_12_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2275, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6659, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4984);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_13_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2276, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5215, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6658, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4983);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_14_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2277, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6657, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4982);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_15_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2278, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6656, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4981);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_16_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2279, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6655, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4980);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_17_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2280, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6654, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4979);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_18_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2281, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6653, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4978);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_19_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2282, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6652, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4977);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_20_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2283, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6651, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4976);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_21_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2284, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6650, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4975);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_22_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2285, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6649, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4974);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_23_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2286, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6648, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4973);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_24_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2287, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5214, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6647, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4972);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_25_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2288, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6646, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4971);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_26_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2289, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6645, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4970);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_27_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2290, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6644, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4969);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_28_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2291, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6643, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4968);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_29_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2292, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6642, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4967);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_30_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2293, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6641, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4966);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_1_31_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2294, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5213, Q => 
                           DLX_INST_DATA_PATH_DECODE_RF_n6640, QN => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4965);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2295, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5294, Q => n_1772, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4516);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2296, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285, Q => n_1773, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4515);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2297, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285, Q => n_1774, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4514);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2298, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285, Q => n_1775, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4513);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2299, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285, Q => n_1776, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4512);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2300, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285, Q => n_1777, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4511);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2301, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285, Q => n_1778, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4510);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2302, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285, Q => n_1779, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4509);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2303, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285, Q => n_1780, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4508);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n2304, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285, Q => n_1781, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4507);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_10_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2305, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285, Q => n_1782, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4506);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_11_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2306, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5285, Q => n_1783, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4505);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_12_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2307, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284, Q => n_1784, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4504);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_13_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2308, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284, Q => n_1785, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4503);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_14_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2309, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284, Q => n_1786, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4502);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_15_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2310, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284, Q => n_1787, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4501);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_16_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2311, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284, Q => n_1788, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4500);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_17_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2312, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284, Q => n_1789, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4499);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_18_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2313, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284, Q => n_1790, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4498);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_19_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2314, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284, Q => n_1791, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4497);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_20_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2315, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284, Q => n_1792, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4496);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_21_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2316, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284, Q => n_1793, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4495);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_22_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2317, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5284, Q => n_1794, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4494);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_23_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2318, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283, Q => n_1795, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4493);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_24_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2319, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283, Q => n_1796, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4492);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_25_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2320, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283, Q => n_1797, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4491);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_26_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2321, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283, Q => n_1798, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4490);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_27_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2322, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283, Q => n_1799, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4489);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_28_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2323, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283, Q => n_1800, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4488);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_29_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2324, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283, Q => n_1801, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4487);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_30_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2325, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283, Q => n_1802, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4486);
   DLX_INST_DATA_PATH_DECODE_RF_REGISTERS_reg_0_31_inst : DFF_X1 port map( D =>
                           DLX_INST_DATA_PATH_DECODE_RF_n2326, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5283, Q => n_1803, QN 
                           => DLX_INST_DATA_PATH_DECODE_RF_n4485);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_0_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4099, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204, Q => 
                           DLX_INST_DATA_PATH_B_outs_0_port, QN => n_1804);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_1_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4100, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204, Q => 
                           DLX_INST_DATA_PATH_B_outs_1_port, QN => n_1805);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_2_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4101, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5204, Q => 
                           DLX_INST_DATA_PATH_B_outs_2_port, QN => n_1806);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_3_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4102, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203, Q => 
                           DLX_INST_DATA_PATH_B_outs_3_port, QN => n_1807);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_4_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4103, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203, Q => 
                           DLX_INST_DATA_PATH_B_outs_4_port, QN => n_1808);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_5_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4104, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5203, Q => 
                           DLX_INST_DATA_PATH_B_outs_5_port, QN => n_1809);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_6_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4105, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202, Q => 
                           DLX_INST_DATA_PATH_B_outs_6_port, QN => n_1810);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_7_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4106, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202, Q => 
                           DLX_INST_DATA_PATH_B_outs_7_port, QN => n_1811);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_8_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4107, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202, Q => 
                           DLX_INST_DATA_PATH_B_outs_8_port, QN => n_1812);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_9_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4108, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5202, Q => 
                           DLX_INST_DATA_PATH_B_outs_9_port, QN => n_1813);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_10_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4109, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201, Q => 
                           DLX_INST_DATA_PATH_B_outs_10_port, QN => n_1814);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_11_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4110, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201, Q => 
                           DLX_INST_DATA_PATH_B_outs_11_port, QN => n_1815);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_12_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4111, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201, Q => 
                           DLX_INST_DATA_PATH_B_outs_12_port, QN => n_1816);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_13_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4112, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5201, Q => 
                           DLX_INST_DATA_PATH_B_outs_13_port, QN => n_1817);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_14_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4113, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200, Q => 
                           DLX_INST_DATA_PATH_B_outs_14_port, QN => n_1818);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_15_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4114, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200, Q => 
                           DLX_INST_DATA_PATH_B_outs_15_port, QN => n_1819);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_16_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4115, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5200, Q => 
                           DLX_INST_DATA_PATH_B_outs_16_port, QN => n_1820);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_17_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4116, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199, Q => 
                           DLX_INST_DATA_PATH_B_outs_17_port, QN => n_1821);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_18_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4117, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199, Q => 
                           DLX_INST_DATA_PATH_B_outs_18_port, QN => n_1822);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_19_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4118, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199, Q => 
                           DLX_INST_DATA_PATH_B_outs_19_port, QN => n_1823);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_20_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4119, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5199, Q => 
                           DLX_INST_DATA_PATH_B_outs_20_port, QN => n_1824);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_21_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4120, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198, Q => 
                           DLX_INST_DATA_PATH_B_outs_21_port, QN => n_1825);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_22_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4121, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198, Q => 
                           DLX_INST_DATA_PATH_B_outs_22_port, QN => n_1826);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_23_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4122, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198, Q => 
                           DLX_INST_DATA_PATH_B_outs_23_port, QN => n_1827);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_24_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4123, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5198, Q => 
                           DLX_INST_DATA_PATH_B_outs_24_port, QN => n_1828);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_25_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4124, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197, Q => 
                           DLX_INST_DATA_PATH_B_outs_25_port, QN => n_1829);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_26_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4125, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197, Q => 
                           DLX_INST_DATA_PATH_B_outs_26_port, QN => n_1830);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_27_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4126, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5197, Q => 
                           DLX_INST_DATA_PATH_B_outs_27_port, QN => n_1831);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_28_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4127, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196, Q => 
                           DLX_INST_DATA_PATH_B_outs_28_port, QN => n_1832);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_29_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4128, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196, Q => 
                           DLX_INST_DATA_PATH_B_outs_29_port, QN => n_1833);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_30_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4129, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196, Q => 
                           DLX_INST_DATA_PATH_B_outs_30_port, QN => n_1834);
   DLX_INST_DATA_PATH_DECODE_RF_OUT2_reg_31_inst : DFF_X1 port map( D => 
                           DLX_INST_DATA_PATH_DECODE_RF_n4130, CK => 
                           DLX_INST_DATA_PATH_DECODE_RF_n5196, Q => 
                           DLX_INST_DATA_PATH_B_outs_31_port, QN => n_1835);
   DLX_INST_DATA_PATH_EXECUTE_U3 : BUF_X1 port map( A => DLX_INST_DATA_PATH_n4,
                           Z => DLX_INST_DATA_PATH_EXECUTE_n4);
   DLX_INST_DATA_PATH_EXECUTE_U2 : BUF_X1 port map( A => DLX_INST_DATA_PATH_n3,
                           Z => DLX_INST_DATA_PATH_EXECUTE_n3);
   DLX_INST_DATA_PATH_EXECUTE_alu1 : alu port map( FUNC(3) => 
                           DLX_INST_ALU_OPCODE_signal_0_port, FUNC(2) => 
                           DLX_INST_ALU_OPCODE_signal_1_port, FUNC(1) => 
                           DLX_INST_ALU_OPCODE_signal_2_port, FUNC(0) => 
                           DLX_INST_ALU_OPCODE_signal_3_port, A(31) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_31_port, A(30) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_30_port, 
                           A(29) => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_29_port
                           , A(28) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_28_port, A(27) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_27_port, 
                           A(26) => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_26_port
                           , A(25) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_25_port, A(24) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_24_port, 
                           A(23) => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_23_port
                           , A(22) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_22_port, A(21) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_21_port, 
                           A(20) => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_20_port
                           , A(19) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_19_port, A(18) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_18_port, 
                           A(17) => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_17_port
                           , A(16) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_16_port, A(15) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_15_port, 
                           A(14) => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_14_port
                           , A(13) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_13_port, A(12) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_12_port, 
                           A(11) => DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_11_port
                           , A(10) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_10_port, A(9) =>
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_9_port, A(8) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_8_port, A(7) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_7_port, A(6) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_6_port, A(5) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_5_port, A(4) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_4_port, A(3) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_3_port, A(2) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_2_port, A(1) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_1_port, A(0) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_0_port, B(31) =>
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_31_port, B(30) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_30_port, 
                           B(29) => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_29_port
                           , B(28) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_28_port, B(27) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_27_port, 
                           B(26) => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_26_port
                           , B(25) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_25_port, B(24) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_24_port, 
                           B(23) => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_23_port
                           , B(22) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_22_port, B(21) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_21_port, 
                           B(20) => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_20_port
                           , B(19) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_19_port, B(18) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_18_port, 
                           B(17) => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_17_port
                           , B(16) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_16_port, B(15) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_15_port, 
                           B(14) => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_14_port
                           , B(13) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_13_port, B(12) 
                           => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_12_port, 
                           B(11) => DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_11_port
                           , B(10) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_10_port, B(9) =>
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_9_port, B(8) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_8_port, B(7) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_7_port, B(6) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_6_port, B(5) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_5_port, B(4) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_4_port, B(3) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_3_port, B(2) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_2_port, B(1) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_1_port, B(0) => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_0_port, 
                           OUTALU(31) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_31_port, 
                           OUTALU(30) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_30_port, 
                           OUTALU(29) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_29_port, 
                           OUTALU(28) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_28_port, 
                           OUTALU(27) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_27_port, 
                           OUTALU(26) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_26_port, 
                           OUTALU(25) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_25_port, 
                           OUTALU(24) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_24_port, 
                           OUTALU(23) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_23_port, 
                           OUTALU(22) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_22_port, 
                           OUTALU(21) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_21_port, 
                           OUTALU(20) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_20_port, 
                           OUTALU(19) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_19_port, 
                           OUTALU(18) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_18_port, 
                           OUTALU(17) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_17_port, 
                           OUTALU(16) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_16_port, 
                           OUTALU(15) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_15_port, 
                           OUTALU(14) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_14_port, 
                           OUTALU(13) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_13_port, 
                           OUTALU(12) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_12_port, 
                           OUTALU(11) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_11_port, 
                           OUTALU(10) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_10_port, 
                           OUTALU(9) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_9_port, 
                           OUTALU(8) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_8_port, 
                           OUTALU(7) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_7_port, 
                           OUTALU(6) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_6_port, 
                           OUTALU(5) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_5_port, 
                           OUTALU(4) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_4_port, 
                           OUTALU(3) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_3_port, 
                           OUTALU(2) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_2_port, 
                           OUTALU(1) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_1_port, 
                           OUTALU(0) => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_0_port);
   DLX_INST_DATA_PATH_EXECUTE_Logic1_port <= '1';
   DLX_INST_DATA_PATH_EXECUTE_zerodec_U11 : NOR4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_A_outs_27_port, A2 => 
                           DLX_INST_DATA_PATH_A_outs_26_port, A3 => 
                           DLX_INST_DATA_PATH_A_outs_25_port, A4 => 
                           DLX_INST_DATA_PATH_A_outs_24_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n17);
   DLX_INST_DATA_PATH_EXECUTE_zerodec_U10 : NOR4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_A_outs_30_port, A2 => 
                           DLX_INST_DATA_PATH_A_outs_2_port, A3 => 
                           DLX_INST_DATA_PATH_A_outs_29_port, A4 => 
                           DLX_INST_DATA_PATH_A_outs_28_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n18);
   DLX_INST_DATA_PATH_EXECUTE_zerodec_U9 : NOR4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_A_outs_5_port, A2 => 
                           DLX_INST_DATA_PATH_A_outs_4_port, A3 => 
                           DLX_INST_DATA_PATH_A_outs_3_port, A4 => 
                           DLX_INST_DATA_PATH_A_outs_31_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n19);
   DLX_INST_DATA_PATH_EXECUTE_zerodec_U8 : NOR4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_A_outs_9_port, A2 => 
                           DLX_INST_DATA_PATH_A_outs_8_port, A3 => 
                           DLX_INST_DATA_PATH_A_outs_7_port, A4 => 
                           DLX_INST_DATA_PATH_A_outs_6_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n20);
   DLX_INST_DATA_PATH_EXECUTE_zerodec_U7 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n17, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n18, A3 => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n19, A4 => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n20, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n11);
   DLX_INST_DATA_PATH_EXECUTE_zerodec_U6 : NOR4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_A_outs_12_port, A2 => 
                           DLX_INST_DATA_PATH_A_outs_11_port, A3 => 
                           DLX_INST_DATA_PATH_A_outs_10_port, A4 => 
                           DLX_INST_DATA_PATH_A_outs_0_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n13);
   DLX_INST_DATA_PATH_EXECUTE_zerodec_U5 : NOR4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_A_outs_16_port, A2 => 
                           DLX_INST_DATA_PATH_A_outs_15_port, A3 => 
                           DLX_INST_DATA_PATH_A_outs_14_port, A4 => 
                           DLX_INST_DATA_PATH_A_outs_13_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n14);
   DLX_INST_DATA_PATH_EXECUTE_zerodec_U4 : NOR4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_A_outs_1_port, A2 => 
                           DLX_INST_DATA_PATH_A_outs_19_port, A3 => 
                           DLX_INST_DATA_PATH_A_outs_18_port, A4 => 
                           DLX_INST_DATA_PATH_A_outs_17_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n15);
   DLX_INST_DATA_PATH_EXECUTE_zerodec_U3 : NOR4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_A_outs_23_port, A2 => 
                           DLX_INST_DATA_PATH_A_outs_22_port, A3 => 
                           DLX_INST_DATA_PATH_A_outs_21_port, A4 => 
                           DLX_INST_DATA_PATH_A_outs_20_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n16);
   DLX_INST_DATA_PATH_EXECUTE_zerodec_U2 : NAND4_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n13, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n14, A3 => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n15, A4 => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n16, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n12);
   DLX_INST_DATA_PATH_EXECUTE_zerodec_U1 : NOR2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_zerodec_n12, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ZERO_DEC_OUT);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U32 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_0_port, B => 
                           DLX_INST_DATA_PATH_A_outs_0_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_0_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U31 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_10_port, B => 
                           DLX_INST_DATA_PATH_A_outs_10_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_10_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U30 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_11_port, B => 
                           DLX_INST_DATA_PATH_A_outs_11_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_11_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U29 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_12_port, B => 
                           DLX_INST_DATA_PATH_A_outs_12_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_12_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U28 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_13_port, B => 
                           DLX_INST_DATA_PATH_A_outs_13_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_13_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U27 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_14_port, B => 
                           DLX_INST_DATA_PATH_A_outs_14_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_14_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U26 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_15_port, B => 
                           DLX_INST_DATA_PATH_A_outs_15_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_15_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U25 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_16_port, B => 
                           DLX_INST_DATA_PATH_A_outs_16_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_16_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U24 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_17_port, B => 
                           DLX_INST_DATA_PATH_A_outs_17_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_17_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U23 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_18_port, B => 
                           DLX_INST_DATA_PATH_A_outs_18_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_18_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U22 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_19_port, B => 
                           DLX_INST_DATA_PATH_A_outs_19_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_19_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U21 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_1_port, B => 
                           DLX_INST_DATA_PATH_A_outs_1_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_1_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U20 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_20_port, B => 
                           DLX_INST_DATA_PATH_A_outs_20_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_20_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U19 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_21_port, B => 
                           DLX_INST_DATA_PATH_A_outs_21_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_21_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U18 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_22_port, B => 
                           DLX_INST_DATA_PATH_A_outs_22_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_22_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U17 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_23_port, B => 
                           DLX_INST_DATA_PATH_A_outs_23_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_23_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U16 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_24_port, B => 
                           DLX_INST_DATA_PATH_A_outs_24_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_24_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U15 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_25_port, B => 
                           DLX_INST_DATA_PATH_A_outs_25_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_25_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U14 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_26_port, B => 
                           DLX_INST_DATA_PATH_A_outs_26_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_26_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U13 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_27_port, B => 
                           DLX_INST_DATA_PATH_A_outs_27_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_27_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U12 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_28_port, B => 
                           DLX_INST_DATA_PATH_A_outs_28_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_28_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U11 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_29_port, B => 
                           DLX_INST_DATA_PATH_A_outs_29_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_29_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U10 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_2_port, B => 
                           DLX_INST_DATA_PATH_A_outs_2_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_2_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U9 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_30_port, B => 
                           DLX_INST_DATA_PATH_A_outs_30_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_30_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U8 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_31_port, B => 
                           DLX_INST_DATA_PATH_A_outs_31_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_31_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U7 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_3_port, B => 
                           DLX_INST_DATA_PATH_A_outs_3_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_3_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U6 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_4_port, B => 
                           DLX_INST_DATA_PATH_A_outs_4_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_4_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U5 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_5_port, B => 
                           DLX_INST_DATA_PATH_A_outs_5_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_5_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U4 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_6_port, B => 
                           DLX_INST_DATA_PATH_A_outs_6_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_6_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_7_port, B => 
                           DLX_INST_DATA_PATH_A_outs_7_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_7_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U2 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_8_port, B => 
                           DLX_INST_DATA_PATH_A_outs_8_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_8_port);
   DLX_INST_DATA_PATH_EXECUTE_mux1_U1 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_NPC2_OUTs_9_port, B => 
                           DLX_INST_DATA_PATH_A_outs_9_port, S => 
                           DLX_INST_MUXA_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX1_OUT_9_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U32 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_0_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_0_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_0_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U31 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_10_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_10_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_10_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U30 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_11_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_11_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_11_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U29 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_12_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_12_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_12_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U28 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_13_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_13_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_13_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U27 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_14_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_14_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_14_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U26 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_15_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_15_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_15_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U25 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_16_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_16_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_16_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U24 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_17_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_17_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_17_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U23 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_18_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_18_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_18_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U22 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_19_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_19_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_19_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U21 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_1_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_1_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_1_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U20 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_20_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_20_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_20_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U19 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_21_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_21_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_21_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U18 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_22_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_22_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_22_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U17 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_23_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_23_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_23_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U16 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_24_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_24_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_24_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U15 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_25_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_25_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_25_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U14 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_26_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_26_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_26_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U13 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_27_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_27_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_27_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U12 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_28_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_28_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_28_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U11 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_29_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_29_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_29_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U10 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_2_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_2_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_2_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U9 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_30_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_30_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_30_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U8 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_31_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_31_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_31_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U7 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_3_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_3_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_3_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U6 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_4_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_4_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_4_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U5 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_5_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_5_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_5_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U4 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_6_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_6_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_6_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_7_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_7_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_7_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U2 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_8_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_8_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_8_port);
   DLX_INST_DATA_PATH_EXECUTE_mux2_U1 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_B_outs_9_port, B => 
                           DLX_INST_DATA_PATH_Imm_outs_9_port, S => 
                           DLX_INST_MUXB_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_MUX2_OUT_9_port);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_U8 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n16, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_U7 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n16, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_U6 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n16, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_U5 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n12, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n11);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_U4 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n12, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_U3 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n12, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_U2 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_n4, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n16);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_U1 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_n3, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n12);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_0_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_0_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_0_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_0_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_0_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_0_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_0_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_0_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_0_n2, Q => 
                           ADDRESS_DRAM_signal_0_port, QN => n_1836);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_1_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_1_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_1_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_1_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_1_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_1_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_1_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_1_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_1_n2, Q => 
                           ADDRESS_DRAM_signal_1_port, QN => n_1837);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_2_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_2_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_2_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_2_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_2_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_2_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_2_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_2_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_2_n2, Q => 
                           ADDRESS_DRAM_signal_2_port, QN => n_1838);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_3_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_3_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_3_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_3_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_3_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_3_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_3_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_3_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_3_n2, Q => 
                           ADDRESS_DRAM_signal_3_port, QN => n_1839);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_4_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_4_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_4_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_4_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_4_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_4_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_4_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_4_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_4_n2, Q => 
                           ADDRESS_DRAM_signal_4_port, QN => n_1840);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_5_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_5_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_5_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_5_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_5_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_5_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_5_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_5_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_5_n2, Q => 
                           ADDRESS_DRAM_signal_5_port, QN => n_1841);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_6_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_6_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_6_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_6_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_6_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_6_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_6_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_6_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_6_n2, Q => 
                           ADDRESS_DRAM_signal_6_port, QN => n_1842);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_7_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_7_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_7_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_7_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_7_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_7_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_7_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_7_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_7_n2, Q => 
                           ADDRESS_DRAM_signal_7_port, QN => n_1843);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_8_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_8_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_8_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_8_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_8_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_8_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_8_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_8_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_8_n2, Q => 
                           ADDRESS_DRAM_signal_8_port, QN => n_1844);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_9_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_9_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_9_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_9_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_9_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_9_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_9_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_9_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_9_n2, Q => 
                           ADDRESS_DRAM_signal_9_port, QN => n_1845);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_10_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_10_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_10_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_10_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_10_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_10_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_10_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_10_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_10_n2, Q => 
                           ADDRESS_DRAM_signal_10_port, QN => n_1846);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_11_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_11_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_11_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_11_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_11_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n9, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_11_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_11_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_11_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_11_n2, Q => 
                           ADDRESS_DRAM_signal_11_port, QN => n_1847);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_12_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_12_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_12_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_12_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_12_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_12_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_12_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_12_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_12_n2, Q => 
                           ADDRESS_DRAM_signal_12_port, QN => n_1848);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_13_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_13_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_13_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_13_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_13_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_13_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_13_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_13_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_13_n2, Q => 
                           ADDRESS_DRAM_signal_13_port, QN => n_1849);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_14_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_14_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_14_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_14_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_14_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_14_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_14_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_14_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_14_n2, Q => 
                           ADDRESS_DRAM_signal_14_port, QN => n_1850);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_15_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_15_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_15_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_15_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_15_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_15_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_15_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_15_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_15_n2, Q => 
                           ADDRESS_DRAM_signal_15_port, QN => n_1851);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_16_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_16_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_16_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_16_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_16_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_16_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_16_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_16_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_16_n2, Q => 
                           ADDRESS_DRAM_signal_16_port, QN => n_1852);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_17_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_17_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_17_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_17_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_17_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_17_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_17_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_17_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_17_n2, Q => 
                           ADDRESS_DRAM_signal_17_port, QN => n_1853);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_18_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_18_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_18_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_18_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_18_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_18_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_18_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_18_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_18_n2, Q => 
                           ADDRESS_DRAM_signal_18_port, QN => n_1854);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_19_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_19_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_19_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_19_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_19_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_19_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_19_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_19_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_19_n2, Q => 
                           ADDRESS_DRAM_signal_19_port, QN => n_1855);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_20_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_20_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_20_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_20_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_20_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_20_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_20_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_20_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_20_n2, Q => 
                           ADDRESS_DRAM_signal_20_port, QN => n_1856);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_21_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_21_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_21_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_21_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_21_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_21_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_21_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_21_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_21_n2, Q => 
                           ADDRESS_DRAM_signal_21_port, QN => n_1857);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_22_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_22_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_22_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_22_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_22_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_22_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_22_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_22_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_22_n2, Q => 
                           ADDRESS_DRAM_signal_22_port, QN => n_1858);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_23_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_23_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_23_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_23_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_23_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n10, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_23_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_23_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_23_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_23_n2, Q => 
                           ADDRESS_DRAM_signal_23_port, QN => n_1859);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_24_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_24_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_24_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_24_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_24_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n11, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_24_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_24_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_24_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_24_n2, Q => 
                           ADDRESS_DRAM_signal_24_port, QN => n_1860);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_25_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_25_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_25_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_25_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_25_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n11, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_25_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_25_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_25_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_25_n2, Q => 
                           ADDRESS_DRAM_signal_25_port, QN => n_1861);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_26_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_26_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_26_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_26_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_26_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n11, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_26_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_26_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_26_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_26_n2, Q => 
                           ADDRESS_DRAM_signal_26_port, QN => n_1862);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_27_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_27_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_27_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_27_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_27_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n11, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_27_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_27_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_27_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_27_n2, Q => 
                           ADDRESS_DRAM_signal_27_port, QN => n_1863);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_28_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_28_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_28_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_28_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_28_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n11, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_28_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_28_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_28_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_28_n2, Q => 
                           ADDRESS_DRAM_signal_28_port, QN => n_1864);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_29_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_29_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_29_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_29_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_29_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n11, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_29_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_29_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_29_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_29_n2, Q => 
                           ADDRESS_DRAM_signal_29_port, QN => n_1865);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_30_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_30_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_30_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_30_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_30_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n11, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_30_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_30_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_30_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_30_n2, Q => 
                           ADDRESS_DRAM_signal_30_port, QN => n_1866);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_31_U3 : MUX2_X1 port map( A => 
                           ADDRESS_DRAM_signal_31_port, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ALU_output_31_port, S => 
                           DLX_INST_ALU_OUTREG_EN_signal, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_31_n1);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_31_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n11, A2 => 
                           DLX_INST_ALU_OUTREG_EN_signal, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_31_n2);
   DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_31_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_31_n1, CK =>
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_ALUoutput_FF_31_n2, Q => 
                           ADDRESS_DRAM_signal_31_port, QN => n_1867);
   DLX_INST_DATA_PATH_EXECUTE_IR3_U8 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n16, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n15);
   DLX_INST_DATA_PATH_EXECUTE_IR3_U7 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n16, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14);
   DLX_INST_DATA_PATH_EXECUTE_IR3_U6 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n16, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13);
   DLX_INST_DATA_PATH_EXECUTE_IR3_U5 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n12, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n11);
   DLX_INST_DATA_PATH_EXECUTE_IR3_U4 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n12, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10);
   DLX_INST_DATA_PATH_EXECUTE_IR3_U3 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n12, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9);
   DLX_INST_DATA_PATH_EXECUTE_IR3_U2 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_n4, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n16);
   DLX_INST_DATA_PATH_EXECUTE_IR3_U1 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_n3, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n12);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_0_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_0_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_0_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_0_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_0_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_0_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_0_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_0_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_0_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_0_port, QN => n_1868);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_1_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_1_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_1_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_1_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_1_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_1_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_1_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_1_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_1_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_1_port, QN => n_1869);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_2_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_2_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_2_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_2_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_2_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_2_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_2_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_2_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_2_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_2_port, QN => n_1870);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_3_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_3_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_3_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_3_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_3_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_3_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_3_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_3_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_3_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_3_port, QN => n_1871);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_4_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_4_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_4_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_4_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_4_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_4_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_4_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_4_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_4_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_4_port, QN => n_1872);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_5_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_5_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_5_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_5_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_5_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_5_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_5_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_5_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_5_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_5_port, QN => n_1873);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_6_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_6_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_6_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_6_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_6_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_6_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_6_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_6_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_6_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_6_port, QN => n_1874);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_7_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_7_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_7_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_7_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_7_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_7_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_7_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_7_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_7_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_7_port, QN => n_1875);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_8_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_8_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_8_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_8_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_8_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_8_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_8_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_8_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_8_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_8_port, QN => n_1876);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_9_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_9_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_9_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_9_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_9_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_9_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_9_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_9_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_9_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_9_port, QN => n_1877);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_10_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_10_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_10_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_10_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_10_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_10_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_10_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_10_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n13, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_10_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_10_port, QN => n_1878);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_11_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_11_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_11_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_11_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_11_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_11_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_11_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_11_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_11_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_11_port, QN => n_1879);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_12_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_12_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_12_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_12_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_12_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_12_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_12_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_12_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_12_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_12_port, QN => n_1880);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_13_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_13_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_13_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_13_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_13_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_13_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_13_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_13_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_13_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_13_port, QN => n_1881);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_14_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_14_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_14_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_14_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_14_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_14_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_14_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_14_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_14_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_14_port, QN => n_1882);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_15_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_15_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_15_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_15_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_15_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_15_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_15_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_15_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_15_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_15_port, QN => n_1883);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_16_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_16_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_16_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_16_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_16_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_16_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_16_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_16_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_16_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_16_port, QN => n_1884);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_17_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_17_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_17_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_17_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_17_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_17_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_17_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_17_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_17_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_17_port, QN => n_1885);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_18_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_18_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_18_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_18_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_18_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_18_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_18_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_18_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_18_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_18_port, QN => n_1886);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_19_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_19_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_19_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_19_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_19_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_19_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_19_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_19_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_19_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_19_port, QN => n_1887);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_20_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_20_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_20_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_20_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_20_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_20_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_20_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_20_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_20_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_20_port, QN => n_1888);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_21_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_21_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_21_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_21_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_21_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_21_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_21_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_21_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n14, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_21_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_21_port, QN => n_1889);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_22_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_22_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_22_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_22_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_22_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_22_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_22_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_22_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_22_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_22_port, QN => n_1890);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_23_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_23_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_23_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_23_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_23_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_23_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_23_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_23_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_23_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_23_port, QN => n_1891);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_24_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_24_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_24_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_24_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_24_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_24_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_24_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_24_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_24_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_24_port, QN => n_1892);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_25_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_25_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_25_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_25_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_25_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_25_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_25_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_25_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_25_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_25_port, QN => n_1893);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_26_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_26_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_26_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_26_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_26_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_26_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_26_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_26_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_26_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_26_port, QN => n_1894);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_27_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_27_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_27_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_27_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_27_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_27_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_27_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_27_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_27_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_27_port, QN => n_1895);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_28_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_28_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_28_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_28_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_28_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_28_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_28_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_28_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_28_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_28_port, QN => n_1896);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_29_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_29_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_29_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_29_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_29_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_29_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_29_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_29_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_29_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_29_port, QN => n_1897);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_30_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_30_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_30_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_30_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_30_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_30_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_30_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_30_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_30_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_30_port, QN => n_1898);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_31_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT3s_31_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT2s_31_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_31_n1);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_31_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_31_n2);
   DLX_INST_DATA_PATH_EXECUTE_IR3_FF_31_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_31_n1, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_n15, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_IR3_FF_31_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT3s_31_port, QN => n_1899);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_U8 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n16, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_U7 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n16, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_U6 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n16, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_U5 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n12, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n11);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_U4 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n12, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_U3 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n12, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_U2 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_n4, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n16);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_U1 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_EXECUTE_n3, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n12);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_0_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_0_port, B => 
                           DLX_INST_DATA_PATH_B_outs_0_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_0_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_0_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_0_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_0_Q_reg : DFFR_X1 port map( D =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_0_n1, CK
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13, RN 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_0_n2,
                           Q => DATAwrite_DRAM_signal_0_port, QN => n_1900);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_1_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_1_port, B => 
                           DLX_INST_DATA_PATH_B_outs_1_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_1_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_1_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_1_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_1_Q_reg : DFFR_X1 port map( D =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_1_n1, CK
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13, RN 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_1_n2,
                           Q => DATAwrite_DRAM_signal_1_port, QN => n_1901);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_2_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_2_port, B => 
                           DLX_INST_DATA_PATH_B_outs_2_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_2_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_2_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_2_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_2_Q_reg : DFFR_X1 port map( D =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_2_n1, CK
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13, RN 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_2_n2,
                           Q => DATAwrite_DRAM_signal_2_port, QN => n_1902);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_3_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_3_port, B => 
                           DLX_INST_DATA_PATH_B_outs_3_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_3_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_3_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_3_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_3_Q_reg : DFFR_X1 port map( D =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_3_n1, CK
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13, RN 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_3_n2,
                           Q => DATAwrite_DRAM_signal_3_port, QN => n_1903);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_4_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_4_port, B => 
                           DLX_INST_DATA_PATH_B_outs_4_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_4_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_4_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_4_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_4_Q_reg : DFFR_X1 port map( D =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_4_n1, CK
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13, RN 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_4_n2,
                           Q => DATAwrite_DRAM_signal_4_port, QN => n_1904);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_5_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_5_port, B => 
                           DLX_INST_DATA_PATH_B_outs_5_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_5_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_5_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_5_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_5_Q_reg : DFFR_X1 port map( D =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_5_n1, CK
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13, RN 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_5_n2,
                           Q => DATAwrite_DRAM_signal_5_port, QN => n_1905);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_6_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_6_port, B => 
                           DLX_INST_DATA_PATH_B_outs_6_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_6_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_6_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_6_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_6_Q_reg : DFFR_X1 port map( D =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_6_n1, CK
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13, RN 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_6_n2,
                           Q => DATAwrite_DRAM_signal_6_port, QN => n_1906);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_7_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_7_port, B => 
                           DLX_INST_DATA_PATH_B_outs_7_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_7_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_7_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_7_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_7_Q_reg : DFFR_X1 port map( D =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_7_n1, CK
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13, RN 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_7_n2,
                           Q => DATAwrite_DRAM_signal_7_port, QN => n_1907);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_8_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_8_port, B => 
                           DLX_INST_DATA_PATH_B_outs_8_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_8_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_8_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_8_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_8_Q_reg : DFFR_X1 port map( D =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_8_n1, CK
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13, RN 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_8_n2,
                           Q => DATAwrite_DRAM_signal_8_port, QN => n_1908);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_9_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_9_port, B => 
                           DLX_INST_DATA_PATH_B_outs_9_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_9_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_9_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_9_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_9_Q_reg : DFFR_X1 port map( D =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_9_n1, CK
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13, RN 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_9_n2,
                           Q => DATAwrite_DRAM_signal_9_port, QN => n_1909);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_10_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_10_port, B => 
                           DLX_INST_DATA_PATH_B_outs_10_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_10_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_10_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_10_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_10_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_10_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n13
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_10_n2, Q
                           => DATAwrite_DRAM_signal_10_port, QN => n_1910);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_11_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_11_port, B => 
                           DLX_INST_DATA_PATH_B_outs_11_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_11_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_11_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n9, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_11_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_11_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_11_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_11_n2, Q
                           => DATAwrite_DRAM_signal_11_port, QN => n_1911);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_12_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_12_port, B => 
                           DLX_INST_DATA_PATH_B_outs_12_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_12_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_12_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_12_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_12_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_12_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_12_n2, Q
                           => DATAwrite_DRAM_signal_12_port, QN => n_1912);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_13_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_13_port, B => 
                           DLX_INST_DATA_PATH_B_outs_13_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_13_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_13_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_13_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_13_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_13_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_13_n2, Q
                           => DATAwrite_DRAM_signal_13_port, QN => n_1913);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_14_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_14_port, B => 
                           DLX_INST_DATA_PATH_B_outs_14_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_14_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_14_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_14_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_14_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_14_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_14_n2, Q
                           => DATAwrite_DRAM_signal_14_port, QN => n_1914);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_15_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_15_port, B => 
                           DLX_INST_DATA_PATH_B_outs_15_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_15_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_15_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_15_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_15_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_15_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_15_n2, Q
                           => DATAwrite_DRAM_signal_15_port, QN => n_1915);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_16_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_16_port, B => 
                           DLX_INST_DATA_PATH_B_outs_16_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_16_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_16_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_16_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_16_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_16_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_16_n2, Q
                           => DATAwrite_DRAM_signal_16_port, QN => n_1916);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_17_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_17_port, B => 
                           DLX_INST_DATA_PATH_B_outs_17_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_17_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_17_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_17_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_17_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_17_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_17_n2, Q
                           => DATAwrite_DRAM_signal_17_port, QN => n_1917);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_18_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_18_port, B => 
                           DLX_INST_DATA_PATH_B_outs_18_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_18_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_18_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_18_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_18_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_18_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_18_n2, Q
                           => DATAwrite_DRAM_signal_18_port, QN => n_1918);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_19_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_19_port, B => 
                           DLX_INST_DATA_PATH_B_outs_19_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_19_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_19_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_19_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_19_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_19_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_19_n2, Q
                           => DATAwrite_DRAM_signal_19_port, QN => n_1919);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_20_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_20_port, B => 
                           DLX_INST_DATA_PATH_B_outs_20_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_20_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_20_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_20_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_20_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_20_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_20_n2, Q
                           => DATAwrite_DRAM_signal_20_port, QN => n_1920);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_21_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_21_port, B => 
                           DLX_INST_DATA_PATH_B_outs_21_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_21_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_21_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_21_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_21_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_21_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n14
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_21_n2, Q
                           => DATAwrite_DRAM_signal_21_port, QN => n_1921);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_22_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_22_port, B => 
                           DLX_INST_DATA_PATH_B_outs_22_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_22_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_22_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_22_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_22_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_22_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_22_n2, Q
                           => DATAwrite_DRAM_signal_22_port, QN => n_1922);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_23_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_23_port, B => 
                           DLX_INST_DATA_PATH_B_outs_23_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_23_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_23_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n10, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_23_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_23_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_23_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_23_n2, Q
                           => DATAwrite_DRAM_signal_23_port, QN => n_1923);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_24_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_24_port, B => 
                           DLX_INST_DATA_PATH_B_outs_24_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_24_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_24_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_24_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_24_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_24_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_24_n2, Q
                           => DATAwrite_DRAM_signal_24_port, QN => n_1924);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_25_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_25_port, B => 
                           DLX_INST_DATA_PATH_B_outs_25_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_25_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_25_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_25_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_25_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_25_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_25_n2, Q
                           => DATAwrite_DRAM_signal_25_port, QN => n_1925);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_26_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_26_port, B => 
                           DLX_INST_DATA_PATH_B_outs_26_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_26_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_26_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_26_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_26_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_26_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_26_n2, Q
                           => DATAwrite_DRAM_signal_26_port, QN => n_1926);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_27_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_27_port, B => 
                           DLX_INST_DATA_PATH_B_outs_27_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_27_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_27_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_27_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_27_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_27_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_27_n2, Q
                           => DATAwrite_DRAM_signal_27_port, QN => n_1927);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_28_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_28_port, B => 
                           DLX_INST_DATA_PATH_B_outs_28_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_28_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_28_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_28_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_28_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_28_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_28_n2, Q
                           => DATAwrite_DRAM_signal_28_port, QN => n_1928);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_29_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_29_port, B => 
                           DLX_INST_DATA_PATH_B_outs_29_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_29_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_29_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_29_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_29_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_29_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_29_n2, Q
                           => DATAwrite_DRAM_signal_29_port, QN => n_1929);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_30_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_30_port, B => 
                           DLX_INST_DATA_PATH_B_outs_30_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_30_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_30_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_30_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_30_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_30_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_30_n2, Q
                           => DATAwrite_DRAM_signal_30_port, QN => n_1930);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_31_U3 : MUX2_X1 port map( A => 
                           DATAwrite_DRAM_signal_31_port, B => 
                           DLX_INST_DATA_PATH_B_outs_31_port, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_31_n1);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_31_U2 : NAND2_X1 port map( A1 =>
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_n11, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_31_n2);
   DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_31_Q_reg : DFFR_X1 port map( D 
                           => DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_31_n1
                           , CK => DLX_INST_DATA_PATH_EXECUTE_B_outregister_n15
                           , RN => 
                           DLX_INST_DATA_PATH_EXECUTE_B_outregister_FF_31_n2, Q
                           => DATAwrite_DRAM_signal_31_port, QN => n_1931);
   DLX_INST_DATA_PATH_EXECUTE_XNOR_2_U1 : XNOR2_X1 port map( A => 
                           DLX_INST_EQ_COND_signal, B => 
                           DLX_INST_DATA_PATH_EXECUTE_ZERO_DEC_OUT, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_XNOR_OUT);
   DLX_INST_DATA_PATH_EXECUTE_COND_U3 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_EXECUTE_n3, A2 => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_EXECUTE_COND_n3);
   DLX_INST_DATA_PATH_EXECUTE_COND_U2 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_COND_OUTs, B => 
                           DLX_INST_DATA_PATH_EXECUTE_XNOR_OUT, S => 
                           DLX_INST_DATA_PATH_EXECUTE_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_EXECUTE_COND_n4);
   DLX_INST_DATA_PATH_EXECUTE_COND_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_EXECUTE_COND_n4, CK => 
                           DLX_INST_DATA_PATH_EXECUTE_n4, RN => 
                           DLX_INST_DATA_PATH_EXECUTE_COND_n3, Q => 
                           DLX_INST_DATA_PATH_COND_OUTs, QN => n_1932);
   DLX_INST_DATA_PATH_MEMORY_U4 : BUF_X1 port map( A => DLX_INST_DATA_PATH_n4, 
                           Z => DLX_INST_DATA_PATH_MEMORY_n4);
   DLX_INST_DATA_PATH_MEMORY_U3 : BUF_X1 port map( A => DLX_INST_DATA_PATH_n3, 
                           Z => DLX_INST_DATA_PATH_MEMORY_n3);
   DLX_INST_DATA_PATH_MEMORY_Logic0_port <= '0';
   DLX_INST_DATA_PATH_MEMORY_Logic1_port <= '1';
   DLX_INST_DATA_PATH_MEMORY_JUMPMUX_U1 : MUX2_X2 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_Logic0_port, B => 
                           DLX_INST_DATA_PATH_COND_OUTs, S => 
                           DLX_INST_JUMP_EN_signal, Z => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U32 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_0_port, B => 
                           ADDRESS_DRAM_signal_0_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_0_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U31 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_10_port, B => 
                           ADDRESS_DRAM_signal_10_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_10_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U30 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_11_port, B => 
                           ADDRESS_DRAM_signal_11_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_11_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U29 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_12_port, B => 
                           ADDRESS_DRAM_signal_12_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_12_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U28 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_13_port, B => 
                           ADDRESS_DRAM_signal_13_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_13_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U27 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_14_port, B => 
                           ADDRESS_DRAM_signal_14_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_14_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U26 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_15_port, B => 
                           ADDRESS_DRAM_signal_15_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_15_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U25 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_16_port, B => 
                           ADDRESS_DRAM_signal_16_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_16_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U24 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_17_port, B => 
                           ADDRESS_DRAM_signal_17_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_17_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U23 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_18_port, B => 
                           ADDRESS_DRAM_signal_18_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_18_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U22 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_19_port, B => 
                           ADDRESS_DRAM_signal_19_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_19_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U21 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_1_port, B => 
                           ADDRESS_DRAM_signal_1_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_1_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U20 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_20_port, B => 
                           ADDRESS_DRAM_signal_20_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_20_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U19 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_21_port, B => 
                           ADDRESS_DRAM_signal_21_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_21_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U18 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_22_port, B => 
                           ADDRESS_DRAM_signal_22_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_22_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U17 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_23_port, B => 
                           ADDRESS_DRAM_signal_23_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_23_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U16 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_24_port, B => 
                           ADDRESS_DRAM_signal_24_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_24_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U15 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_25_port, B => 
                           ADDRESS_DRAM_signal_25_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_25_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U14 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_26_port, B => 
                           ADDRESS_DRAM_signal_26_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_26_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U13 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_27_port, B => 
                           ADDRESS_DRAM_signal_27_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_27_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U12 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_28_port, B => 
                           ADDRESS_DRAM_signal_28_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_28_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U11 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_29_port, B => 
                           ADDRESS_DRAM_signal_29_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_29_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U10 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_2_port, B => 
                           ADDRESS_DRAM_signal_2_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_2_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U9 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_30_port, B => 
                           ADDRESS_DRAM_signal_30_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_30_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U8 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_31_port, B => 
                           ADDRESS_DRAM_signal_31_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_31_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U7 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_3_port, B => 
                           ADDRESS_DRAM_signal_3_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_3_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U6 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_4_port, B => 
                           ADDRESS_DRAM_signal_4_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_4_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U5 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_5_port, B => 
                           ADDRESS_DRAM_signal_5_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_5_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U4 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_6_port, B => 
                           ADDRESS_DRAM_signal_6_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_6_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_7_port, B => 
                           ADDRESS_DRAM_signal_7_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_7_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U2 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_8_port, B => 
                           ADDRESS_DRAM_signal_8_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_8_port);
   DLX_INST_DATA_PATH_MEMORY_MUX_PC_U1 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ADDERPC_OUTs_9_port, B => 
                           ADDRESS_DRAM_signal_9_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_muxjmp_to_mux, Z => 
                           DLX_INST_DATA_PATH_TO_PC_OUTs_9_port);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_U8 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n16, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_U7 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n16, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_U6 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n16, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_U5 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n12, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n11);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_U4 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n12, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_U3 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n12, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_U2 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_n4, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n16);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_U1 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_n3, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n12);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_0_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_0_port, B => 
                           ADDRESS_DRAM_signal_0_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_0_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_0_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_0_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_0_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_0_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_0_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_0_port, QN => n_1933);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_1_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_1_port, B => 
                           ADDRESS_DRAM_signal_1_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_1_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_1_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_1_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_1_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_1_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_1_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_1_port, QN => n_1934);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_2_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_2_port, B => 
                           ADDRESS_DRAM_signal_2_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_2_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_2_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_2_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_2_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_2_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_2_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_2_port, QN => n_1935);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_3_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_3_port, B => 
                           ADDRESS_DRAM_signal_3_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_3_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_3_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_3_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_3_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_3_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_3_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_3_port, QN => n_1936);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_4_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_4_port, B => 
                           ADDRESS_DRAM_signal_4_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_4_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_4_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_4_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_4_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_4_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_4_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_4_port, QN => n_1937);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_5_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_5_port, B => 
                           ADDRESS_DRAM_signal_5_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_5_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_5_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_5_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_5_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_5_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_5_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_5_port, QN => n_1938);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_6_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_6_port, B => 
                           ADDRESS_DRAM_signal_6_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_6_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_6_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_6_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_6_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_6_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_6_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_6_port, QN => n_1939);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_7_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_7_port, B => 
                           ADDRESS_DRAM_signal_7_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_7_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_7_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_7_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_7_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_7_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_7_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_7_port, QN => n_1940);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_8_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_8_port, B => 
                           ADDRESS_DRAM_signal_8_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_8_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_8_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_8_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_8_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_8_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_8_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_8_port, QN => n_1941);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_9_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_9_port, B => 
                           ADDRESS_DRAM_signal_9_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_9_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_9_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_9_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_9_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_9_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_9_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_9_port, QN => n_1942);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_10_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_10_port, B => 
                           ADDRESS_DRAM_signal_10_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_10_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_10_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_10_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_10_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_10_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_10_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_10_port, QN => n_1943);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_11_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_11_port, B => 
                           ADDRESS_DRAM_signal_11_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_11_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_11_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_11_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_11_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_11_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_11_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_11_port, QN => n_1944);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_12_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_12_port, B => 
                           ADDRESS_DRAM_signal_12_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_12_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_12_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_12_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_12_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_12_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_12_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_12_port, QN => n_1945);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_13_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_13_port, B => 
                           ADDRESS_DRAM_signal_13_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_13_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_13_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_13_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_13_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_13_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_13_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_13_port, QN => n_1946);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_14_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_14_port, B => 
                           ADDRESS_DRAM_signal_14_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_14_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_14_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_14_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_14_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_14_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_14_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_14_port, QN => n_1947);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_15_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_15_port, B => 
                           ADDRESS_DRAM_signal_15_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_15_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_15_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_15_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_15_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_15_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_15_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_15_port, QN => n_1948);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_16_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_16_port, B => 
                           ADDRESS_DRAM_signal_16_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_16_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_16_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_16_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_16_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_16_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_16_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_16_port, QN => n_1949);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_17_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_17_port, B => 
                           ADDRESS_DRAM_signal_17_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_17_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_17_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_17_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_17_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_17_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_17_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_17_port, QN => n_1950);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_18_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_18_port, B => 
                           ADDRESS_DRAM_signal_18_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_18_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_18_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_18_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_18_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_18_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_18_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_18_port, QN => n_1951);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_19_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_19_port, B => 
                           ADDRESS_DRAM_signal_19_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_19_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_19_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_19_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_19_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_19_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_19_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_19_port, QN => n_1952);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_20_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_20_port, B => 
                           ADDRESS_DRAM_signal_20_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_20_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_20_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_20_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_20_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_20_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_20_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_20_port, QN => n_1953);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_21_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_21_port, B => 
                           ADDRESS_DRAM_signal_21_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_21_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_21_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_21_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_21_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_21_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_21_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_21_port, QN => n_1954);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_22_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_22_port, B => 
                           ADDRESS_DRAM_signal_22_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_22_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_22_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_22_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_22_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_22_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_22_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_22_port, QN => n_1955);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_23_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_23_port, B => 
                           ADDRESS_DRAM_signal_23_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_23_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_23_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_23_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_23_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_23_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_23_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_23_port, QN => n_1956);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_24_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_24_port, B => 
                           ADDRESS_DRAM_signal_24_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_24_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_24_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_24_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_24_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_24_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_24_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_24_port, QN => n_1957);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_25_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_25_port, B => 
                           ADDRESS_DRAM_signal_25_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_25_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_25_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_25_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_25_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_25_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_25_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_25_port, QN => n_1958);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_26_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_26_port, B => 
                           ADDRESS_DRAM_signal_26_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_26_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_26_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_26_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_26_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_26_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_26_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_26_port, QN => n_1959);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_27_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_27_port, B => 
                           ADDRESS_DRAM_signal_27_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_27_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_27_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_27_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_27_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_27_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_27_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_27_port, QN => n_1960);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_28_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_28_port, B => 
                           ADDRESS_DRAM_signal_28_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_28_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_28_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_28_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_28_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_28_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_28_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_28_port, QN => n_1961);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_29_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_29_port, B => 
                           ADDRESS_DRAM_signal_29_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_29_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_29_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_29_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_29_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_29_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_29_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_29_port, QN => n_1962);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_30_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_30_port, B => 
                           ADDRESS_DRAM_signal_30_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_30_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_30_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_30_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_30_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_30_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_30_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_30_port, QN => n_1963);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_31_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_31_port, B => 
                           ADDRESS_DRAM_signal_31_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_31_n1);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_31_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_31_n2);
   DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_31_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_31_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_ALU_OUT2r_FF_31_n2, Q => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_31_port, QN => n_1964);
   DLX_INST_DATA_PATH_MEMORY_IR4_U8 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n16, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n15);
   DLX_INST_DATA_PATH_MEMORY_IR4_U7 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n16, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14);
   DLX_INST_DATA_PATH_MEMORY_IR4_U6 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n16, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13);
   DLX_INST_DATA_PATH_MEMORY_IR4_U5 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n12, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n11);
   DLX_INST_DATA_PATH_MEMORY_IR4_U4 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n12, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10);
   DLX_INST_DATA_PATH_MEMORY_IR4_U3 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n12, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9);
   DLX_INST_DATA_PATH_MEMORY_IR4_U2 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_n4, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n16);
   DLX_INST_DATA_PATH_MEMORY_IR4_U1 : BUF_X1 port map( A => 
                           DLX_INST_DATA_PATH_MEMORY_n3, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n12);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_0_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_0_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_0_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_0_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_0_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_0_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_0_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_0_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_0_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_0_port, QN => n_1965);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_1_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_1_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_1_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_1_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_1_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_1_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_1_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_1_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_1_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_1_port, QN => n_1966);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_2_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_2_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_2_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_2_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_2_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_2_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_2_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_2_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_2_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_2_port, QN => n_1967);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_3_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_3_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_3_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_3_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_3_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_3_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_3_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_3_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_3_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_3_port, QN => n_1968);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_4_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_4_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_4_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_4_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_4_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_4_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_4_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_4_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_4_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_4_port, QN => n_1969);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_5_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_5_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_5_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_5_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_5_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_5_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_5_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_5_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_5_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_5_port, QN => n_1970);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_6_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_6_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_6_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_6_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_6_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_6_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_6_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_6_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_6_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_6_port, QN => n_1971);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_7_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_7_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_7_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_7_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_7_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_7_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_7_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_7_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_7_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_7_port, QN => n_1972);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_8_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_8_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_8_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_8_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_8_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_8_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_8_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_8_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_8_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_8_port, QN => n_1973);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_9_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_9_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_9_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_9_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_9_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_9_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_9_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_9_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_9_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_9_port, QN => n_1974);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_10_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_10_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_10_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_10_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_10_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_10_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_10_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_10_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n13, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_10_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_10_port, QN => n_1975);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_11_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_11_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_11_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_11_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_11_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n9, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_11_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_11_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_11_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_11_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_11_port, QN => n_1976);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_12_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_12_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_12_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_12_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_12_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_12_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_12_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_12_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_12_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_12_port, QN => n_1977);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_13_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_13_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_13_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_13_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_13_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_13_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_13_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_13_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_13_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_13_port, QN => n_1978);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_14_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_14_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_14_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_14_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_14_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_14_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_14_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_14_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_14_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_14_port, QN => n_1979);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_15_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_15_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_15_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_15_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_15_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_15_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_15_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_15_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_15_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_15_port, QN => n_1980);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_16_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_16_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_16_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_16_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_16_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_16_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_16_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_16_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_16_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_16_port, QN => n_1981);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_17_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_17_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_17_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_17_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_17_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_17_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_17_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_17_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_17_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_17_port, QN => n_1982);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_18_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_18_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_18_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_18_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_18_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_18_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_18_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_18_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_18_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_18_port, QN => n_1983);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_19_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_19_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_19_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_19_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_19_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_19_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_19_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_19_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_19_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_19_port, QN => n_1984);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_20_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_20_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_20_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_20_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_20_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_20_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_20_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_20_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_20_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_20_port, QN => n_1985);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_21_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_21_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_21_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_21_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_21_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_21_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_21_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_21_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n14, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_21_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_21_port, QN => n_1986);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_22_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_22_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_22_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_22_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_22_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_22_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_22_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_22_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_22_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_22_port, QN => n_1987);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_23_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_23_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_23_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_23_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_23_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n10, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_23_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_23_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_23_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_23_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_23_port, QN => n_1988);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_24_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_24_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_24_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_24_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_24_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_24_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_24_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_24_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_24_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_24_port, QN => n_1989);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_25_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_25_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_25_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_25_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_25_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_25_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_25_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_25_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_25_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_25_port, QN => n_1990);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_26_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_26_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_26_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_26_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_26_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_26_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_26_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_26_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_26_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_26_port, QN => n_1991);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_27_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_27_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_27_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_27_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_27_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_27_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_27_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_27_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_27_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_27_port, QN => n_1992);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_28_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_28_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_28_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_28_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_28_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_28_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_28_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_28_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_28_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_28_port, QN => n_1993);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_29_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_29_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_29_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_29_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_29_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_29_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_29_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_29_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_29_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_29_port, QN => n_1994);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_30_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_30_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_30_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_30_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_30_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_30_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_30_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_30_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_30_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_30_port, QN => n_1995);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_31_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_IR_OUT4s_31_port, B => 
                           DLX_INST_DATA_PATH_IR_OUT3s_31_port, S => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, Z => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_31_n1);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_31_U2 : NAND2_X1 port map( A1 => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n11, A2 => 
                           DLX_INST_DATA_PATH_MEMORY_Logic1_port, ZN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_31_n2);
   DLX_INST_DATA_PATH_MEMORY_IR4_FF_31_Q_reg : DFFR_X1 port map( D => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_31_n1, CK => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_n15, RN => 
                           DLX_INST_DATA_PATH_MEMORY_IR4_FF_31_n2, Q => 
                           DLX_INST_DATA_PATH_IR_OUT4s_31_port, QN => n_1996);
   DLX_INST_DATA_PATH_WB_MUXWB_U32 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_0_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_0_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_0_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U31 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_10_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_10_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_10_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U30 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_11_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_11_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_11_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U29 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_12_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_12_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_12_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U28 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_13_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_13_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_13_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U27 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_14_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_14_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_14_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U26 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_15_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_15_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_15_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U25 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_16_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_16_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_16_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U24 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_17_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_17_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_17_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U23 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_18_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_18_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_18_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U22 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_19_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_19_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_19_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U21 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_1_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_1_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_1_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U20 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_20_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_20_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_20_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U19 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_21_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_21_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_21_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U18 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_22_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_22_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_22_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U17 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_23_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_23_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_23_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U16 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_24_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_24_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_24_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U15 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_25_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_25_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_25_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U14 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_26_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_26_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_26_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U13 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_27_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_27_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_27_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U12 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_28_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_28_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_28_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U11 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_29_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_29_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_29_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U10 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_2_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_2_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_2_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U9 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_30_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_30_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_30_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U8 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_31_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_31_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_31_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U7 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_3_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_3_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_3_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U6 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_4_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_4_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_4_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U5 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_5_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_5_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_5_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U4 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_6_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_6_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_6_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U3 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_7_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_7_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_7_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U2 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_8_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_8_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_8_port);
   DLX_INST_DATA_PATH_WB_MUXWB_U1 : MUX2_X1 port map( A => 
                           DLX_INST_DATA_PATH_LMD_OUTs_9_port, B => 
                           DLX_INST_DATA_PATH_ALU_OUT2s_9_port, S => 
                           DLX_INST_WB_MUX_SEL_signal, Z => 
                           DLX_INST_DATA_PATH_DATAIN_RFs_9_port);

end SYN_STRUCTURAL;
