
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_dlx is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (LLS, LRS, ADDS, SUBS, ANDS, ORS, XORS, SNES, SLES, SGES, NOP);
attribute ENUM_ENCODING of aluOp : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";

end CONV_PACK_dlx;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_1;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_1;

architecture SYN_STRUCTURAL of RCA_NBITS4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_2;

architecture SYN_STRUCTURAL of RCA_NBITS4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_2;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_3;

architecture SYN_STRUCTURAL of RCA_NBITS4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_4;

architecture SYN_STRUCTURAL of RCA_NBITS4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_3;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_5;

architecture SYN_STRUCTURAL of RCA_NBITS4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_6;

architecture SYN_STRUCTURAL of RCA_NBITS4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_4;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_7;

architecture SYN_STRUCTURAL of RCA_NBITS4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_8;

architecture SYN_STRUCTURAL of RCA_NBITS4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_5;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_9;

architecture SYN_STRUCTURAL of RCA_NBITS4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_10;

architecture SYN_STRUCTURAL of RCA_NBITS4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_6;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_11;

architecture SYN_STRUCTURAL of RCA_NBITS4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_12;

architecture SYN_STRUCTURAL of RCA_NBITS4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_7;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_13;

architecture SYN_STRUCTURAL of RCA_NBITS4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_14;

architecture SYN_STRUCTURAL of RCA_NBITS4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_bits4_0;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits4_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_15;

architecture SYN_STRUCTURAL of RCA_NBITS4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBITS4_0;

architecture SYN_STRUCTURAL of RCA_NBITS4_0 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_1 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_1;

architecture SYN_BEHAVIORAL of G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_2 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_2;

architecture SYN_BEHAVIORAL of G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_3 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_3;

architecture SYN_BEHAVIORAL of G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_4 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_4;

architecture SYN_BEHAVIORAL of G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_1 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_1;

architecture SYN_BEHAVIORAL of PG_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_2 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_2;

architecture SYN_BEHAVIORAL of PG_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_5 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_5;

architecture SYN_BEHAVIORAL of G_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_6 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_6;

architecture SYN_BEHAVIORAL of G_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_3 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_3;

architecture SYN_BEHAVIORAL of PG_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_4 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_4;

architecture SYN_BEHAVIORAL of PG_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_5 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_5;

architecture SYN_BEHAVIORAL of PG_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_7 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_7;

architecture SYN_BEHAVIORAL of G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_6 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_6;

architecture SYN_BEHAVIORAL of PG_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_7 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_7;

architecture SYN_BEHAVIORAL of PG_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_8 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_8;

architecture SYN_BEHAVIORAL of PG_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_9 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_9;

architecture SYN_BEHAVIORAL of PG_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_10 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_10;

architecture SYN_BEHAVIORAL of PG_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_11 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_11;

architecture SYN_BEHAVIORAL of PG_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_12 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_12;

architecture SYN_BEHAVIORAL of PG_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_8 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_8;

architecture SYN_BEHAVIORAL of G_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_13 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_13;

architecture SYN_BEHAVIORAL of PG_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_14 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_14;

architecture SYN_BEHAVIORAL of PG_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_15 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_15;

architecture SYN_BEHAVIORAL of PG_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_16 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_16;

architecture SYN_BEHAVIORAL of PG_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_17 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_17;

architecture SYN_BEHAVIORAL of PG_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_18 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_18;

architecture SYN_BEHAVIORAL of PG_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_19 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_19;

architecture SYN_BEHAVIORAL of PG_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_20 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_20;

architecture SYN_BEHAVIORAL of PG_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_21 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_21;

architecture SYN_BEHAVIORAL of PG_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_22 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_22;

architecture SYN_BEHAVIORAL of PG_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_23 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_23;

architecture SYN_BEHAVIORAL of PG_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_24 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_24;

architecture SYN_BEHAVIORAL of PG_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_25 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_25;

architecture SYN_BEHAVIORAL of PG_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_26 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_26;

architecture SYN_BEHAVIORAL of PG_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_0 is

   port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out std_logic);

end PG_0;

architecture SYN_BEHAVIORAL of PG_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);
   U3 : AND2_X1 port map( A1 => p_k1j, A2 => p_ik, ZN => P_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_0 is

   port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);

end G_0;

architecture SYN_BEHAVIORAL of G_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => p_ik, B2 => g_k1j, A => g_ik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_1 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_1;

architecture SYN_BEHAVIORAL of pg_generator_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_2 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_2;

architecture SYN_BEHAVIORAL of pg_generator_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_3 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_3;

architecture SYN_BEHAVIORAL of pg_generator_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_4 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_4;

architecture SYN_BEHAVIORAL of pg_generator_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_5 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_5;

architecture SYN_BEHAVIORAL of pg_generator_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_6 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_6;

architecture SYN_BEHAVIORAL of pg_generator_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_7 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_7;

architecture SYN_BEHAVIORAL of pg_generator_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_8 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_8;

architecture SYN_BEHAVIORAL of pg_generator_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_9 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_9;

architecture SYN_BEHAVIORAL of pg_generator_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_10 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_10;

architecture SYN_BEHAVIORAL of pg_generator_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_11 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_11;

architecture SYN_BEHAVIORAL of pg_generator_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_12 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_12;

architecture SYN_BEHAVIORAL of pg_generator_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_13 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_13;

architecture SYN_BEHAVIORAL of pg_generator_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_14 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_14;

architecture SYN_BEHAVIORAL of pg_generator_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_15 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_15;

architecture SYN_BEHAVIORAL of pg_generator_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_16 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_16;

architecture SYN_BEHAVIORAL of pg_generator_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_17 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_17;

architecture SYN_BEHAVIORAL of pg_generator_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_18 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_18;

architecture SYN_BEHAVIORAL of pg_generator_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_19 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_19;

architecture SYN_BEHAVIORAL of pg_generator_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_20 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_20;

architecture SYN_BEHAVIORAL of pg_generator_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_21 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_21;

architecture SYN_BEHAVIORAL of pg_generator_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_22 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_22;

architecture SYN_BEHAVIORAL of pg_generator_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_23 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_23;

architecture SYN_BEHAVIORAL of pg_generator_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_24 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_24;

architecture SYN_BEHAVIORAL of pg_generator_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_25 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_25;

architecture SYN_BEHAVIORAL of pg_generator_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_26 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_26;

architecture SYN_BEHAVIORAL of pg_generator_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_27 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_27;

architecture SYN_BEHAVIORAL of pg_generator_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_28 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_28;

architecture SYN_BEHAVIORAL of pg_generator_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_29 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_29;

architecture SYN_BEHAVIORAL of pg_generator_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_30 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_30;

architecture SYN_BEHAVIORAL of pg_generator_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_31 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_31;

architecture SYN_BEHAVIORAL of pg_generator_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity pg_generator_0 is

   port( A, B : in std_logic;  P, G : out std_logic);

end pg_generator_0;

architecture SYN_BEHAVIORAL of pg_generator_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_1;

architecture SYN_STRUCTURAL of CarrySelect_1 is

   component MUX21_GENERIC_bits4_1
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1000, n_1001 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1000);
   RCA2 : RCA_NBITS4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1001);
   MUX21_GEN : MUX21_GENERIC_bits4_1 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_2;

architecture SYN_STRUCTURAL of CarrySelect_2 is

   component MUX21_GENERIC_bits4_2
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1002, n_1003 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1002);
   RCA2 : RCA_NBITS4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1003);
   MUX21_GEN : MUX21_GENERIC_bits4_2 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_3;

architecture SYN_STRUCTURAL of CarrySelect_3 is

   component MUX21_GENERIC_bits4_3
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1004, n_1005 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1004);
   RCA2 : RCA_NBITS4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1005);
   MUX21_GEN : MUX21_GENERIC_bits4_3 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_4;

architecture SYN_STRUCTURAL of CarrySelect_4 is

   component MUX21_GENERIC_bits4_4
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1006, n_1007 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1006);
   RCA2 : RCA_NBITS4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1007);
   MUX21_GEN : MUX21_GENERIC_bits4_4 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_5;

architecture SYN_STRUCTURAL of CarrySelect_5 is

   component MUX21_GENERIC_bits4_5
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1008, n_1009 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1008);
   RCA2 : RCA_NBITS4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1009);
   MUX21_GEN : MUX21_GENERIC_bits4_5 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_6;

architecture SYN_STRUCTURAL of CarrySelect_6 is

   component MUX21_GENERIC_bits4_6
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1010, n_1011 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1010);
   RCA2 : RCA_NBITS4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1011);
   MUX21_GEN : MUX21_GENERIC_bits4_6 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_7;

architecture SYN_STRUCTURAL of CarrySelect_7 is

   component MUX21_GENERIC_bits4_7
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1012, n_1013 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1012);
   RCA2 : RCA_NBITS4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1013);
   MUX21_GEN : MUX21_GENERIC_bits4_7 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CarrySelect_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end CarrySelect_0;

architecture SYN_STRUCTURAL of CarrySelect_0 is

   component MUX21_GENERIC_bits4_0
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBITS4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBITS4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, 
      sum2_3_port, sum2_2_port, sum2_1_port, sum2_0_port, n_1014, n_1015 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RCA1 : RCA_NBITS4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1014);
   RCA2 : RCA_NBITS4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum2_3_port, S(2) => sum2_2_port, S(1) => 
                           sum2_1_port, S(0) => sum2_0_port, Co => n_1015);
   MUX21_GEN : MUX21_GENERIC_bits4_0 port map( A(3) => sum2_3_port, A(2) => 
                           sum2_2_port, A(1) => sum2_1_port, A(0) => 
                           sum2_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity logic_and_shift_N32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end logic_and_shift_N32_DW01_ash_0;

architecture SYN_mx2 of logic_and_shift_N32_DW01_ash_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal temp_int_SH_4_port, temp_int_SH_3_port, temp_int_SH_2_port, 
      temp_int_SH_1_port, temp_int_SH_0_port, SHMAG_5_port, ML_int_1_31_port, 
      ML_int_1_30_port, ML_int_1_29_port, ML_int_1_28_port, ML_int_1_27_port, 
      ML_int_1_26_port, ML_int_1_25_port, ML_int_1_24_port, ML_int_1_23_port, 
      ML_int_1_22_port, ML_int_1_21_port, ML_int_1_20_port, ML_int_1_19_port, 
      ML_int_1_18_port, ML_int_1_17_port, ML_int_1_16_port, ML_int_1_15_port, 
      ML_int_1_14_port, ML_int_1_13_port, ML_int_1_12_port, ML_int_1_11_port, 
      ML_int_1_10_port, ML_int_1_9_port, ML_int_1_8_port, ML_int_1_7_port, 
      ML_int_1_6_port, ML_int_1_5_port, ML_int_1_4_port, ML_int_1_3_port, 
      ML_int_1_2_port, ML_int_1_1_port, ML_int_1_0_port, ML_int_2_31_port, 
      ML_int_2_30_port, ML_int_2_29_port, ML_int_2_28_port, ML_int_2_27_port, 
      ML_int_2_26_port, ML_int_2_25_port, ML_int_2_24_port, ML_int_2_23_port, 
      ML_int_2_22_port, ML_int_2_21_port, ML_int_2_20_port, ML_int_2_19_port, 
      ML_int_2_18_port, ML_int_2_17_port, ML_int_2_16_port, ML_int_2_15_port, 
      ML_int_2_14_port, ML_int_2_13_port, ML_int_2_12_port, ML_int_2_11_port, 
      ML_int_2_10_port, ML_int_2_9_port, ML_int_2_8_port, ML_int_2_7_port, 
      ML_int_2_6_port, ML_int_2_5_port, ML_int_2_4_port, ML_int_2_3_port, 
      ML_int_2_2_port, ML_int_2_1_port, ML_int_2_0_port, ML_int_3_31_port, 
      ML_int_3_30_port, ML_int_3_29_port, ML_int_3_28_port, ML_int_3_27_port, 
      ML_int_3_26_port, ML_int_3_25_port, ML_int_3_24_port, ML_int_3_23_port, 
      ML_int_3_22_port, ML_int_3_21_port, ML_int_3_20_port, ML_int_3_19_port, 
      ML_int_3_18_port, ML_int_3_17_port, ML_int_3_16_port, ML_int_3_15_port, 
      ML_int_3_14_port, ML_int_3_13_port, ML_int_3_12_port, ML_int_3_11_port, 
      ML_int_3_10_port, ML_int_3_9_port, ML_int_3_8_port, ML_int_3_7_port, 
      ML_int_3_6_port, ML_int_3_5_port, ML_int_3_4_port, ML_int_3_3_port, 
      ML_int_3_2_port, ML_int_3_1_port, ML_int_3_0_port, ML_int_4_31_port, 
      ML_int_4_30_port, ML_int_4_29_port, ML_int_4_28_port, ML_int_4_27_port, 
      ML_int_4_26_port, ML_int_4_25_port, ML_int_4_24_port, ML_int_4_23_port, 
      ML_int_4_22_port, ML_int_4_21_port, ML_int_4_20_port, ML_int_4_19_port, 
      ML_int_4_18_port, ML_int_4_17_port, ML_int_4_16_port, ML_int_4_15_port, 
      ML_int_4_14_port, ML_int_4_13_port, ML_int_4_12_port, ML_int_4_11_port, 
      ML_int_4_10_port, ML_int_4_9_port, ML_int_4_8_port, ML_int_5_31_port, 
      ML_int_5_30_port, ML_int_5_29_port, ML_int_5_28_port, ML_int_5_27_port, 
      ML_int_5_26_port, ML_int_5_25_port, ML_int_5_24_port, ML_int_5_23_port, 
      ML_int_5_22_port, ML_int_5_21_port, ML_int_5_20_port, ML_int_5_19_port, 
      ML_int_5_18_port, ML_int_5_17_port, ML_int_5_16_port, n28, n29, n30, n31,
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_31_port);
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_30_port);
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_29_port);
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_28_port);
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_27_port);
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_26_port);
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_25_port);
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => temp_int_SH_4_port, Z => ML_int_5_24_port);
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => n71, S => 
                           temp_int_SH_4_port, Z => ML_int_5_23_port);
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => n67, S => 
                           temp_int_SH_4_port, Z => ML_int_5_22_port);
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => n69, S => 
                           temp_int_SH_4_port, Z => ML_int_5_21_port);
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => n65, S => 
                           temp_int_SH_4_port, Z => ML_int_5_20_port);
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => n70, S => 
                           temp_int_SH_4_port, Z => ML_int_5_19_port);
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => n66, S => 
                           temp_int_SH_4_port, Z => ML_int_5_18_port);
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => n68, S => 
                           temp_int_SH_4_port, Z => ML_int_5_17_port);
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => n64, S => 
                           temp_int_SH_4_port, Z => ML_int_5_16_port);
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => temp_int_SH_3_port, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           temp_int_SH_3_port, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           temp_int_SH_3_port, Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => temp_int_SH_2_port, Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => temp_int_SH_1_port, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           temp_int_SH_1_port, Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => temp_int_SH_0_port,
                           Z => ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => temp_int_SH_0_port,
                           Z => ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => temp_int_SH_0_port,
                           Z => ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => temp_int_SH_0_port,
                           Z => ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => temp_int_SH_0_port,
                           Z => ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => temp_int_SH_0_port,
                           Z => ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => temp_int_SH_0_port,
                           Z => ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => temp_int_SH_0_port,
                           Z => ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => temp_int_SH_0_port,
                           Z => ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => temp_int_SH_0_port,
                           Z => ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => temp_int_SH_0_port,
                           Z => ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => temp_int_SH_0_port,
                           Z => ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => temp_int_SH_0_port,
                           Z => ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => temp_int_SH_0_port,
                           Z => ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => temp_int_SH_0_port,
                           Z => ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => temp_int_SH_0_port,
                           Z => ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => temp_int_SH_0_port,
                           Z => ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => temp_int_SH_0_port,
                           Z => ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => temp_int_SH_0_port,
                           Z => ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => temp_int_SH_0_port,
                           Z => ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => temp_int_SH_0_port,
                           Z => ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => temp_int_SH_0_port, 
                           Z => ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => temp_int_SH_0_port, Z 
                           => ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => temp_int_SH_0_port, Z 
                           => ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => temp_int_SH_0_port, Z 
                           => ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => temp_int_SH_0_port, Z 
                           => ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => temp_int_SH_0_port, Z 
                           => ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => temp_int_SH_0_port, Z 
                           => ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => temp_int_SH_0_port, Z 
                           => ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => temp_int_SH_0_port, Z 
                           => ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => temp_int_SH_0_port, Z 
                           => ML_int_1_1_port);
   U3 : NAND2_X2 port map( A1 => n38, A2 => n44, ZN => temp_int_SH_1_port);
   U4 : NAND2_X2 port map( A1 => n38, A2 => n45, ZN => temp_int_SH_0_port);
   U5 : NAND2_X2 port map( A1 => n38, A2 => n42, ZN => temp_int_SH_3_port);
   U6 : NAND2_X2 port map( A1 => n38, A2 => n43, ZN => temp_int_SH_2_port);
   U94 : NAND3_X1 port map( A1 => SH(11), A2 => SH(10), A3 => SH(12), ZN => n51
                           );
   U96 : NAND3_X1 port map( A1 => SH(17), A2 => SH(16), A3 => SH(18), ZN => n52
                           );
   U98 : NAND3_X1 port map( A1 => SH(23), A2 => SH(22), A3 => SH(24), ZN => n53
                           );
   U100 : NAND3_X1 port map( A1 => SH(29), A2 => SH(28), A3 => SH(6), ZN => n54
                           );
   U104 : NAND3_X1 port map( A1 => n79, A2 => n80, A3 => n78, ZN => n60);
   U106 : NAND3_X1 port map( A1 => n88, A2 => n89, A3 => n87, ZN => n61);
   U108 : NAND3_X1 port map( A1 => n85, A2 => n86, A3 => n84, ZN => n62);
   U110 : NAND3_X1 port map( A1 => n82, A2 => n83, A3 => n81, ZN => n63);
   U7 : INV_X1 port map( A => n37, ZN => n64);
   U8 : INV_X1 port map( A => n36, ZN => n68);
   U9 : INV_X1 port map( A => n35, ZN => n66);
   U10 : INV_X1 port map( A => n33, ZN => n70);
   U11 : INV_X1 port map( A => n32, ZN => n65);
   U12 : INV_X1 port map( A => n31, ZN => n69);
   U13 : INV_X1 port map( A => n30, ZN => n67);
   U14 : INV_X1 port map( A => n29, ZN => n71);
   U15 : INV_X1 port map( A => n28, ZN => n76);
   U16 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => n75, ZN => n33);
   U17 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => n75, ZN => n32);
   U18 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => n75, ZN => n31);
   U19 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => n75, ZN => n30);
   U20 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => n75, ZN => n29);
   U21 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => n75, ZN => n37);
   U22 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => n75, ZN => n36);
   U23 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => n75, ZN => n35);
   U24 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => n74, ZN => 
                           ML_int_3_3_port);
   U25 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => n74, ZN => 
                           ML_int_3_0_port);
   U26 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => n74, ZN => 
                           ML_int_3_1_port);
   U27 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => n74, ZN => 
                           ML_int_3_2_port);
   U28 : NAND2_X1 port map( A1 => n34, A2 => n77, ZN => n28);
   U29 : INV_X1 port map( A => temp_int_SH_4_port, ZN => n77);
   U30 : INV_X1 port map( A => temp_int_SH_3_port, ZN => n75);
   U31 : INV_X1 port map( A => temp_int_SH_2_port, ZN => n74);
   U32 : INV_X1 port map( A => temp_int_SH_1_port, ZN => n73);
   U33 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => n73, ZN => 
                           ML_int_2_0_port);
   U34 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => n73, ZN => 
                           ML_int_2_1_port);
   U35 : NAND2_X1 port map( A1 => SH(0), A2 => n40, ZN => n45);
   U36 : NAND2_X1 port map( A1 => SH(1), A2 => n40, ZN => n44);
   U37 : NAND2_X1 port map( A1 => SH(2), A2 => n40, ZN => n43);
   U38 : NAND2_X1 port map( A1 => SH(3), A2 => n40, ZN => n42);
   U39 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => temp_int_SH_4_port);
   U40 : NAND2_X1 port map( A1 => SH(4), A2 => n40, ZN => n39);
   U41 : NOR4_X1 port map( A1 => n60, A2 => SH(28), A3 => SH(6), A4 => SH(29), 
                           ZN => n59);
   U42 : AND2_X1 port map( A1 => SHMAG_5_port, A2 => n90, ZN => n34);
   U43 : AND2_X1 port map( A1 => n38, A2 => n41, ZN => SHMAG_5_port);
   U44 : NAND2_X1 port map( A1 => SH(5), A2 => n40, ZN => n41);
   U45 : NOR4_X1 port map( A1 => n61, A2 => SH(22), A3 => SH(24), A4 => SH(23),
                           ZN => n58);
   U46 : NOR4_X1 port map( A1 => n51, A2 => n83, A3 => n81, A4 => n82, ZN => 
                           n50);
   U47 : NOR4_X1 port map( A1 => n52, A2 => n86, A3 => n84, A4 => n85, ZN => 
                           n49);
   U48 : NAND2_X1 port map( A1 => SH(30), A2 => n46, ZN => n40);
   U49 : NAND4_X1 port map( A1 => n47, A2 => n48, A3 => n49, A4 => n50, ZN => 
                           n46);
   U50 : NOR4_X1 port map( A1 => n54, A2 => n80, A3 => n78, A4 => n79, ZN => 
                           n47);
   U51 : NOR4_X1 port map( A1 => n53, A2 => n89, A3 => n87, A4 => n88, ZN => 
                           n48);
   U52 : NAND2_X1 port map( A1 => n55, A2 => n90, ZN => n38);
   U53 : NAND4_X1 port map( A1 => n56, A2 => n57, A3 => n58, A4 => n59, ZN => 
                           n55);
   U54 : NOR4_X1 port map( A1 => n63, A2 => SH(10), A3 => SH(12), A4 => SH(11),
                           ZN => n56);
   U55 : NOR4_X1 port map( A1 => n62, A2 => SH(16), A3 => SH(18), A4 => SH(17),
                           ZN => n57);
   U56 : INV_X1 port map( A => SH(30), ZN => n90);
   U57 : INV_X1 port map( A => SH(26), ZN => n88);
   U58 : INV_X1 port map( A => SH(13), ZN => n81);
   U59 : INV_X1 port map( A => SH(25), ZN => n87);
   U60 : INV_X1 port map( A => SH(14), ZN => n82);
   U61 : INV_X1 port map( A => SH(27), ZN => n89);
   U62 : INV_X1 port map( A => SH(15), ZN => n83);
   U63 : INV_X1 port map( A => SH(8), ZN => n79);
   U64 : INV_X1 port map( A => SH(20), ZN => n85);
   U65 : INV_X1 port map( A => SH(19), ZN => n84);
   U66 : INV_X1 port map( A => SH(7), ZN => n78);
   U67 : INV_X1 port map( A => SH(21), ZN => n86);
   U68 : INV_X1 port map( A => SH(9), ZN => n80);
   U69 : AND2_X1 port map( A1 => A(0), A2 => n72, ZN => ML_int_1_0_port);
   U70 : INV_X1 port map( A => temp_int_SH_0_port, ZN => n72);
   U71 : NOR2_X1 port map( A1 => n28, A2 => n37, ZN => B(0));
   U72 : NOR2_X1 port map( A1 => n28, A2 => n36, ZN => B(1));
   U73 : NOR2_X1 port map( A1 => n28, A2 => n35, ZN => B(2));
   U74 : NOR2_X1 port map( A1 => n28, A2 => n33, ZN => B(3));
   U75 : NOR2_X1 port map( A1 => n28, A2 => n32, ZN => B(4));
   U76 : NOR2_X1 port map( A1 => n28, A2 => n31, ZN => B(5));
   U77 : NOR2_X1 port map( A1 => n28, A2 => n30, ZN => B(6));
   U78 : NOR2_X1 port map( A1 => n28, A2 => n29, ZN => B(7));
   U79 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n76, ZN => B(8));
   U80 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n76, ZN => B(9));
   U81 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n76, ZN => B(10));
   U82 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n76, ZN => B(11));
   U83 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n76, ZN => B(12));
   U84 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n76, ZN => B(13));
   U85 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n76, ZN => B(14));
   U86 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n76, ZN => B(15));
   U87 : AND2_X1 port map( A1 => ML_int_5_16_port, A2 => n34, ZN => B(16));
   U88 : AND2_X1 port map( A1 => ML_int_5_17_port, A2 => n34, ZN => B(17));
   U89 : AND2_X1 port map( A1 => ML_int_5_18_port, A2 => n34, ZN => B(18));
   U90 : AND2_X1 port map( A1 => ML_int_5_19_port, A2 => n34, ZN => B(19));
   U91 : AND2_X1 port map( A1 => ML_int_5_20_port, A2 => n34, ZN => B(20));
   U92 : AND2_X1 port map( A1 => ML_int_5_21_port, A2 => n34, ZN => B(21));
   U93 : AND2_X1 port map( A1 => ML_int_5_22_port, A2 => n34, ZN => B(22));
   U95 : AND2_X1 port map( A1 => ML_int_5_23_port, A2 => n34, ZN => B(23));
   U97 : AND2_X1 port map( A1 => ML_int_5_24_port, A2 => n34, ZN => B(24));
   U99 : AND2_X1 port map( A1 => ML_int_5_25_port, A2 => n34, ZN => B(25));
   U101 : AND2_X1 port map( A1 => ML_int_5_26_port, A2 => n34, ZN => B(26));
   U102 : AND2_X1 port map( A1 => ML_int_5_27_port, A2 => n34, ZN => B(27));
   U103 : AND2_X1 port map( A1 => ML_int_5_28_port, A2 => n34, ZN => B(28));
   U105 : AND2_X1 port map( A1 => ML_int_5_29_port, A2 => n34, ZN => B(29));
   U107 : AND2_X1 port map( A1 => ML_int_5_30_port, A2 => n34, ZN => B(30));
   U109 : AND2_X1 port map( A1 => ML_int_5_31_port, A2 => n34, ZN => B(31));

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity logic_and_shift_N32_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end logic_and_shift_N32_DW_rash_0;

architecture SYN_mx2 of logic_and_shift_N32_DW_rash_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247 : std_logic;

begin
   
   U3 : NOR2_X2 port map( A1 => n238, A2 => SH(1), ZN => n116);
   U4 : NOR2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n117);
   U81 : MUX2_X1 port map( A => n193, B => n102, S => SH(4), Z => n94);
   U89 : MUX2_X1 port map( A => n112, B => n214, S => SH(4), Z => n111);
   U113 : MUX2_X1 port map( A => n133, B => n213, S => SH(4), Z => n132);
   U151 : MUX2_X1 port map( A => n125, B => n107, S => SH(2), Z => n120);
   U195 : MUX2_X1 port map( A => n178, B => n210, S => SH(4), Z => n177);
   U5 : NOR2_X1 port map( A1 => n243, A2 => SH(3), ZN => n123);
   U6 : NOR2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n122);
   U7 : NOR2_X1 port map( A1 => n246, A2 => n242, ZN => n67);
   U8 : INV_X1 port map( A => n100, ZN => n237);
   U9 : INV_X1 port map( A => n101, ZN => n239);
   U10 : NAND2_X1 port map( A1 => n122, A2 => n163, ZN => n62);
   U11 : INV_X1 port map( A => n117, ZN => n240);
   U12 : INV_X1 port map( A => n116, ZN => n236);
   U13 : AOI222_X1 port map( A1 => n222, A2 => n123, B1 => n231, B2 => n241, C1
                           => n74, C2 => n122, ZN => n91);
   U14 : AOI222_X1 port map( A1 => n224, A2 => n123, B1 => n233, B2 => n241, C1
                           => n66, C2 => n122, ZN => n88);
   U15 : AOI222_X1 port map( A1 => n227, A2 => n123, B1 => n234, B2 => n241, C1
                           => n127, C2 => n122, ZN => n82);
   U16 : INV_X1 port map( A => n163, ZN => n246);
   U17 : AOI221_X1 port map( B1 => n74, B2 => n123, C1 => n75, C2 => n122, A =>
                           n179, ZN => n141);
   U18 : OAI22_X1 port map( A1 => n104, A2 => n119, B1 => n105, B2 => n129, ZN 
                           => n179);
   U19 : AOI221_X1 port map( B1 => n66, B2 => n123, C1 => n70, C2 => n122, A =>
                           n140, ZN => n134);
   U20 : OAI22_X1 port map( A1 => n104, A2 => n118, B1 => n105, B2 => n128, ZN 
                           => n140);
   U21 : AOI221_X1 port map( B1 => n127, B2 => n123, C1 => n84, C2 => n122, A 
                           => n138, ZN => n113);
   U22 : OAI22_X1 port map( A1 => n104, A2 => n108, B1 => n105, B2 => n139, ZN 
                           => n138);
   U23 : AND2_X1 port map( A1 => n161, A2 => n243, ZN => n69);
   U24 : NOR2_X1 port map( A1 => n64, A2 => n245, ZN => n144);
   U25 : AOI22_X1 port map( A1 => n222, A2 => n122, B1 => n231, B2 => n123, ZN 
                           => n72);
   U26 : AOI22_X1 port map( A1 => n224, A2 => n122, B1 => n233, B2 => n123, ZN 
                           => n63);
   U27 : AOI22_X1 port map( A1 => n227, A2 => n122, B1 => n234, B2 => n123, ZN 
                           => n121);
   U28 : INV_X1 port map( A => n142, ZN => n244);
   U29 : INV_X1 port map( A => n123, ZN => n242);
   U30 : INV_X1 port map( A => n122, ZN => n245);
   U31 : INV_X1 port map( A => n105, ZN => n241);
   U32 : INV_X1 port map( A => n118, ZN => n233);
   U33 : INV_X1 port map( A => n108, ZN => n234);
   U34 : INV_X1 port map( A => n119, ZN => n231);
   U35 : OAI21_X1 port map( B1 => n97, B2 => n98, A => n99, ZN => n95);
   U36 : OAI22_X1 port map( A1 => n100, A2 => n191, B1 => n101, B2 => n192, ZN 
                           => n97);
   U37 : OAI22_X1 port map( A1 => n240, A2 => n189, B1 => n236, B2 => n190, ZN 
                           => n98);
   U38 : INV_X1 port map( A => n93, ZN => n204);
   U39 : INV_X1 port map( A => n129, ZN => n222);
   U40 : INV_X1 port map( A => n128, ZN => n224);
   U41 : INV_X1 port map( A => n139, ZN => n227);
   U42 : INV_X1 port map( A => n126, ZN => n219);
   U43 : INV_X1 port map( A => n85, ZN => n207);
   U44 : INV_X1 port map( A => n61, ZN => n197);
   U45 : INV_X1 port map( A => n86, ZN => n199);
   U46 : INV_X1 port map( A => n71, ZN => n195);
   U47 : INV_X1 port map( A => n68, ZN => n206);
   U48 : INV_X1 port map( A => n79, ZN => n208);
   U49 : INV_X1 port map( A => n80, ZN => n202);
   U50 : INV_X1 port map( A => n124, ZN => n220);
   U51 : OAI222_X1 port map( A1 => n125, A2 => n242, B1 => n107, B2 => n105, C1
                           => n126, C2 => n245, ZN => n124);
   U52 : INV_X1 port map( A => n107, ZN => n235);
   U53 : INV_X1 port map( A => n103, ZN => n193);
   U54 : OAI222_X1 port map( A1 => n242, A2 => n76, B1 => n104, B2 => n208, C1 
                           => n105, C2 => n80, ZN => n103);
   U55 : AOI222_X1 port map( A1 => n116, A2 => A(30), B1 => n237, B2 => A(31), 
                           C1 => n117, C2 => A(29), ZN => n118);
   U56 : AOI221_X1 port map( B1 => n239, B2 => A(27), C1 => n237, C2 => A(26), 
                           A => n180, ZN => n129);
   U57 : OAI22_X1 port map( A1 => n225, A2 => n236, B1 => n223, B2 => n240, ZN 
                           => n180);
   U58 : AOI221_X1 port map( B1 => n239, B2 => A(28), C1 => n237, C2 => A(27), 
                           A => n150, ZN => n128);
   U59 : OAI22_X1 port map( A1 => n226, A2 => n236, B1 => n225, B2 => n240, ZN 
                           => n150);
   U60 : INV_X1 port map( A => A(26), ZN => n226);
   U61 : AOI221_X1 port map( B1 => n239, B2 => A(29), C1 => n237, C2 => A(28), 
                           A => n228, ZN => n139);
   U62 : INV_X1 port map( A => n165, ZN => n228);
   U63 : AOI22_X1 port map( A1 => A(27), A2 => n116, B1 => A(26), B2 => n117, 
                           ZN => n165);
   U64 : AOI221_X1 port map( B1 => n239, B2 => A(12), C1 => n237, C2 => A(11), 
                           A => n136, ZN => n61);
   U65 : OAI22_X1 port map( A1 => n200, A2 => n236, B1 => n198, B2 => n240, ZN 
                           => n136);
   U66 : AOI221_X1 port map( B1 => n239, B2 => A(13), C1 => n237, C2 => A(12), 
                           A => n166, ZN => n86);
   U67 : OAI22_X1 port map( A1 => n201, A2 => n236, B1 => n200, B2 => n240, ZN 
                           => n166);
   U68 : INV_X1 port map( A => A(11), ZN => n201);
   U69 : AOI221_X1 port map( B1 => n239, B2 => A(31), C1 => n237, C2 => A(30), 
                           A => n232, ZN => n119);
   U70 : INV_X1 port map( A => n181, ZN => n232);
   U71 : AOI22_X1 port map( A1 => A(29), A2 => n116, B1 => A(28), B2 => n117, 
                           ZN => n181);
   U72 : AOI221_X1 port map( B1 => n239, B2 => A(26), C1 => n237, C2 => A(25), 
                           A => n158, ZN => n126);
   U73 : OAI22_X1 port map( A1 => n223, A2 => n236, B1 => n221, B2 => n240, ZN 
                           => n158);
   U74 : AOI221_X1 port map( B1 => n239, B2 => A(11), C1 => n237, C2 => A(10), 
                           A => n186, ZN => n71);
   U75 : OAI22_X1 port map( A1 => n198, A2 => n236, B1 => n196, B2 => n240, ZN 
                           => n186);
   U76 : AOI221_X1 port map( B1 => n239, B2 => A(15), C1 => n237, C2 => A(14), 
                           A => n205, ZN => n93);
   U77 : INV_X1 port map( A => n185, ZN => n205);
   U78 : AOI22_X1 port map( A1 => A(13), A2 => n116, B1 => A(12), B2 => n117, 
                           ZN => n185);
   U79 : AOI221_X1 port map( B1 => n239, B2 => A(14), C1 => n237, C2 => A(13), 
                           A => n203, ZN => n80);
   U80 : INV_X1 port map( A => n157, ZN => n203);
   U82 : AOI22_X1 port map( A1 => A(12), A2 => n116, B1 => A(11), B2 => n117, 
                           ZN => n157);
   U83 : NAND2_X1 port map( A1 => SH(1), A2 => SH(0), ZN => n101);
   U84 : NAND2_X1 port map( A1 => SH(1), A2 => n238, ZN => n100);
   U85 : AOI221_X1 port map( B1 => n239, B2 => A(30), C1 => n237, C2 => A(29), 
                           A => n230, ZN => n125);
   U86 : INV_X1 port map( A => n154, ZN => n230);
   U87 : AOI22_X1 port map( A1 => A(28), A2 => n116, B1 => A(27), B2 => n117, 
                           ZN => n154);
   U88 : OAI221_X1 port map( B1 => n101, B2 => n216, C1 => n100, C2 => n215, A 
                           => n147, ZN => n70);
   U90 : INV_X1 port map( A => A(19), ZN => n215);
   U91 : AOI22_X1 port map( A1 => A(18), A2 => n116, B1 => A(17), B2 => n117, 
                           ZN => n147);
   U92 : OAI221_X1 port map( B1 => n101, B2 => n217, C1 => n100, C2 => n216, A 
                           => n160, ZN => n84);
   U93 : AOI22_X1 port map( A1 => A(19), A2 => n116, B1 => A(18), B2 => n117, 
                           ZN => n160);
   U94 : OAI221_X1 port map( B1 => n236, B2 => n212, C1 => n211, C2 => n240, A 
                           => n182, ZN => n75);
   U95 : AOI22_X1 port map( A1 => A(19), A2 => n239, B1 => A(18), B2 => n237, 
                           ZN => n182);
   U96 : OAI221_X1 port map( B1 => n101, B2 => n218, C1 => n100, C2 => n217, A 
                           => n156, ZN => n78);
   U97 : AOI22_X1 port map( A1 => A(20), A2 => n116, B1 => A(19), B2 => n117, 
                           ZN => n156);
   U98 : OAI221_X1 port map( B1 => n101, B2 => n221, C1 => n100, C2 => n218, A 
                           => n183, ZN => n74);
   U99 : AOI22_X1 port map( A1 => A(21), A2 => n116, B1 => A(20), B2 => n117, 
                           ZN => n183);
   U100 : OAI221_X1 port map( B1 => n101, B2 => n223, C1 => n100, C2 => n221, A
                           => n148, ZN => n66);
   U101 : AOI22_X1 port map( A1 => A(22), A2 => n116, B1 => A(21), B2 => n117, 
                           ZN => n148);
   U102 : OAI221_X1 port map( B1 => n101, B2 => n225, C1 => n100, C2 => n223, A
                           => n164, ZN => n127);
   U103 : AOI22_X1 port map( A1 => A(23), A2 => n116, B1 => A(22), B2 => n117, 
                           ZN => n164);
   U104 : NAND2_X1 port map( A1 => SH(3), A2 => n243, ZN => n105);
   U105 : AOI221_X1 port map( B1 => n239, B2 => A(8), C1 => n237, C2 => A(7), A
                           => n135, ZN => n87);
   U106 : OAI22_X1 port map( A1 => n192, A2 => n236, B1 => n191, B2 => n240, ZN
                           => n135);
   U107 : AOI221_X1 port map( B1 => n239, B2 => A(9), C1 => n237, C2 => A(8), A
                           => n114, ZN => n81);
   U108 : OAI22_X1 port map( A1 => n194, A2 => n236, B1 => n192, B2 => n240, ZN
                           => n114);
   U109 : AOI221_X1 port map( B1 => n239, B2 => A(7), C1 => n237, C2 => A(6), A
                           => n184, ZN => n90);
   U110 : OAI22_X1 port map( A1 => n191, A2 => n236, B1 => n190, B2 => n240, ZN
                           => n184);
   U111 : NAND2_X1 port map( A1 => SH(4), A2 => n247, ZN => n64);
   U112 : INV_X1 port map( A => n96, ZN => n247);
   U114 : AOI221_X1 port map( B1 => n239, B2 => A(10), C1 => n237, C2 => A(9), 
                           A => n106, ZN => n76);
   U115 : OAI22_X1 port map( A1 => n196, A2 => n236, B1 => n194, B2 => n240, ZN
                           => n106);
   U116 : AOI222_X1 port map( A1 => n78, A2 => n122, B1 => n219, B2 => n123, C1
                           => n229, C2 => SH(3), ZN => n102);
   U117 : INV_X1 port map( A => n120, ZN => n229);
   U118 : OAI221_X1 port map( B1 => n101, B2 => n211, C1 => n100, C2 => n209, A
                           => n149, ZN => n68);
   U119 : AOI22_X1 port map( A1 => A(14), A2 => n116, B1 => A(13), B2 => n117, 
                           ZN => n149);
   U120 : OAI221_X1 port map( B1 => n101, B2 => n212, C1 => n211, C2 => n100, A
                           => n162, ZN => n85);
   U121 : AOI22_X1 port map( A1 => n116, A2 => A(15), B1 => n117, B2 => A(14), 
                           ZN => n162);
   U122 : OAI221_X1 port map( B1 => n211, B2 => n236, C1 => n209, C2 => n240, A
                           => n155, ZN => n79);
   U123 : AOI22_X1 port map( A1 => A(18), A2 => n239, B1 => A(17), B2 => n237, 
                           ZN => n155);
   U124 : NAND2_X1 port map( A1 => SH(3), A2 => SH(2), ZN => n104);
   U125 : AOI22_X1 port map( A1 => n117, A2 => A(30), B1 => n116, B2 => A(31), 
                           ZN => n108);
   U126 : NOR4_X1 port map( A1 => n172, A2 => SH(29), A3 => SH(5), A4 => SH(30)
                           , ZN => n171);
   U127 : OR4_X1 port map( A1 => SH(7), A2 => SH(6), A3 => SH(9), A4 => SH(8), 
                           ZN => n172);
   U128 : NOR2_X1 port map( A1 => n245, A2 => SH(4), ZN => n99);
   U129 : NAND4_X1 port map( A1 => n168, A2 => n169, A3 => n170, A4 => n171, ZN
                           => n96);
   U130 : NOR4_X1 port map( A1 => n175, A2 => SH(10), A3 => SH(12), A4 => 
                           SH(11), ZN => n168);
   U131 : NOR4_X1 port map( A1 => n174, A2 => SH(16), A3 => SH(18), A4 => 
                           SH(17), ZN => n169);
   U132 : NOR4_X1 port map( A1 => n173, A2 => SH(23), A3 => SH(25), A4 => 
                           SH(24), ZN => n170);
   U133 : NAND2_X1 port map( A1 => n161, A2 => SH(2), ZN => n142);
   U134 : OAI221_X1 port map( B1 => n101, B2 => n189, C1 => n100, C2 => n188, A
                           => n187, ZN => n176);
   U135 : INV_X1 port map( A => A(2), ZN => n188);
   U136 : AOI22_X1 port map( A1 => A(1), A2 => n116, B1 => A(0), B2 => n117, ZN
                           => n187);
   U137 : OAI221_X1 port map( B1 => n101, B2 => n190, C1 => n100, C2 => n189, A
                           => n137, ZN => n131);
   U138 : AOI22_X1 port map( A1 => A(2), A2 => n116, B1 => A(1), B2 => n117, ZN
                           => n137);
   U139 : OAI221_X1 port map( B1 => n101, B2 => n191, C1 => n100, C2 => n190, A
                           => n115, ZN => n110);
   U140 : AOI22_X1 port map( A1 => A(3), A2 => n116, B1 => A(2), B2 => n117, ZN
                           => n115);
   U141 : NOR3_X1 port map( A1 => n64, A2 => SH(3), A3 => n120, ZN => n153);
   U142 : NOR2_X1 port map( A1 => n96, A2 => SH(4), ZN => n163);
   U143 : NAND2_X1 port map( A1 => A(31), A2 => n117, ZN => n107);
   U144 : INV_X1 port map( A => A(4), ZN => n190);
   U145 : INV_X1 port map( A => A(5), ZN => n191);
   U146 : INV_X1 port map( A => A(24), ZN => n223);
   U147 : INV_X1 port map( A => A(16), ZN => n211);
   U148 : INV_X1 port map( A => SH(2), ZN => n243);
   U149 : INV_X1 port map( A => A(3), ZN => n189);
   U150 : INV_X1 port map( A => A(6), ZN => n192);
   U152 : INV_X1 port map( A => A(23), ZN => n221);
   U153 : INV_X1 port map( A => A(25), ZN => n225);
   U154 : INV_X1 port map( A => SH(0), ZN => n238);
   U155 : INV_X1 port map( A => A(20), ZN => n216);
   U156 : INV_X1 port map( A => A(21), ZN => n217);
   U157 : INV_X1 port map( A => A(22), ZN => n218);
   U158 : INV_X1 port map( A => A(7), ZN => n194);
   U159 : INV_X1 port map( A => A(8), ZN => n196);
   U160 : INV_X1 port map( A => A(9), ZN => n198);
   U161 : INV_X1 port map( A => A(10), ZN => n200);
   U162 : INV_X1 port map( A => A(17), ZN => n212);
   U163 : INV_X1 port map( A => A(15), ZN => n209);
   U164 : INV_X1 port map( A => n141, ZN => n210);
   U165 : OAI222_X1 port map( A1 => n71, A2 => n105, B1 => n93, B2 => n104, C1 
                           => n90, C2 => n242, ZN => n178);
   U166 : INV_X1 port map( A => n134, ZN => n213);
   U167 : OAI222_X1 port map( A1 => n61, A2 => n105, B1 => n206, B2 => n104, C1
                           => n87, C2 => n242, ZN => n133);
   U168 : INV_X1 port map( A => n113, ZN => n214);
   U169 : OAI222_X1 port map( A1 => n86, A2 => n105, B1 => n207, B2 => n104, C1
                           => n81, C2 => n242, ZN => n112);
   U170 : OR4_X1 port map( A1 => SH(20), A2 => SH(19), A3 => SH(22), A4 => 
                           SH(21), ZN => n174);
   U171 : AND2_X1 port map( A1 => SH(3), A2 => n163, ZN => n161);
   U172 : OR3_X1 port map( A1 => SH(28), A2 => SH(27), A3 => SH(26), ZN => n173
                           );
   U173 : OR3_X1 port map( A1 => SH(15), A2 => SH(14), A3 => SH(13), ZN => n175
                           );
   U174 : NOR2_X1 port map( A1 => n167, A2 => n96, ZN => B(0));
   U175 : AOI21_X1 port map( B1 => n99, B2 => n176, A => n177, ZN => n167);
   U176 : NOR2_X1 port map( A1 => n130, A2 => n96, ZN => B(1));
   U177 : AOI21_X1 port map( B1 => n99, B2 => n131, A => n132, ZN => n130);
   U178 : NOR2_X1 port map( A1 => n109, A2 => n96, ZN => B(2));
   U179 : AOI21_X1 port map( B1 => n99, B2 => n110, A => n111, ZN => n109);
   U180 : AOI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => B(3));
   U181 : OAI221_X1 port map( B1 => n90, B2 => n62, C1 => n91, C2 => n64, A => 
                           n92, ZN => B(4));
   U182 : AOI222_X1 port map( A1 => n244, A2 => n75, B1 => n67, B2 => n195, C1 
                           => n69, C2 => n204, ZN => n92);
   U183 : OAI221_X1 port map( B1 => n87, B2 => n62, C1 => n88, C2 => n64, A => 
                           n89, ZN => B(5));
   U184 : AOI222_X1 port map( A1 => n244, A2 => n70, B1 => n67, B2 => n197, C1 
                           => n69, C2 => n68, ZN => n89);
   U185 : OAI221_X1 port map( B1 => n81, B2 => n62, C1 => n82, C2 => n64, A => 
                           n83, ZN => B(6));
   U186 : AOI222_X1 port map( A1 => n244, A2 => n84, B1 => n67, B2 => n199, C1 
                           => n69, C2 => n85, ZN => n83);
   U187 : OAI221_X1 port map( B1 => n76, B2 => n62, C1 => n220, C2 => n64, A =>
                           n77, ZN => B(7));
   U188 : AOI222_X1 port map( A1 => n244, A2 => n78, B1 => n67, B2 => n202, C1 
                           => n69, C2 => n79, ZN => n77);
   U189 : OAI221_X1 port map( B1 => n71, B2 => n62, C1 => n72, C2 => n64, A => 
                           n73, ZN => B(8));
   U190 : AOI222_X1 port map( A1 => n244, A2 => n74, B1 => n67, B2 => n204, C1 
                           => n69, C2 => n75, ZN => n73);
   U191 : OAI221_X1 port map( B1 => n61, B2 => n62, C1 => n63, C2 => n64, A => 
                           n65, ZN => B(9));
   U192 : AOI222_X1 port map( A1 => n244, A2 => n66, B1 => n67, B2 => n68, C1 
                           => n69, C2 => n70, ZN => n65);
   U193 : OAI221_X1 port map( B1 => n86, B2 => n62, C1 => n121, C2 => n64, A =>
                           n159, ZN => B(10));
   U194 : AOI222_X1 port map( A1 => n244, A2 => n127, B1 => n67, B2 => n85, C1 
                           => n69, C2 => n84, ZN => n159);
   U196 : OAI221_X1 port map( B1 => n126, B2 => n142, C1 => n80, C2 => n62, A 
                           => n152, ZN => B(11));
   U197 : AOI221_X1 port map( B1 => n69, B2 => n78, C1 => n67, C2 => n79, A => 
                           n153, ZN => n152);
   U198 : OAI221_X1 port map( B1 => n129, B2 => n142, C1 => n93, C2 => n62, A 
                           => n151, ZN => B(12));
   U199 : AOI222_X1 port map( A1 => n69, A2 => n74, B1 => n144, B2 => n231, C1 
                           => n67, C2 => n75, ZN => n151);
   U200 : OAI221_X1 port map( B1 => n128, B2 => n142, C1 => n206, C2 => n62, A 
                           => n146, ZN => B(13));
   U201 : AOI222_X1 port map( A1 => n69, A2 => n66, B1 => n144, B2 => n233, C1 
                           => n67, C2 => n70, ZN => n146);
   U202 : OAI221_X1 port map( B1 => n139, B2 => n142, C1 => n207, C2 => n62, A 
                           => n145, ZN => B(14));
   U203 : AOI222_X1 port map( A1 => n69, A2 => n127, B1 => n144, B2 => n234, C1
                           => n67, C2 => n84, ZN => n145);
   U204 : OAI221_X1 port map( B1 => n125, B2 => n142, C1 => n208, C2 => n62, A 
                           => n143, ZN => B(15));
   U205 : AOI222_X1 port map( A1 => n69, A2 => n219, B1 => n144, B2 => n235, C1
                           => n67, C2 => n78, ZN => n143);
   U206 : NOR2_X1 port map( A1 => n141, A2 => n246, ZN => B(16));
   U207 : NOR2_X1 port map( A1 => n134, A2 => n246, ZN => B(17));
   U208 : NOR2_X1 port map( A1 => n113, A2 => n246, ZN => B(18));
   U209 : NOR2_X1 port map( A1 => n102, A2 => n246, ZN => B(19));
   U210 : NOR2_X1 port map( A1 => n91, A2 => n246, ZN => B(20));
   U211 : NOR2_X1 port map( A1 => n88, A2 => n246, ZN => B(21));
   U212 : NOR2_X1 port map( A1 => n82, A2 => n246, ZN => B(22));
   U213 : NOR2_X1 port map( A1 => n220, A2 => n246, ZN => B(23));
   U214 : NOR2_X1 port map( A1 => n72, A2 => n246, ZN => B(24));
   U215 : NOR2_X1 port map( A1 => n63, A2 => n246, ZN => B(25));
   U216 : NOR2_X1 port map( A1 => n121, A2 => n246, ZN => B(26));
   U217 : NOR3_X1 port map( A1 => n246, A2 => SH(3), A3 => n120, ZN => B(27));
   U218 : NOR2_X1 port map( A1 => n119, A2 => n62, ZN => B(28));
   U219 : NOR2_X1 port map( A1 => n118, A2 => n62, ZN => B(29));
   U220 : NOR2_X1 port map( A1 => n108, A2 => n62, ZN => B(30));
   U221 : NOR2_X1 port map( A1 => n62, A2 => n107, ZN => B(31));

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_1 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_1;

architecture SYN_ASYNCH_FD of FD_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1020 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1020);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_2 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_2;

architecture SYN_ASYNCH_FD of FD_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1021 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1021);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_3 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_3;

architecture SYN_ASYNCH_FD of FD_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1022 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1022);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_4 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_4;

architecture SYN_ASYNCH_FD of FD_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1023 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1023);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_5 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_5;

architecture SYN_ASYNCH_FD of FD_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1024 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1024);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_6 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_6;

architecture SYN_ASYNCH_FD of FD_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1025 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1025);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_7 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_7;

architecture SYN_ASYNCH_FD of FD_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1026 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1026);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_8 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_8;

architecture SYN_ASYNCH_FD of FD_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1027 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1027);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_9 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_9;

architecture SYN_ASYNCH_FD of FD_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1028 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1028);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_10 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_10;

architecture SYN_ASYNCH_FD of FD_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1029 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1029);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_11 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_11;

architecture SYN_ASYNCH_FD of FD_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1030 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1030);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_12 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_12;

architecture SYN_ASYNCH_FD of FD_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1031 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1031);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_13 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_13;

architecture SYN_ASYNCH_FD of FD_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1032 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1032);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_14 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_14;

architecture SYN_ASYNCH_FD of FD_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1033 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1033);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_15 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_15;

architecture SYN_ASYNCH_FD of FD_15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1034 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1034);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_16 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_16;

architecture SYN_ASYNCH_FD of FD_16 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1035 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1035);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_17 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_17;

architecture SYN_ASYNCH_FD of FD_17 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1036 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1036);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_18 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_18;

architecture SYN_ASYNCH_FD of FD_18 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1037 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1037);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_19 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_19;

architecture SYN_ASYNCH_FD of FD_19 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1038 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1038);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_20 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_20;

architecture SYN_ASYNCH_FD of FD_20 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1039 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1039);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_21 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_21;

architecture SYN_ASYNCH_FD of FD_21 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1040 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1040);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_22 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_22;

architecture SYN_ASYNCH_FD of FD_22 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1041 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1041);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_23 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_23;

architecture SYN_ASYNCH_FD of FD_23 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1042 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1042);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_24 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_24;

architecture SYN_ASYNCH_FD of FD_24 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1043 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1043);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_25 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_25;

architecture SYN_ASYNCH_FD of FD_25 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1044 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1044);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_26 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_26;

architecture SYN_ASYNCH_FD of FD_26 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1045 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1045);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_27 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_27;

architecture SYN_ASYNCH_FD of FD_27 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1046 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1046);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_28 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_28;

architecture SYN_ASYNCH_FD of FD_28 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1047 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1047);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_29 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_29;

architecture SYN_ASYNCH_FD of FD_29 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1048 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1048);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_30 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_30;

architecture SYN_ASYNCH_FD of FD_30 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1049 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1049);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_31 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_31;

architecture SYN_ASYNCH_FD of FD_31 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1050 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1050);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_32 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_32;

architecture SYN_ASYNCH_FD of FD_32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1051 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1051);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_33 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_33;

architecture SYN_ASYNCH_FD of FD_33 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1052 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1052);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_34 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_34;

architecture SYN_ASYNCH_FD of FD_34 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1053 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1053);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_35 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_35;

architecture SYN_ASYNCH_FD of FD_35 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1054 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1054);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_36 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_36;

architecture SYN_ASYNCH_FD of FD_36 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1055 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1055);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_37 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_37;

architecture SYN_ASYNCH_FD of FD_37 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1056 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1056);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_38 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_38;

architecture SYN_ASYNCH_FD of FD_38 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1057 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1057);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_39 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_39;

architecture SYN_ASYNCH_FD of FD_39 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1058 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1058);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_40 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_40;

architecture SYN_ASYNCH_FD of FD_40 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1059 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1059);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_41 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_41;

architecture SYN_ASYNCH_FD of FD_41 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1060 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1060);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_42 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_42;

architecture SYN_ASYNCH_FD of FD_42 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1061 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1061);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_43 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_43;

architecture SYN_ASYNCH_FD of FD_43 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1062 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1062);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_44 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_44;

architecture SYN_ASYNCH_FD of FD_44 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1063 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1063);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_45 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_45;

architecture SYN_ASYNCH_FD of FD_45 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1064 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1064);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_46 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_46;

architecture SYN_ASYNCH_FD of FD_46 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1065 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1065);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_47 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_47;

architecture SYN_ASYNCH_FD of FD_47 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1066 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1066);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_48 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_48;

architecture SYN_ASYNCH_FD of FD_48 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1067 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1067);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_49 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_49;

architecture SYN_ASYNCH_FD of FD_49 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1068 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1068);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_50 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_50;

architecture SYN_ASYNCH_FD of FD_50 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1069 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1069);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_51 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_51;

architecture SYN_ASYNCH_FD of FD_51 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1070 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1070);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_52 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_52;

architecture SYN_ASYNCH_FD of FD_52 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1071 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1071);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_53 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_53;

architecture SYN_ASYNCH_FD of FD_53 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1072 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1072);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_54 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_54;

architecture SYN_ASYNCH_FD of FD_54 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1073 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1073);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_55 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_55;

architecture SYN_ASYNCH_FD of FD_55 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1074 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1074);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_56 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_56;

architecture SYN_ASYNCH_FD of FD_56 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1075 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1075);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_57 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_57;

architecture SYN_ASYNCH_FD of FD_57 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1076 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1076);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_58 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_58;

architecture SYN_ASYNCH_FD of FD_58 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1077 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1077);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_59 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_59;

architecture SYN_ASYNCH_FD of FD_59 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1078 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1078);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_60 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_60;

architecture SYN_ASYNCH_FD of FD_60 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1079 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1079);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_61 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_61;

architecture SYN_ASYNCH_FD of FD_61 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1080 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1080);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_62 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_62;

architecture SYN_ASYNCH_FD of FD_62 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1081 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1081);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_63 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_63;

architecture SYN_ASYNCH_FD of FD_63 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1082 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1082);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_64 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_64;

architecture SYN_ASYNCH_FD of FD_64 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1083 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1083);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_65 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_65;

architecture SYN_ASYNCH_FD of FD_65 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1084 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1084);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_66 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_66;

architecture SYN_ASYNCH_FD of FD_66 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1085 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1085);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_67 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_67;

architecture SYN_ASYNCH_FD of FD_67 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1086 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1086);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_68 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_68;

architecture SYN_ASYNCH_FD of FD_68 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1087 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1087);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_69 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_69;

architecture SYN_ASYNCH_FD of FD_69 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1088 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1088);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_70 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_70;

architecture SYN_ASYNCH_FD of FD_70 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1089 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1089);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_71 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_71;

architecture SYN_ASYNCH_FD of FD_71 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1090 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1090);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_72 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_72;

architecture SYN_ASYNCH_FD of FD_72 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1091 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1091);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_73 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_73;

architecture SYN_ASYNCH_FD of FD_73 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1092 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1092);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_74 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_74;

architecture SYN_ASYNCH_FD of FD_74 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1093 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1093);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_75 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_75;

architecture SYN_ASYNCH_FD of FD_75 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1094 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1094);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_76 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_76;

architecture SYN_ASYNCH_FD of FD_76 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1095 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1095);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_77 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_77;

architecture SYN_ASYNCH_FD of FD_77 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1096 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1096);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_78 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_78;

architecture SYN_ASYNCH_FD of FD_78 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1097 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1097);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_79 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_79;

architecture SYN_ASYNCH_FD of FD_79 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1098 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1098);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_80 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_80;

architecture SYN_ASYNCH_FD of FD_80 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1099 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1099);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_81 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_81;

architecture SYN_ASYNCH_FD of FD_81 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1100 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1100);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_82 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_82;

architecture SYN_ASYNCH_FD of FD_82 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1101 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1101);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_83 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_83;

architecture SYN_ASYNCH_FD of FD_83 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1102 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1102);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_84 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_84;

architecture SYN_ASYNCH_FD of FD_84 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1103 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1103);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_85 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_85;

architecture SYN_ASYNCH_FD of FD_85 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1104 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1104);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_86 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_86;

architecture SYN_ASYNCH_FD of FD_86 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1105 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1105);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_87 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_87;

architecture SYN_ASYNCH_FD of FD_87 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1106 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1106);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_88 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_88;

architecture SYN_ASYNCH_FD of FD_88 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1107 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1107);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_89 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_89;

architecture SYN_ASYNCH_FD of FD_89 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1108 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1108);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_90 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_90;

architecture SYN_ASYNCH_FD of FD_90 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1109 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1109);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_91 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_91;

architecture SYN_ASYNCH_FD of FD_91 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1110 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1110);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_92 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_92;

architecture SYN_ASYNCH_FD of FD_92 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1111 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1111);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_93 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_93;

architecture SYN_ASYNCH_FD of FD_93 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1112 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1112);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_94 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_94;

architecture SYN_ASYNCH_FD of FD_94 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1113 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1113);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_95 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_95;

architecture SYN_ASYNCH_FD of FD_95 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1114 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1114);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_96 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_96;

architecture SYN_ASYNCH_FD of FD_96 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1115 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1115);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_97 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_97;

architecture SYN_ASYNCH_FD of FD_97 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1116 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1116);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_98 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_98;

architecture SYN_ASYNCH_FD of FD_98 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1117 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1117);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_99 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_99;

architecture SYN_ASYNCH_FD of FD_99 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1118 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1118);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_100 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_100;

architecture SYN_ASYNCH_FD of FD_100 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1119 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1119);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_101 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_101;

architecture SYN_ASYNCH_FD of FD_101 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1120 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1120);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_102 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_102;

architecture SYN_ASYNCH_FD of FD_102 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1121 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1121);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_103 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_103;

architecture SYN_ASYNCH_FD of FD_103 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1122 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1122);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_104 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_104;

architecture SYN_ASYNCH_FD of FD_104 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1123 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1123);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_105 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_105;

architecture SYN_ASYNCH_FD of FD_105 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1124 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1124);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_106 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_106;

architecture SYN_ASYNCH_FD of FD_106 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1125 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1125);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_107 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_107;

architecture SYN_ASYNCH_FD of FD_107 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1126 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1126);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_108 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_108;

architecture SYN_ASYNCH_FD of FD_108 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1127 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1127);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_109 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_109;

architecture SYN_ASYNCH_FD of FD_109 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1128 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1128);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_110 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_110;

architecture SYN_ASYNCH_FD of FD_110 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1129 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1129);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_111 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_111;

architecture SYN_ASYNCH_FD of FD_111 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1130 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1130);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_112 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_112;

architecture SYN_ASYNCH_FD of FD_112 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1131 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1131);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_113 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_113;

architecture SYN_ASYNCH_FD of FD_113 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1132 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1132);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_114 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_114;

architecture SYN_ASYNCH_FD of FD_114 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1133 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1133);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_115 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_115;

architecture SYN_ASYNCH_FD of FD_115 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1134 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1134);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_116 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_116;

architecture SYN_ASYNCH_FD of FD_116 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1135 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1135);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_117 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_117;

architecture SYN_ASYNCH_FD of FD_117 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1136 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1136);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_118 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_118;

architecture SYN_ASYNCH_FD of FD_118 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1137 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1137);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_119 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_119;

architecture SYN_ASYNCH_FD of FD_119 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1138 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1138);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_120 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_120;

architecture SYN_ASYNCH_FD of FD_120 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1139 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1139);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_121 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_121;

architecture SYN_ASYNCH_FD of FD_121 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1140 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1140);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_122 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_122;

architecture SYN_ASYNCH_FD of FD_122 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1141 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1141);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_123 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_123;

architecture SYN_ASYNCH_FD of FD_123 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1142 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1142);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_124 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_124;

architecture SYN_ASYNCH_FD of FD_124 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1143 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1143);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_125 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_125;

architecture SYN_ASYNCH_FD of FD_125 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1144 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1144);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_126 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_126;

architecture SYN_ASYNCH_FD of FD_126 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1145 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1145);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_127 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_127;

architecture SYN_ASYNCH_FD of FD_127 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1146 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1146);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_128 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_128;

architecture SYN_ASYNCH_FD of FD_128 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1147 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1147);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_129 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_129;

architecture SYN_ASYNCH_FD of FD_129 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1148 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1148);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_130 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_130;

architecture SYN_ASYNCH_FD of FD_130 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1149 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1149);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_131 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_131;

architecture SYN_ASYNCH_FD of FD_131 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1150 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1150);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_132 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_132;

architecture SYN_ASYNCH_FD of FD_132 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1151 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1151);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_133 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_133;

architecture SYN_ASYNCH_FD of FD_133 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1152 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1152);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_134 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_134;

architecture SYN_ASYNCH_FD of FD_134 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1153 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1153);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_135 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_135;

architecture SYN_ASYNCH_FD of FD_135 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1154 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1154);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_136 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_136;

architecture SYN_ASYNCH_FD of FD_136 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1155 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1155);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_137 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_137;

architecture SYN_ASYNCH_FD of FD_137 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1156 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1156);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_138 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_138;

architecture SYN_ASYNCH_FD of FD_138 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1157 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1157);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_139 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_139;

architecture SYN_ASYNCH_FD of FD_139 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1158 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1158);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_140 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_140;

architecture SYN_ASYNCH_FD of FD_140 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1159 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1159);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_141 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_141;

architecture SYN_ASYNCH_FD of FD_141 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1160 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1160);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_142 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_142;

architecture SYN_ASYNCH_FD of FD_142 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1161 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1161);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_143 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_143;

architecture SYN_ASYNCH_FD of FD_143 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1162 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1162);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_144 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_144;

architecture SYN_ASYNCH_FD of FD_144 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1163 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1163);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_145 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_145;

architecture SYN_ASYNCH_FD of FD_145 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1164 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1164);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_146 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_146;

architecture SYN_ASYNCH_FD of FD_146 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1165 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1165);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_147 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_147;

architecture SYN_ASYNCH_FD of FD_147 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1166 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1166);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_148 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_148;

architecture SYN_ASYNCH_FD of FD_148 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1167 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1167);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_149 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_149;

architecture SYN_ASYNCH_FD of FD_149 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1168 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1168);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_150 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_150;

architecture SYN_ASYNCH_FD of FD_150 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1169 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1169);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_151 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_151;

architecture SYN_ASYNCH_FD of FD_151 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1170 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1170);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_152 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_152;

architecture SYN_ASYNCH_FD of FD_152 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1171 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1171);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_153 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_153;

architecture SYN_ASYNCH_FD of FD_153 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1172 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1172);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_154 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_154;

architecture SYN_ASYNCH_FD of FD_154 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1173 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1173);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_155 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_155;

architecture SYN_ASYNCH_FD of FD_155 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1174 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1174);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_156 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_156;

architecture SYN_ASYNCH_FD of FD_156 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1175 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1175);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_157 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_157;

architecture SYN_ASYNCH_FD of FD_157 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1176 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1176);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_158 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_158;

architecture SYN_ASYNCH_FD of FD_158 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1177 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1177);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_159 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_159;

architecture SYN_ASYNCH_FD of FD_159 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1178 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1178);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_160 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_160;

architecture SYN_ASYNCH_FD of FD_160 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1179 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1179);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_161 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_161;

architecture SYN_ASYNCH_FD of FD_161 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1180 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1180);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_162 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_162;

architecture SYN_ASYNCH_FD of FD_162 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1181 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1181);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_163 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_163;

architecture SYN_ASYNCH_FD of FD_163 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1182 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1182);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_164 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_164;

architecture SYN_ASYNCH_FD of FD_164 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1183 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1183);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_165 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_165;

architecture SYN_ASYNCH_FD of FD_165 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1184 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1184);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_166 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_166;

architecture SYN_ASYNCH_FD of FD_166 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1185 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1185);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_167 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_167;

architecture SYN_ASYNCH_FD of FD_167 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1186 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1186);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_168 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_168;

architecture SYN_ASYNCH_FD of FD_168 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1187 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1187);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_169 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_169;

architecture SYN_ASYNCH_FD of FD_169 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1188 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1188);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_170 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_170;

architecture SYN_ASYNCH_FD of FD_170 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1189 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1189);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_171 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_171;

architecture SYN_ASYNCH_FD of FD_171 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1190 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1190);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_172 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_172;

architecture SYN_ASYNCH_FD of FD_172 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1191 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1191);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_173 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_173;

architecture SYN_ASYNCH_FD of FD_173 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1192 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1192);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_174 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_174;

architecture SYN_ASYNCH_FD of FD_174 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1193 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1193);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_175 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_175;

architecture SYN_ASYNCH_FD of FD_175 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1194 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1194);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_176 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_176;

architecture SYN_ASYNCH_FD of FD_176 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1195 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1195);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_177 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_177;

architecture SYN_ASYNCH_FD of FD_177 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1196 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1196);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_178 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_178;

architecture SYN_ASYNCH_FD of FD_178 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1197 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1197);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_179 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_179;

architecture SYN_ASYNCH_FD of FD_179 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1198 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1198);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_180 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_180;

architecture SYN_ASYNCH_FD of FD_180 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1199 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1199);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_181 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_181;

architecture SYN_ASYNCH_FD of FD_181 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1200 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1200);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_182 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_182;

architecture SYN_ASYNCH_FD of FD_182 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1201 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1201);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_183 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_183;

architecture SYN_ASYNCH_FD of FD_183 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1202 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1202);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_184 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_184;

architecture SYN_ASYNCH_FD of FD_184 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1203 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1203);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_185 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_185;

architecture SYN_ASYNCH_FD of FD_185 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1204 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1204);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_186 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_186;

architecture SYN_ASYNCH_FD of FD_186 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1205 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1205);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_187 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_187;

architecture SYN_ASYNCH_FD of FD_187 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1206 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1206);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_188 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_188;

architecture SYN_ASYNCH_FD of FD_188 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1207 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1207);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_189 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_189;

architecture SYN_ASYNCH_FD of FD_189 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1208 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1208);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_190 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_190;

architecture SYN_ASYNCH_FD of FD_190 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1209 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1209);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_191 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_191;

architecture SYN_ASYNCH_FD of FD_191 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1210 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1210);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_192 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_192;

architecture SYN_ASYNCH_FD of FD_192 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1211 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1211);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_193 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_193;

architecture SYN_ASYNCH_FD of FD_193 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1212 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1212);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_194 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_194;

architecture SYN_ASYNCH_FD of FD_194 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1213 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1213);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_195 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_195;

architecture SYN_ASYNCH_FD of FD_195 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1214 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1214);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_196 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_196;

architecture SYN_ASYNCH_FD of FD_196 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1215 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1215);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_197 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_197;

architecture SYN_ASYNCH_FD of FD_197 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1216 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1216);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_198 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_198;

architecture SYN_ASYNCH_FD of FD_198 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1217 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1217);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_199 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_199;

architecture SYN_ASYNCH_FD of FD_199 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1218 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1218);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_200 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_200;

architecture SYN_ASYNCH_FD of FD_200 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1219 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1219);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_201 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_201;

architecture SYN_ASYNCH_FD of FD_201 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1220 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1220);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_202 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_202;

architecture SYN_ASYNCH_FD of FD_202 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1221 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1221);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_203 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_203;

architecture SYN_ASYNCH_FD of FD_203 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1222 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1222);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_204 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_204;

architecture SYN_ASYNCH_FD of FD_204 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1223 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1223);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_205 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_205;

architecture SYN_ASYNCH_FD of FD_205 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1224 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1224);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_206 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_206;

architecture SYN_ASYNCH_FD of FD_206 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1225 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1225);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_207 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_207;

architecture SYN_ASYNCH_FD of FD_207 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1226 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1226);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_208 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_208;

architecture SYN_ASYNCH_FD of FD_208 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1227 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1227);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_209 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_209;

architecture SYN_ASYNCH_FD of FD_209 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1228 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1228);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_210 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_210;

architecture SYN_ASYNCH_FD of FD_210 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1229 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1229);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_211 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_211;

architecture SYN_ASYNCH_FD of FD_211 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1230 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1230);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_212 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_212;

architecture SYN_ASYNCH_FD of FD_212 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1231 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1231);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_213 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_213;

architecture SYN_ASYNCH_FD of FD_213 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1232 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1232);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_214 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_214;

architecture SYN_ASYNCH_FD of FD_214 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1233 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1233);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_215 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_215;

architecture SYN_ASYNCH_FD of FD_215 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1234 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1234);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_216 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_216;

architecture SYN_ASYNCH_FD of FD_216 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1235 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1235);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_217 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_217;

architecture SYN_ASYNCH_FD of FD_217 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1236 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1236);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_218 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_218;

architecture SYN_ASYNCH_FD of FD_218 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1237 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1237);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_219 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_219;

architecture SYN_ASYNCH_FD of FD_219 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1238 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1238);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_220 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_220;

architecture SYN_ASYNCH_FD of FD_220 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1239 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1239);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_221 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_221;

architecture SYN_ASYNCH_FD of FD_221 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1240 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1240);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_222 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_222;

architecture SYN_ASYNCH_FD of FD_222 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1241 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1241);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_223 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_223;

architecture SYN_ASYNCH_FD of FD_223 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1242 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1242);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_224 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_224;

architecture SYN_ASYNCH_FD of FD_224 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1243 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1243);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_225 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_225;

architecture SYN_ASYNCH_FD of FD_225 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1244 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1244);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_226 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_226;

architecture SYN_ASYNCH_FD of FD_226 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1245 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1245);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_227 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_227;

architecture SYN_ASYNCH_FD of FD_227 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1246 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1246);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_228 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_228;

architecture SYN_ASYNCH_FD of FD_228 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1247 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1247);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_229 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_229;

architecture SYN_ASYNCH_FD of FD_229 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1248 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1248);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_230 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_230;

architecture SYN_ASYNCH_FD of FD_230 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1249 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1249);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_231 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_231;

architecture SYN_ASYNCH_FD of FD_231 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1250 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1250);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_232 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_232;

architecture SYN_ASYNCH_FD of FD_232 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1251 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1251);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_233 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_233;

architecture SYN_ASYNCH_FD of FD_233 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1252 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1252);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_234 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_234;

architecture SYN_ASYNCH_FD of FD_234 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1253 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1253);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_235 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_235;

architecture SYN_ASYNCH_FD of FD_235 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1254 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1254);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_236 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_236;

architecture SYN_ASYNCH_FD of FD_236 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1255 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1255);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_237 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_237;

architecture SYN_ASYNCH_FD of FD_237 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1256 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1256);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_238 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_238;

architecture SYN_ASYNCH_FD of FD_238 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1257 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1257);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_239 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_239;

architecture SYN_ASYNCH_FD of FD_239 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1258 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1258);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_240 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_240;

architecture SYN_ASYNCH_FD of FD_240 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1259 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1259);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_241 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_241;

architecture SYN_ASYNCH_FD of FD_241 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1260 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1260);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_242 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_242;

architecture SYN_ASYNCH_FD of FD_242 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1261 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1261);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_243 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_243;

architecture SYN_ASYNCH_FD of FD_243 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1262 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1262);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_244 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_244;

architecture SYN_ASYNCH_FD of FD_244 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1263 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1263);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_245 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_245;

architecture SYN_ASYNCH_FD of FD_245 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1264 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1264);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_246 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_246;

architecture SYN_ASYNCH_FD of FD_246 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1265 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1265);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_247 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_247;

architecture SYN_ASYNCH_FD of FD_247 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1266 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1266);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_248 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_248;

architecture SYN_ASYNCH_FD of FD_248 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1267 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1267);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_249 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_249;

architecture SYN_ASYNCH_FD of FD_249 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1268 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1268);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_250 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_250;

architecture SYN_ASYNCH_FD of FD_250 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1269 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1269);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_251 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_251;

architecture SYN_ASYNCH_FD of FD_251 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1270 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1270);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_252 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_252;

architecture SYN_ASYNCH_FD of FD_252 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1271 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1271);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_253 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_253;

architecture SYN_ASYNCH_FD of FD_253 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1272 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1272);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_254 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_254;

architecture SYN_ASYNCH_FD of FD_254 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1273 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1273);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_255 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_255;

architecture SYN_ASYNCH_FD of FD_255 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1274 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1274);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_256 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_256;

architecture SYN_ASYNCH_FD of FD_256 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1275 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1275);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_257 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_257;

architecture SYN_ASYNCH_FD of FD_257 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1276 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1276);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_258 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_258;

architecture SYN_ASYNCH_FD of FD_258 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1277 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1277);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_259 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_259;

architecture SYN_ASYNCH_FD of FD_259 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1278 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1278);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_260 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_260;

architecture SYN_ASYNCH_FD of FD_260 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1279 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1279);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_261 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_261;

architecture SYN_ASYNCH_FD of FD_261 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1280 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1280);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_262 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_262;

architecture SYN_ASYNCH_FD of FD_262 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1281 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1281);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_263 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_263;

architecture SYN_ASYNCH_FD of FD_263 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1282 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1282);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_264 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_264;

architecture SYN_ASYNCH_FD of FD_264 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1283 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1283);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_265 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_265;

architecture SYN_ASYNCH_FD of FD_265 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1284 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1284);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_266 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_266;

architecture SYN_ASYNCH_FD of FD_266 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1285 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1285);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_267 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_267;

architecture SYN_ASYNCH_FD of FD_267 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1286 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1286);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_268 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_268;

architecture SYN_ASYNCH_FD of FD_268 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1287 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1287);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_269 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_269;

architecture SYN_ASYNCH_FD of FD_269 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1288 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1288);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_270 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_270;

architecture SYN_ASYNCH_FD of FD_270 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1289 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1289);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_271 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_271;

architecture SYN_ASYNCH_FD of FD_271 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1290 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1290);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_272 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_272;

architecture SYN_ASYNCH_FD of FD_272 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1291 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1291);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_273 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_273;

architecture SYN_ASYNCH_FD of FD_273 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1292 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1292);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_274 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_274;

architecture SYN_ASYNCH_FD of FD_274 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1293 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1293);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_275 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_275;

architecture SYN_ASYNCH_FD of FD_275 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1294 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1294);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_276 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_276;

architecture SYN_ASYNCH_FD of FD_276 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1295 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1295);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_277 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_277;

architecture SYN_ASYNCH_FD of FD_277 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1296 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1296);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_278 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_278;

architecture SYN_ASYNCH_FD of FD_278 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1297 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1297);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_279 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_279;

architecture SYN_ASYNCH_FD of FD_279 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1298 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1298);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_280 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_280;

architecture SYN_ASYNCH_FD of FD_280 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1299 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1299);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_281 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_281;

architecture SYN_ASYNCH_FD of FD_281 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1300 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1300);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_282 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_282;

architecture SYN_ASYNCH_FD of FD_282 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1301 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1301);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_283 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_283;

architecture SYN_ASYNCH_FD of FD_283 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1302 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1302);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_284 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_284;

architecture SYN_ASYNCH_FD of FD_284 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1303 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1303);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_285 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_285;

architecture SYN_ASYNCH_FD of FD_285 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1304 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1304);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_286 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_286;

architecture SYN_ASYNCH_FD of FD_286 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1305 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1305);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_287 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_287;

architecture SYN_ASYNCH_FD of FD_287 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1306 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1306);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_288 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_288;

architecture SYN_ASYNCH_FD of FD_288 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1307 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1307);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_289 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_289;

architecture SYN_ASYNCH_FD of FD_289 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1308 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1308);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_290 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_290;

architecture SYN_ASYNCH_FD of FD_290 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1309 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1309);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_291 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_291;

architecture SYN_ASYNCH_FD of FD_291 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1310 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1310);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_292 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_292;

architecture SYN_ASYNCH_FD of FD_292 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1311 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1311);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_293 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_293;

architecture SYN_ASYNCH_FD of FD_293 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1312 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1312);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_294 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_294;

architecture SYN_ASYNCH_FD of FD_294 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1313 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1313);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_295 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_295;

architecture SYN_ASYNCH_FD of FD_295 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1314 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1314);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_296 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_296;

architecture SYN_ASYNCH_FD of FD_296 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1315 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1315);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_297 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_297;

architecture SYN_ASYNCH_FD of FD_297 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1316 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1316);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_298 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_298;

architecture SYN_ASYNCH_FD of FD_298 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1317 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1317);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_299 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_299;

architecture SYN_ASYNCH_FD of FD_299 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1318 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1318);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_300 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_300;

architecture SYN_ASYNCH_FD of FD_300 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1319 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1319);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_301 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_301;

architecture SYN_ASYNCH_FD of FD_301 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1320 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1320);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_302 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_302;

architecture SYN_ASYNCH_FD of FD_302 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1321 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1321);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_303 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_303;

architecture SYN_ASYNCH_FD of FD_303 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1322 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1322);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_304 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_304;

architecture SYN_ASYNCH_FD of FD_304 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1323 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1323);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_305 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_305;

architecture SYN_ASYNCH_FD of FD_305 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1324 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1324);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_306 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_306;

architecture SYN_ASYNCH_FD of FD_306 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1325 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1325);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_307 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_307;

architecture SYN_ASYNCH_FD of FD_307 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1326 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1326);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_308 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_308;

architecture SYN_ASYNCH_FD of FD_308 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1327 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1327);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_309 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_309;

architecture SYN_ASYNCH_FD of FD_309 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1328 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1328);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_310 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_310;

architecture SYN_ASYNCH_FD of FD_310 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1329 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1329);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_311 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_311;

architecture SYN_ASYNCH_FD of FD_311 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1330 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1330);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_312 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_312;

architecture SYN_ASYNCH_FD of FD_312 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1331 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1331);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_313 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_313;

architecture SYN_ASYNCH_FD of FD_313 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1332 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1332);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_314 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_314;

architecture SYN_ASYNCH_FD of FD_314 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1333 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1333);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_315 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_315;

architecture SYN_ASYNCH_FD of FD_315 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1334 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1334);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_316 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_316;

architecture SYN_ASYNCH_FD of FD_316 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1335 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1335);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_317 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_317;

architecture SYN_ASYNCH_FD of FD_317 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1336 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1336);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_318 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_318;

architecture SYN_ASYNCH_FD of FD_318 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1337 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1337);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_319 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_319;

architecture SYN_ASYNCH_FD of FD_319 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1338 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1338);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_320 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_320;

architecture SYN_ASYNCH_FD of FD_320 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1339 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1339);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_321 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_321;

architecture SYN_ASYNCH_FD of FD_321 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1340 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1340);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_322 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_322;

architecture SYN_ASYNCH_FD of FD_322 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1341 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1341);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_323 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_323;

architecture SYN_ASYNCH_FD of FD_323 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1342 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1342);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_324 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_324;

architecture SYN_ASYNCH_FD of FD_324 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1343 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1343);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_325 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_325;

architecture SYN_ASYNCH_FD of FD_325 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1344 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1344);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_326 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_326;

architecture SYN_ASYNCH_FD of FD_326 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1345 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1345);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_327 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_327;

architecture SYN_ASYNCH_FD of FD_327 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1346 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1346);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_328 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_328;

architecture SYN_ASYNCH_FD of FD_328 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1347 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1347);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_329 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_329;

architecture SYN_ASYNCH_FD of FD_329 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1348 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1348);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_330 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_330;

architecture SYN_ASYNCH_FD of FD_330 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1349 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1349);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_331 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_331;

architecture SYN_ASYNCH_FD of FD_331 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1350 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1350);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_332 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_332;

architecture SYN_ASYNCH_FD of FD_332 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1351 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1351);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_333 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_333;

architecture SYN_ASYNCH_FD of FD_333 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1352 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1352);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_334 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_334;

architecture SYN_ASYNCH_FD of FD_334 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1353 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1353);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_335 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_335;

architecture SYN_ASYNCH_FD of FD_335 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1354 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1354);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_336 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_336;

architecture SYN_ASYNCH_FD of FD_336 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1355 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1355);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_337 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_337;

architecture SYN_ASYNCH_FD of FD_337 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1356 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1356);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_338 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_338;

architecture SYN_ASYNCH_FD of FD_338 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1357 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1357);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_339 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_339;

architecture SYN_ASYNCH_FD of FD_339 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1358 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1358);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_340 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_340;

architecture SYN_ASYNCH_FD of FD_340 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1359 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1359);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_341 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_341;

architecture SYN_ASYNCH_FD of FD_341 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1360 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1360);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_342 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_342;

architecture SYN_ASYNCH_FD of FD_342 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1361 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1361);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_343 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_343;

architecture SYN_ASYNCH_FD of FD_343 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1362 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1362);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_344 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_344;

architecture SYN_ASYNCH_FD of FD_344 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1363 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1363);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_345 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_345;

architecture SYN_ASYNCH_FD of FD_345 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1364 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1364);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_346 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_346;

architecture SYN_ASYNCH_FD of FD_346 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1365 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1365);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_347 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_347;

architecture SYN_ASYNCH_FD of FD_347 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1366 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1366);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_348 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_348;

architecture SYN_ASYNCH_FD of FD_348 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1367 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1367);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_349 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_349;

architecture SYN_ASYNCH_FD of FD_349 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1368 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1368);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_350 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_350;

architecture SYN_ASYNCH_FD of FD_350 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1369 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1369);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_351 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_351;

architecture SYN_ASYNCH_FD of FD_351 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1370 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1370);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_352 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_352;

architecture SYN_ASYNCH_FD of FD_352 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1371 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1371);
   U2 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n2);
   U3 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_1;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U5 : MUX2_X1 port map( A => B(4), B => A(4), S => S, Z => Y(4));
   U6 : MUX2_X1 port map( A => B(5), B => A(5), S => S, Z => Y(5));
   U7 : MUX2_X1 port map( A => B(6), B => A(6), S => S, Z => Y(6));
   U8 : MUX2_X1 port map( A => B(7), B => A(7), S => S, Z => Y(7));
   U9 : MUX2_X1 port map( A => B(8), B => A(8), S => S, Z => Y(8));
   U10 : MUX2_X1 port map( A => B(9), B => A(9), S => S, Z => Y(9));
   U11 : MUX2_X1 port map( A => B(10), B => A(10), S => S, Z => Y(10));
   U12 : MUX2_X1 port map( A => B(11), B => A(11), S => S, Z => Y(11));
   U13 : MUX2_X1 port map( A => B(12), B => A(12), S => S, Z => Y(12));
   U14 : MUX2_X1 port map( A => B(13), B => A(13), S => S, Z => Y(13));
   U15 : MUX2_X1 port map( A => B(14), B => A(14), S => S, Z => Y(14));
   U16 : MUX2_X1 port map( A => B(15), B => A(15), S => S, Z => Y(15));
   U17 : MUX2_X1 port map( A => B(16), B => A(16), S => S, Z => Y(16));
   U18 : MUX2_X1 port map( A => B(17), B => A(17), S => S, Z => Y(17));
   U19 : MUX2_X1 port map( A => B(18), B => A(18), S => S, Z => Y(18));
   U20 : MUX2_X1 port map( A => B(19), B => A(19), S => S, Z => Y(19));
   U21 : MUX2_X1 port map( A => B(20), B => A(20), S => S, Z => Y(20));
   U22 : MUX2_X1 port map( A => B(21), B => A(21), S => S, Z => Y(21));
   U23 : MUX2_X1 port map( A => B(22), B => A(22), S => S, Z => Y(22));
   U24 : MUX2_X1 port map( A => B(23), B => A(23), S => S, Z => Y(23));
   U25 : MUX2_X1 port map( A => B(24), B => A(24), S => S, Z => Y(24));
   U26 : MUX2_X1 port map( A => B(25), B => A(25), S => S, Z => Y(25));
   U27 : MUX2_X1 port map( A => B(26), B => A(26), S => S, Z => Y(26));
   U28 : MUX2_X1 port map( A => B(27), B => A(27), S => S, Z => Y(27));
   U29 : MUX2_X1 port map( A => B(28), B => A(28), S => S, Z => Y(28));
   U30 : MUX2_X1 port map( A => B(29), B => A(29), S => S, Z => Y(29));
   U31 : MUX2_X1 port map( A => B(30), B => A(30), S => S, Z => Y(30));
   U32 : MUX2_X1 port map( A => B(31), B => A(31), S => S, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_1 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_1;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_3
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_4
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_5
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_6
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_7
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_8
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_9
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_10
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_11
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_12
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_13
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_14
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_15
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_16
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_17
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_18
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_19
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_20
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_21
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_22
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_23
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_24
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_25
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_26
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_27
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_28
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_29
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_30
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_31
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_32
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_32 port map( D => data_in(0), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_31 port map( D => data_in(1), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_30 port map( D => data_in(2), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_29 port map( D => data_in(3), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_28 port map( D => data_in(4), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_27 port map( D => data_in(5), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_26 port map( D => data_in(6), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_25 port map( D => data_in(7), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_24 port map( D => data_in(8), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_23 port map( D => data_in(9), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_22 port map( D => data_in(10), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_21 port map( D => data_in(11), CK => n14, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_20 port map( D => data_in(12), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(12));
   FF_13 : FD_19 port map( D => data_in(13), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(13));
   FF_14 : FD_18 port map( D => data_in(14), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(14));
   FF_15 : FD_17 port map( D => data_in(15), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(15));
   FF_16 : FD_16 port map( D => data_in(16), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(16));
   FF_17 : FD_15 port map( D => data_in(17), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(17));
   FF_18 : FD_14 port map( D => data_in(18), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(18));
   FF_19 : FD_13 port map( D => data_in(19), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(19));
   FF_20 : FD_12 port map( D => data_in(20), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(20));
   FF_21 : FD_11 port map( D => data_in(21), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(21));
   FF_22 : FD_10 port map( D => data_in(22), CK => n15, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(22));
   FF_23 : FD_9 port map( D => data_in(23), CK => n15, RESET => n10, ENABLE => 
                           ENABLE, Q => data_out(23));
   FF_24 : FD_8 port map( D => data_in(24), CK => n15, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(24));
   FF_25 : FD_7 port map( D => data_in(25), CK => n15, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(25));
   FF_26 : FD_6 port map( D => data_in(26), CK => n15, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(26));
   FF_27 : FD_5 port map( D => data_in(27), CK => n15, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(27));
   FF_28 : FD_4 port map( D => data_in(28), CK => n15, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(28));
   FF_29 : FD_3 port map( D => data_in(29), CK => n15, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(29));
   FF_30 : FD_2 port map( D => data_in(30), CK => n15, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(30));
   FF_31 : FD_1 port map( D => data_in(31), CK => n15, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => CK, Z => n16);
   U3 : BUF_X1 port map( A => n12, Z => n9);
   U4 : BUF_X1 port map( A => n12, Z => n10);
   U5 : BUF_X1 port map( A => n12, Z => n11);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_2 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_2;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_33
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_34
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_35
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_36
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_37
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_38
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_39
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_40
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_41
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_42
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_43
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_44
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_45
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_46
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_47
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_48
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_49
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_50
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_51
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_52
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_53
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_54
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_55
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_56
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_57
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_58
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_59
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_60
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_61
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_62
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_63
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_64
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_64 port map( D => data_in(0), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_63 port map( D => data_in(1), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_62 port map( D => data_in(2), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_61 port map( D => data_in(3), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_60 port map( D => data_in(4), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_59 port map( D => data_in(5), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_58 port map( D => data_in(6), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_57 port map( D => data_in(7), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_56 port map( D => data_in(8), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_55 port map( D => data_in(9), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_54 port map( D => data_in(10), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_53 port map( D => data_in(11), CK => n14, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_52 port map( D => data_in(12), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(12));
   FF_13 : FD_51 port map( D => data_in(13), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(13));
   FF_14 : FD_50 port map( D => data_in(14), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(14));
   FF_15 : FD_49 port map( D => data_in(15), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(15));
   FF_16 : FD_48 port map( D => data_in(16), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(16));
   FF_17 : FD_47 port map( D => data_in(17), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(17));
   FF_18 : FD_46 port map( D => data_in(18), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(18));
   FF_19 : FD_45 port map( D => data_in(19), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(19));
   FF_20 : FD_44 port map( D => data_in(20), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(20));
   FF_21 : FD_43 port map( D => data_in(21), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(21));
   FF_22 : FD_42 port map( D => data_in(22), CK => n15, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(22));
   FF_23 : FD_41 port map( D => data_in(23), CK => n15, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(23));
   FF_24 : FD_40 port map( D => data_in(24), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(24));
   FF_25 : FD_39 port map( D => data_in(25), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(25));
   FF_26 : FD_38 port map( D => data_in(26), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(26));
   FF_27 : FD_37 port map( D => data_in(27), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(27));
   FF_28 : FD_36 port map( D => data_in(28), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(28));
   FF_29 : FD_35 port map( D => data_in(29), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(29));
   FF_30 : FD_34 port map( D => data_in(30), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(30));
   FF_31 : FD_33 port map( D => data_in(31), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => CK, Z => n16);
   U3 : BUF_X1 port map( A => n12, Z => n9);
   U4 : BUF_X1 port map( A => n12, Z => n10);
   U5 : BUF_X1 port map( A => n12, Z => n11);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_2;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U2 : MUX2_X1 port map( A => B(4), B => A(4), S => S, Z => Y(4));
   U3 : MUX2_X1 port map( A => B(5), B => A(5), S => S, Z => Y(5));
   U4 : MUX2_X1 port map( A => B(7), B => A(7), S => S, Z => Y(7));
   U5 : MUX2_X1 port map( A => B(9), B => A(9), S => S, Z => Y(9));
   U6 : MUX2_X1 port map( A => B(11), B => A(11), S => S, Z => Y(11));
   U7 : MUX2_X1 port map( A => B(17), B => A(17), S => S, Z => Y(17));
   U8 : MUX2_X1 port map( A => B(19), B => A(19), S => S, Z => Y(19));
   U9 : MUX2_X1 port map( A => B(21), B => A(21), S => S, Z => Y(21));
   U10 : MUX2_X1 port map( A => B(30), B => A(30), S => S, Z => Y(30));
   U11 : MUX2_X1 port map( A => B(31), B => A(31), S => S, Z => Y(31));
   U12 : MUX2_X1 port map( A => B(29), B => A(29), S => S, Z => Y(29));
   U13 : MUX2_X1 port map( A => B(28), B => A(28), S => S, Z => Y(28));
   U14 : MUX2_X1 port map( A => B(27), B => A(27), S => S, Z => Y(27));
   U15 : MUX2_X1 port map( A => B(26), B => A(26), S => S, Z => Y(26));
   U16 : MUX2_X1 port map( A => B(25), B => A(25), S => S, Z => Y(25));
   U17 : MUX2_X1 port map( A => B(24), B => A(24), S => S, Z => Y(24));
   U18 : MUX2_X1 port map( A => B(23), B => A(23), S => S, Z => Y(23));
   U19 : MUX2_X1 port map( A => B(22), B => A(22), S => S, Z => Y(22));
   U20 : MUX2_X1 port map( A => B(20), B => A(20), S => S, Z => Y(20));
   U21 : MUX2_X1 port map( A => B(18), B => A(18), S => S, Z => Y(18));
   U22 : MUX2_X1 port map( A => B(16), B => A(16), S => S, Z => Y(16));
   U23 : MUX2_X1 port map( A => B(15), B => A(15), S => S, Z => Y(15));
   U24 : MUX2_X1 port map( A => B(14), B => A(14), S => S, Z => Y(14));
   U25 : MUX2_X1 port map( A => B(13), B => A(13), S => S, Z => Y(13));
   U26 : MUX2_X1 port map( A => B(12), B => A(12), S => S, Z => Y(12));
   U27 : MUX2_X1 port map( A => B(10), B => A(10), S => S, Z => Y(10));
   U28 : MUX2_X1 port map( A => B(8), B => A(8), S => S, Z => Y(8));
   U29 : MUX2_X1 port map( A => B(6), B => A(6), S => S, Z => Y(6));
   U30 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U31 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U32 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FD_0 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_0;

architecture SYN_ASYNCH_FD of FD_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n3, n4, n_1372 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CK, RN => n3, Q => Q_port, QN => 
                           n_1372);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n4);
   U3 : NAND2_X1 port map( A1 => RESET, A2 => ENABLE, ZN => n3);

end SYN_ASYNCH_FD;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_3 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_3;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_65
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_66
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_67
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_68
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_69
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_70
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_71
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_72
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_73
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_74
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_75
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_76
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_77
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_78
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_79
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_80
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_81
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_82
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_83
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_84
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_85
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_86
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_87
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_88
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_89
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_90
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_91
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_92
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_93
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_94
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_95
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_96
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_96 port map( D => data_in(0), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_95 port map( D => data_in(1), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_94 port map( D => data_in(2), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_93 port map( D => data_in(3), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_92 port map( D => data_in(4), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_91 port map( D => data_in(5), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_90 port map( D => data_in(6), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_89 port map( D => data_in(7), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_88 port map( D => data_in(8), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_87 port map( D => data_in(9), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_86 port map( D => data_in(10), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(10));
   FF_11 : FD_85 port map( D => data_in(11), CK => n14, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(11));
   FF_12 : FD_84 port map( D => data_in(12), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(12));
   FF_13 : FD_83 port map( D => data_in(13), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(13));
   FF_14 : FD_82 port map( D => data_in(14), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(14));
   FF_15 : FD_81 port map( D => data_in(15), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(15));
   FF_16 : FD_80 port map( D => data_in(16), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(16));
   FF_17 : FD_79 port map( D => data_in(17), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(17));
   FF_18 : FD_78 port map( D => data_in(18), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(18));
   FF_19 : FD_77 port map( D => data_in(19), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(19));
   FF_20 : FD_76 port map( D => data_in(20), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(20));
   FF_21 : FD_75 port map( D => data_in(21), CK => n14, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(21));
   FF_22 : FD_74 port map( D => data_in(22), CK => n15, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(22));
   FF_23 : FD_73 port map( D => data_in(23), CK => n15, RESET => n10, ENABLE =>
                           ENABLE, Q => data_out(23));
   FF_24 : FD_72 port map( D => data_in(24), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(24));
   FF_25 : FD_71 port map( D => data_in(25), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(25));
   FF_26 : FD_70 port map( D => data_in(26), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(26));
   FF_27 : FD_69 port map( D => data_in(27), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(27));
   FF_28 : FD_68 port map( D => data_in(28), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(28));
   FF_29 : FD_67 port map( D => data_in(29), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(29));
   FF_30 : FD_66 port map( D => data_in(30), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(30));
   FF_31 : FD_65 port map( D => data_in(31), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => CK, Z => n16);
   U3 : BUF_X1 port map( A => n12, Z => n9);
   U4 : BUF_X1 port map( A => n12, Z => n10);
   U5 : BUF_X1 port map( A => n12, Z => n11);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_4 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_4;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_97
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_98
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_99
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_100
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_101
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_102
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_103
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_104
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_105
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_106
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_107
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_108
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_109
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_110
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_111
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_112
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_113
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_114
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_115
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_116
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_117
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_118
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_119
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_120
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_121
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_122
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_123
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_124
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_125
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_126
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_127
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_128
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_128 port map( D => data_in(0), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_127 port map( D => data_in(1), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_126 port map( D => data_in(2), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_125 port map( D => data_in(3), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_124 port map( D => data_in(4), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_123 port map( D => data_in(5), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_122 port map( D => data_in(6), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_121 port map( D => data_in(7), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_120 port map( D => data_in(8), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_119 port map( D => data_in(9), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_118 port map( D => data_in(10), CK => n13, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(10));
   FF_11 : FD_117 port map( D => data_in(11), CK => n14, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(11));
   FF_12 : FD_116 port map( D => data_in(12), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(12));
   FF_13 : FD_115 port map( D => data_in(13), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(13));
   FF_14 : FD_114 port map( D => data_in(14), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(14));
   FF_15 : FD_113 port map( D => data_in(15), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(15));
   FF_16 : FD_112 port map( D => data_in(16), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(16));
   FF_17 : FD_111 port map( D => data_in(17), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(17));
   FF_18 : FD_110 port map( D => data_in(18), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(18));
   FF_19 : FD_109 port map( D => data_in(19), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(19));
   FF_20 : FD_108 port map( D => data_in(20), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(20));
   FF_21 : FD_107 port map( D => data_in(21), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(21));
   FF_22 : FD_106 port map( D => data_in(22), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(22));
   FF_23 : FD_105 port map( D => data_in(23), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(23));
   FF_24 : FD_104 port map( D => data_in(24), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(24));
   FF_25 : FD_103 port map( D => data_in(25), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(25));
   FF_26 : FD_102 port map( D => data_in(26), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(26));
   FF_27 : FD_101 port map( D => data_in(27), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(27));
   FF_28 : FD_100 port map( D => data_in(28), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(28));
   FF_29 : FD_99 port map( D => data_in(29), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(29));
   FF_30 : FD_98 port map( D => data_in(30), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(30));
   FF_31 : FD_97 port map( D => data_in(31), CK => n15, RESET => n11, ENABLE =>
                           ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => CK, Z => n16);
   U3 : BUF_X1 port map( A => n12, Z => n9);
   U4 : BUF_X1 port map( A => n12, Z => n10);
   U5 : BUF_X1 port map( A => n12, Z => n11);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_5 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_5;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_129
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_130
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_131
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_132
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_133
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_134
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_135
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_136
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_137
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_138
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_139
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_140
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_141
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_142
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_143
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_144
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_145
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_146
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_147
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_148
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_149
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_150
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_151
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_152
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_153
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_154
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_155
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_156
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_157
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_158
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_159
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_160
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_160 port map( D => data_in(0), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_159 port map( D => data_in(1), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_158 port map( D => data_in(2), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_157 port map( D => data_in(3), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_156 port map( D => data_in(4), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_155 port map( D => data_in(5), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_154 port map( D => data_in(6), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_153 port map( D => data_in(7), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_152 port map( D => data_in(8), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_151 port map( D => data_in(9), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_150 port map( D => data_in(10), CK => n13, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(10));
   FF_11 : FD_149 port map( D => data_in(11), CK => n14, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(11));
   FF_12 : FD_148 port map( D => data_in(12), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(12));
   FF_13 : FD_147 port map( D => data_in(13), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(13));
   FF_14 : FD_146 port map( D => data_in(14), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(14));
   FF_15 : FD_145 port map( D => data_in(15), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(15));
   FF_16 : FD_144 port map( D => data_in(16), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(16));
   FF_17 : FD_143 port map( D => data_in(17), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(17));
   FF_18 : FD_142 port map( D => data_in(18), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(18));
   FF_19 : FD_141 port map( D => data_in(19), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(19));
   FF_20 : FD_140 port map( D => data_in(20), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(20));
   FF_21 : FD_139 port map( D => data_in(21), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(21));
   FF_22 : FD_138 port map( D => data_in(22), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(22));
   FF_23 : FD_137 port map( D => data_in(23), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(23));
   FF_24 : FD_136 port map( D => data_in(24), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(24));
   FF_25 : FD_135 port map( D => data_in(25), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(25));
   FF_26 : FD_134 port map( D => data_in(26), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(26));
   FF_27 : FD_133 port map( D => data_in(27), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(27));
   FF_28 : FD_132 port map( D => data_in(28), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(28));
   FF_29 : FD_131 port map( D => data_in(29), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(29));
   FF_30 : FD_130 port map( D => data_in(30), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(30));
   FF_31 : FD_129 port map( D => data_in(31), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => CK, Z => n16);
   U3 : BUF_X1 port map( A => n12, Z => n9);
   U4 : BUF_X1 port map( A => n12, Z => n10);
   U5 : BUF_X1 port map( A => n12, Z => n11);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_3;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U5 : MUX2_X1 port map( A => B(4), B => A(4), S => S, Z => Y(4));
   U6 : MUX2_X1 port map( A => B(5), B => A(5), S => S, Z => Y(5));
   U7 : MUX2_X1 port map( A => B(6), B => A(6), S => S, Z => Y(6));
   U8 : MUX2_X1 port map( A => B(7), B => A(7), S => S, Z => Y(7));
   U9 : MUX2_X1 port map( A => B(8), B => A(8), S => S, Z => Y(8));
   U10 : MUX2_X1 port map( A => B(9), B => A(9), S => S, Z => Y(9));
   U11 : MUX2_X1 port map( A => B(10), B => A(10), S => S, Z => Y(10));
   U12 : MUX2_X1 port map( A => B(11), B => A(11), S => S, Z => Y(11));
   U13 : MUX2_X1 port map( A => B(12), B => A(12), S => S, Z => Y(12));
   U14 : MUX2_X1 port map( A => B(13), B => A(13), S => S, Z => Y(13));
   U15 : MUX2_X1 port map( A => B(14), B => A(14), S => S, Z => Y(14));
   U16 : MUX2_X1 port map( A => B(15), B => A(15), S => S, Z => Y(15));
   U17 : MUX2_X1 port map( A => B(16), B => A(16), S => S, Z => Y(16));
   U18 : MUX2_X1 port map( A => B(17), B => A(17), S => S, Z => Y(17));
   U19 : MUX2_X1 port map( A => B(18), B => A(18), S => S, Z => Y(18));
   U20 : MUX2_X1 port map( A => B(19), B => A(19), S => S, Z => Y(19));
   U21 : MUX2_X1 port map( A => B(20), B => A(20), S => S, Z => Y(20));
   U22 : MUX2_X1 port map( A => B(21), B => A(21), S => S, Z => Y(21));
   U23 : MUX2_X1 port map( A => B(22), B => A(22), S => S, Z => Y(22));
   U24 : MUX2_X1 port map( A => B(23), B => A(23), S => S, Z => Y(23));
   U25 : MUX2_X1 port map( A => B(24), B => A(24), S => S, Z => Y(24));
   U26 : MUX2_X1 port map( A => B(25), B => A(25), S => S, Z => Y(25));
   U27 : MUX2_X1 port map( A => B(26), B => A(26), S => S, Z => Y(26));
   U28 : MUX2_X1 port map( A => B(27), B => A(27), S => S, Z => Y(27));
   U29 : MUX2_X1 port map( A => B(28), B => A(28), S => S, Z => Y(28));
   U30 : MUX2_X1 port map( A => B(29), B => A(29), S => S, Z => Y(29));
   U31 : MUX2_X1 port map( A => B(30), B => A(30), S => S, Z => Y(30));
   U32 : MUX2_X1 port map( A => B(31), B => A(31), S => S, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_bits32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_GENERIC_bits32_0;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_bits32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => S, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => S, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => S, Z => Y(3));
   U5 : MUX2_X1 port map( A => B(4), B => A(4), S => S, Z => Y(4));
   U6 : MUX2_X1 port map( A => B(5), B => A(5), S => S, Z => Y(5));
   U7 : MUX2_X1 port map( A => B(6), B => A(6), S => S, Z => Y(6));
   U8 : MUX2_X1 port map( A => B(7), B => A(7), S => S, Z => Y(7));
   U9 : MUX2_X1 port map( A => B(8), B => A(8), S => S, Z => Y(8));
   U10 : MUX2_X1 port map( A => B(9), B => A(9), S => S, Z => Y(9));
   U11 : MUX2_X1 port map( A => B(10), B => A(10), S => S, Z => Y(10));
   U12 : MUX2_X1 port map( A => B(11), B => A(11), S => S, Z => Y(11));
   U13 : MUX2_X1 port map( A => B(12), B => A(12), S => S, Z => Y(12));
   U14 : MUX2_X1 port map( A => B(13), B => A(13), S => S, Z => Y(13));
   U15 : MUX2_X1 port map( A => B(14), B => A(14), S => S, Z => Y(14));
   U16 : MUX2_X1 port map( A => B(15), B => A(15), S => S, Z => Y(15));
   U17 : MUX2_X1 port map( A => B(16), B => A(16), S => S, Z => Y(16));
   U18 : MUX2_X1 port map( A => B(17), B => A(17), S => S, Z => Y(17));
   U19 : MUX2_X1 port map( A => B(18), B => A(18), S => S, Z => Y(18));
   U20 : MUX2_X1 port map( A => B(19), B => A(19), S => S, Z => Y(19));
   U21 : MUX2_X1 port map( A => B(20), B => A(20), S => S, Z => Y(20));
   U22 : MUX2_X1 port map( A => B(21), B => A(21), S => S, Z => Y(21));
   U23 : MUX2_X1 port map( A => B(22), B => A(22), S => S, Z => Y(22));
   U24 : MUX2_X1 port map( A => B(23), B => A(23), S => S, Z => Y(23));
   U25 : MUX2_X1 port map( A => B(24), B => A(24), S => S, Z => Y(24));
   U26 : MUX2_X1 port map( A => B(25), B => A(25), S => S, Z => Y(25));
   U27 : MUX2_X1 port map( A => B(26), B => A(26), S => S, Z => Y(26));
   U28 : MUX2_X1 port map( A => B(27), B => A(27), S => S, Z => Y(27));
   U29 : MUX2_X1 port map( A => B(28), B => A(28), S => S, Z => Y(28));
   U30 : MUX2_X1 port map( A => B(29), B => A(29), S => S, Z => Y(29));
   U31 : MUX2_X1 port map( A => B(30), B => A(30), S => S, Z => Y(30));
   U32 : MUX2_X1 port map( A => B(31), B => A(31), S => S, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_6 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_6;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_161
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_162
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_163
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_164
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_165
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_166
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_167
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_168
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_169
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_170
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_171
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_172
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_173
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_174
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_175
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_176
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_177
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_178
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_179
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_180
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_181
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_182
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_183
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_184
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_185
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_186
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_187
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_188
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_189
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_190
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_191
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_192
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_192 port map( D => data_in(0), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_191 port map( D => data_in(1), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_190 port map( D => data_in(2), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_189 port map( D => data_in(3), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_188 port map( D => data_in(4), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_187 port map( D => data_in(5), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_186 port map( D => data_in(6), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_185 port map( D => data_in(7), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_184 port map( D => data_in(8), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_183 port map( D => data_in(9), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_182 port map( D => data_in(10), CK => n13, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(10));
   FF_11 : FD_181 port map( D => data_in(11), CK => n14, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(11));
   FF_12 : FD_180 port map( D => data_in(12), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(12));
   FF_13 : FD_179 port map( D => data_in(13), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(13));
   FF_14 : FD_178 port map( D => data_in(14), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(14));
   FF_15 : FD_177 port map( D => data_in(15), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(15));
   FF_16 : FD_176 port map( D => data_in(16), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(16));
   FF_17 : FD_175 port map( D => data_in(17), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(17));
   FF_18 : FD_174 port map( D => data_in(18), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(18));
   FF_19 : FD_173 port map( D => data_in(19), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(19));
   FF_20 : FD_172 port map( D => data_in(20), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(20));
   FF_21 : FD_171 port map( D => data_in(21), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(21));
   FF_22 : FD_170 port map( D => data_in(22), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(22));
   FF_23 : FD_169 port map( D => data_in(23), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(23));
   FF_24 : FD_168 port map( D => data_in(24), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(24));
   FF_25 : FD_167 port map( D => data_in(25), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(25));
   FF_26 : FD_166 port map( D => data_in(26), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(26));
   FF_27 : FD_165 port map( D => data_in(27), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(27));
   FF_28 : FD_164 port map( D => data_in(28), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(28));
   FF_29 : FD_163 port map( D => data_in(29), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(29));
   FF_30 : FD_162 port map( D => data_in(30), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(30));
   FF_31 : FD_161 port map( D => data_in(31), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => CK, Z => n16);
   U2 : BUF_X1 port map( A => RESET, Z => n12);
   U3 : BUF_X1 port map( A => n12, Z => n9);
   U4 : BUF_X1 port map( A => n12, Z => n10);
   U5 : BUF_X1 port map( A => n12, Z => n11);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_7 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_7;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_7 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_193
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_194
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_195
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_196
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_197
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_198
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_199
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_200
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_201
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_202
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_203
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_204
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_205
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_206
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_207
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_208
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_209
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_210
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_211
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_212
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_213
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_214
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_215
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_216
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_217
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_218
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_219
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_220
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_221
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_222
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_223
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_224
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_224 port map( D => data_in(0), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_223 port map( D => data_in(1), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_222 port map( D => data_in(2), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_221 port map( D => data_in(3), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_220 port map( D => data_in(4), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_219 port map( D => data_in(5), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_218 port map( D => data_in(6), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_217 port map( D => data_in(7), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_216 port map( D => data_in(8), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_215 port map( D => data_in(9), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_214 port map( D => data_in(10), CK => n13, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(10));
   FF_11 : FD_213 port map( D => data_in(11), CK => n14, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(11));
   FF_12 : FD_212 port map( D => data_in(12), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(12));
   FF_13 : FD_211 port map( D => data_in(13), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(13));
   FF_14 : FD_210 port map( D => data_in(14), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(14));
   FF_15 : FD_209 port map( D => data_in(15), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(15));
   FF_16 : FD_208 port map( D => data_in(16), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(16));
   FF_17 : FD_207 port map( D => data_in(17), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(17));
   FF_18 : FD_206 port map( D => data_in(18), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(18));
   FF_19 : FD_205 port map( D => data_in(19), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(19));
   FF_20 : FD_204 port map( D => data_in(20), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(20));
   FF_21 : FD_203 port map( D => data_in(21), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(21));
   FF_22 : FD_202 port map( D => data_in(22), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(22));
   FF_23 : FD_201 port map( D => data_in(23), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(23));
   FF_24 : FD_200 port map( D => data_in(24), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(24));
   FF_25 : FD_199 port map( D => data_in(25), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(25));
   FF_26 : FD_198 port map( D => data_in(26), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(26));
   FF_27 : FD_197 port map( D => data_in(27), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(27));
   FF_28 : FD_196 port map( D => data_in(28), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(28));
   FF_29 : FD_195 port map( D => data_in(29), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(29));
   FF_30 : FD_194 port map( D => data_in(30), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(30));
   FF_31 : FD_193 port map( D => data_in(31), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => CK, Z => n16);
   U2 : BUF_X1 port map( A => RESET, Z => n12);
   U3 : BUF_X1 port map( A => n12, Z => n9);
   U4 : BUF_X1 port map( A => n12, Z => n10);
   U5 : BUF_X1 port map( A => n12, Z => n11);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_8 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_8;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_8 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_225
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_226
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_227
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_228
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_229
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_230
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_231
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_232
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_233
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_234
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_235
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_236
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_237
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_238
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_239
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_240
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_241
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_242
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_243
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_244
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_245
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_246
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_247
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_248
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_249
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_250
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_251
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_252
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_253
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_254
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_255
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_256
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_256 port map( D => data_in(0), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_255 port map( D => data_in(1), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_254 port map( D => data_in(2), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_253 port map( D => data_in(3), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_252 port map( D => data_in(4), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_251 port map( D => data_in(5), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_250 port map( D => data_in(6), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_249 port map( D => data_in(7), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_248 port map( D => data_in(8), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_247 port map( D => data_in(9), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_246 port map( D => data_in(10), CK => n13, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(10));
   FF_11 : FD_245 port map( D => data_in(11), CK => n14, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(11));
   FF_12 : FD_244 port map( D => data_in(12), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(12));
   FF_13 : FD_243 port map( D => data_in(13), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(13));
   FF_14 : FD_242 port map( D => data_in(14), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(14));
   FF_15 : FD_241 port map( D => data_in(15), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(15));
   FF_16 : FD_240 port map( D => data_in(16), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(16));
   FF_17 : FD_239 port map( D => data_in(17), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(17));
   FF_18 : FD_238 port map( D => data_in(18), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(18));
   FF_19 : FD_237 port map( D => data_in(19), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(19));
   FF_20 : FD_236 port map( D => data_in(20), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(20));
   FF_21 : FD_235 port map( D => data_in(21), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(21));
   FF_22 : FD_234 port map( D => data_in(22), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(22));
   FF_23 : FD_233 port map( D => data_in(23), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(23));
   FF_24 : FD_232 port map( D => data_in(24), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(24));
   FF_25 : FD_231 port map( D => data_in(25), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(25));
   FF_26 : FD_230 port map( D => data_in(26), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(26));
   FF_27 : FD_229 port map( D => data_in(27), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(27));
   FF_28 : FD_228 port map( D => data_in(28), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(28));
   FF_29 : FD_227 port map( D => data_in(29), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(29));
   FF_30 : FD_226 port map( D => data_in(30), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(30));
   FF_31 : FD_225 port map( D => data_in(31), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => CK, Z => n16);
   U2 : BUF_X1 port map( A => RESET, Z => n12);
   U3 : BUF_X1 port map( A => n12, Z => n9);
   U4 : BUF_X1 port map( A => n12, Z => n10);
   U5 : BUF_X1 port map( A => n12, Z => n11);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_9 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_9;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_9 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_257
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_258
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_259
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_260
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_261
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_262
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_263
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_264
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_265
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_266
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_267
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_268
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_269
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_270
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_271
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_272
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_273
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_274
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_275
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_276
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_277
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_278
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_279
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_280
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_281
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_282
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_283
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_284
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_285
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_286
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_287
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_288
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_288 port map( D => data_in(0), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_287 port map( D => data_in(1), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_286 port map( D => data_in(2), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_285 port map( D => data_in(3), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_284 port map( D => data_in(4), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_283 port map( D => data_in(5), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_282 port map( D => data_in(6), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_281 port map( D => data_in(7), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_280 port map( D => data_in(8), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_279 port map( D => data_in(9), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_278 port map( D => data_in(10), CK => n13, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(10));
   FF_11 : FD_277 port map( D => data_in(11), CK => n14, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(11));
   FF_12 : FD_276 port map( D => data_in(12), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(12));
   FF_13 : FD_275 port map( D => data_in(13), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(13));
   FF_14 : FD_274 port map( D => data_in(14), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(14));
   FF_15 : FD_273 port map( D => data_in(15), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(15));
   FF_16 : FD_272 port map( D => data_in(16), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(16));
   FF_17 : FD_271 port map( D => data_in(17), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(17));
   FF_18 : FD_270 port map( D => data_in(18), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(18));
   FF_19 : FD_269 port map( D => data_in(19), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(19));
   FF_20 : FD_268 port map( D => data_in(20), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(20));
   FF_21 : FD_267 port map( D => data_in(21), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(21));
   FF_22 : FD_266 port map( D => data_in(22), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(22));
   FF_23 : FD_265 port map( D => data_in(23), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(23));
   FF_24 : FD_264 port map( D => data_in(24), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(24));
   FF_25 : FD_263 port map( D => data_in(25), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(25));
   FF_26 : FD_262 port map( D => data_in(26), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(26));
   FF_27 : FD_261 port map( D => data_in(27), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(27));
   FF_28 : FD_260 port map( D => data_in(28), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(28));
   FF_29 : FD_259 port map( D => data_in(29), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(29));
   FF_30 : FD_258 port map( D => data_in(30), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(30));
   FF_31 : FD_257 port map( D => data_in(31), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => CK, Z => n16);
   U3 : BUF_X1 port map( A => n12, Z => n9);
   U4 : BUF_X1 port map( A => n12, Z => n10);
   U5 : BUF_X1 port map( A => n12, Z => n11);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_10 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_10;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_10 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_289
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_290
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_291
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_292
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_293
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_294
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_295
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_296
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_297
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_298
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_299
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_300
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_301
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_302
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_303
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_304
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_305
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_306
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_307
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_308
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_309
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_310
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_311
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_312
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_313
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_314
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_315
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_316
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_317
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_318
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_319
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_320
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_320 port map( D => data_in(0), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_319 port map( D => data_in(1), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_318 port map( D => data_in(2), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_317 port map( D => data_in(3), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_316 port map( D => data_in(4), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_315 port map( D => data_in(5), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_314 port map( D => data_in(6), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_313 port map( D => data_in(7), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_312 port map( D => data_in(8), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_311 port map( D => data_in(9), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_310 port map( D => data_in(10), CK => n13, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(10));
   FF_11 : FD_309 port map( D => data_in(11), CK => n14, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(11));
   FF_12 : FD_308 port map( D => data_in(12), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(12));
   FF_13 : FD_307 port map( D => data_in(13), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(13));
   FF_14 : FD_306 port map( D => data_in(14), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(14));
   FF_15 : FD_305 port map( D => data_in(15), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(15));
   FF_16 : FD_304 port map( D => data_in(16), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(16));
   FF_17 : FD_303 port map( D => data_in(17), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(17));
   FF_18 : FD_302 port map( D => data_in(18), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(18));
   FF_19 : FD_301 port map( D => data_in(19), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(19));
   FF_20 : FD_300 port map( D => data_in(20), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(20));
   FF_21 : FD_299 port map( D => data_in(21), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(21));
   FF_22 : FD_298 port map( D => data_in(22), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(22));
   FF_23 : FD_297 port map( D => data_in(23), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(23));
   FF_24 : FD_296 port map( D => data_in(24), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(24));
   FF_25 : FD_295 port map( D => data_in(25), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(25));
   FF_26 : FD_294 port map( D => data_in(26), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(26));
   FF_27 : FD_293 port map( D => data_in(27), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(27));
   FF_28 : FD_292 port map( D => data_in(28), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(28));
   FF_29 : FD_291 port map( D => data_in(29), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(29));
   FF_30 : FD_290 port map( D => data_in(30), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(30));
   FF_31 : FD_289 port map( D => data_in(31), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => CK, Z => n16);
   U3 : BUF_X1 port map( A => n12, Z => n9);
   U4 : BUF_X1 port map( A => n12, Z => n10);
   U5 : BUF_X1 port map( A => n12, Z => n11);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity register_generic_nbits32_0 is

   port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  data_out : out std_logic_vector (31 downto 0));

end register_generic_nbits32_0;

architecture SYN_ASYNCHRONOUS of register_generic_nbits32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_321
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_322
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_323
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_324
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_325
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_326
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_327
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_328
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_329
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_330
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_331
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_332
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_333
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_334
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_335
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_336
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_337
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_338
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_339
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_340
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_341
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_342
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_343
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_344
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_345
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_346
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_347
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_348
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_349
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_350
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_351
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_352
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16 : std_logic;

begin
   
   FF_0 : FD_352 port map( D => data_in(0), CK => n15, RESET => n11, ENABLE => 
                           ENABLE, Q => data_out(0));
   FF_1 : FD_351 port map( D => data_in(1), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(1));
   FF_2 : FD_350 port map( D => data_in(2), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(2));
   FF_3 : FD_349 port map( D => data_in(3), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(3));
   FF_4 : FD_348 port map( D => data_in(4), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(4));
   FF_5 : FD_347 port map( D => data_in(5), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(5));
   FF_6 : FD_346 port map( D => data_in(6), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(6));
   FF_7 : FD_345 port map( D => data_in(7), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(7));
   FF_8 : FD_344 port map( D => data_in(8), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(8));
   FF_9 : FD_343 port map( D => data_in(9), CK => n13, RESET => n9, ENABLE => 
                           ENABLE, Q => data_out(9));
   FF_10 : FD_342 port map( D => data_in(10), CK => n13, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(10));
   FF_11 : FD_341 port map( D => data_in(11), CK => n13, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(11));
   FF_12 : FD_340 port map( D => data_in(12), CK => n14, RESET => n9, ENABLE =>
                           ENABLE, Q => data_out(12));
   FF_13 : FD_339 port map( D => data_in(13), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(13));
   FF_14 : FD_338 port map( D => data_in(14), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(14));
   FF_15 : FD_337 port map( D => data_in(15), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(15));
   FF_16 : FD_336 port map( D => data_in(16), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(16));
   FF_17 : FD_335 port map( D => data_in(17), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(17));
   FF_18 : FD_334 port map( D => data_in(18), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(18));
   FF_19 : FD_333 port map( D => data_in(19), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(19));
   FF_20 : FD_332 port map( D => data_in(20), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(20));
   FF_21 : FD_331 port map( D => data_in(21), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(21));
   FF_22 : FD_330 port map( D => data_in(22), CK => n14, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(22));
   FF_23 : FD_329 port map( D => data_in(23), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(23));
   FF_24 : FD_328 port map( D => data_in(24), CK => n15, RESET => n10, ENABLE 
                           => ENABLE, Q => data_out(24));
   FF_25 : FD_327 port map( D => data_in(25), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(25));
   FF_26 : FD_326 port map( D => data_in(26), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(26));
   FF_27 : FD_325 port map( D => data_in(27), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(27));
   FF_28 : FD_324 port map( D => data_in(28), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(28));
   FF_29 : FD_323 port map( D => data_in(29), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(29));
   FF_30 : FD_322 port map( D => data_in(30), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(30));
   FF_31 : FD_321 port map( D => data_in(31), CK => n15, RESET => n11, ENABLE 
                           => ENABLE, Q => data_out(31));
   U1 : BUF_X1 port map( A => RESET, Z => n12);
   U2 : BUF_X1 port map( A => CK, Z => n16);
   U3 : BUF_X1 port map( A => n12, Z => n9);
   U4 : BUF_X1 port map( A => n12, Z => n10);
   U5 : BUF_X1 port map( A => n12, Z => n11);
   U6 : BUF_X1 port map( A => n16, Z => n13);
   U7 : BUF_X1 port map( A => n16, Z => n14);
   U8 : BUF_X1 port map( A => n16, Z => n15);

end SYN_ASYNCHRONOUS;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4 is

   port( A, B : in std_logic_vector (32 downto 1);  C0 : in std_logic;  COUT : 
         out std_logic_vector (8 downto 0));

end CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4;

architecture SYN_STRUCTURAL of CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_1
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_2
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_3
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_4
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_1
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_2
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_5
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component G_6
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_3
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_4
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_5
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_7
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_6
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_7
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_8
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_9
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_10
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_11
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_12
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_8
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component PG_13
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_14
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_15
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_16
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_17
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_18
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_19
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_20
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_21
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_22
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_23
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_24
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_25
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_26
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component PG_0
      port( p_ik, g_ik, p_k1j, g_k1j : in std_logic;  P_ij, G_ij : out 
            std_logic);
   end component;
   
   component G_0
      port( p_ik, g_ik, g_k1j : in std_logic;  G_ij : out std_logic);
   end component;
   
   component pg_generator_1
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_2
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_3
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_4
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_5
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_6
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_7
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_8
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_9
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_10
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_11
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_12
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_13
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_14
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_15
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_16
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_17
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_18
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_19
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_20
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_21
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_22
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_23
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_24
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_25
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_26
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_27
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_28
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_29
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_30
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_31
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component pg_generator_0
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   signal COUT_8_port, COUT_7_port, COUT_6_port, COUT_5_port, COUT_4_port, 
      COUT_3_port, COUT_2_port, COUT_1_port, gi_1_port, pi_1_port, 
      gSignal_16_16_port, gSignal_16_15_port, gSignal_16_13_port, 
      gSignal_16_9_port, gSignal_15_15_port, gSignal_14_14_port, 
      gSignal_14_13_port, gSignal_13_13_port, gSignal_12_12_port, 
      gSignal_12_11_port, gSignal_12_9_port, gSignal_11_11_port, 
      gSignal_10_10_port, gSignal_10_9_port, gSignal_9_9_port, gSignal_8_8_port
      , gSignal_8_7_port, gSignal_8_5_port, gSignal_7_7_port, gSignal_6_6_port,
      gSignal_6_5_port, gSignal_5_5_port, gSignal_4_4_port, gSignal_4_3_port, 
      gSignal_3_3_port, gSignal_2_2_port, gSignal_2_1_port, pSignal_16_16_port,
      pSignal_16_15_port, pSignal_16_13_port, pSignal_16_9_port, 
      pSignal_15_15_port, pSignal_14_14_port, pSignal_14_13_port, 
      pSignal_13_13_port, pSignal_12_12_port, pSignal_12_11_port, 
      pSignal_12_9_port, pSignal_11_11_port, pSignal_10_10_port, 
      pSignal_10_9_port, pSignal_9_9_port, pSignal_8_8_port, pSignal_8_7_port, 
      pSignal_8_5_port, pSignal_7_7_port, pSignal_6_6_port, pSignal_6_5_port, 
      pSignal_5_5_port, pSignal_4_4_port, pSignal_4_3_port, pSignal_3_3_port, 
      pSignal_2_2_port, pSignal_32_32_port, pSignal_32_31_port, 
      pSignal_32_29_port, pSignal_32_25_port, pSignal_32_17_port, 
      pSignal_31_31_port, pSignal_30_30_port, pSignal_30_29_port, 
      pSignal_29_29_port, pSignal_28_28_port, pSignal_28_27_port, 
      pSignal_28_25_port, pSignal_28_17_port, pSignal_27_27_port, 
      pSignal_26_26_port, pSignal_26_25_port, pSignal_25_25_port, 
      pSignal_24_24_port, pSignal_24_23_port, pSignal_24_21_port, 
      pSignal_24_17_port, pSignal_23_23_port, pSignal_22_22_port, 
      pSignal_22_21_port, pSignal_21_21_port, pSignal_20_20_port, 
      pSignal_20_19_port, pSignal_20_17_port, pSignal_19_19_port, 
      pSignal_18_18_port, pSignal_18_17_port, pSignal_17_17_port, 
      gSignal_32_32_port, gSignal_32_31_port, gSignal_32_29_port, 
      gSignal_32_25_port, gSignal_32_17_port, gSignal_31_31_port, 
      gSignal_30_30_port, gSignal_30_29_port, gSignal_29_29_port, 
      gSignal_28_28_port, gSignal_28_27_port, gSignal_28_25_port, 
      gSignal_28_17_port, gSignal_27_27_port, gSignal_26_26_port, 
      gSignal_26_25_port, gSignal_25_25_port, gSignal_24_24_port, 
      gSignal_24_23_port, gSignal_24_21_port, gSignal_24_17_port, 
      gSignal_23_23_port, gSignal_22_22_port, gSignal_22_21_port, 
      gSignal_21_21_port, gSignal_20_20_port, gSignal_20_19_port, 
      gSignal_20_17_port, gSignal_19_19_port, gSignal_18_18_port, 
      gSignal_18_17_port, gSignal_17_17_port, n3, n4 : std_logic;

begin
   COUT <= ( COUT_8_port, COUT_7_port, COUT_6_port, COUT_5_port, COUT_4_port, 
      COUT_3_port, COUT_2_port, COUT_1_port, C0 );
   
   pg_inst_1 : pg_generator_0 port map( A => A(1), B => B(1), P => pi_1_port, G
                           => gi_1_port);
   pg_inst_2 : pg_generator_31 port map( A => A(2), B => B(2), P => 
                           pSignal_2_2_port, G => gSignal_2_2_port);
   pg_inst_3 : pg_generator_30 port map( A => A(3), B => B(3), P => 
                           pSignal_3_3_port, G => gSignal_3_3_port);
   pg_inst_4 : pg_generator_29 port map( A => A(4), B => B(4), P => 
                           pSignal_4_4_port, G => gSignal_4_4_port);
   pg_inst_5 : pg_generator_28 port map( A => A(5), B => B(5), P => 
                           pSignal_5_5_port, G => gSignal_5_5_port);
   pg_inst_6 : pg_generator_27 port map( A => A(6), B => B(6), P => 
                           pSignal_6_6_port, G => gSignal_6_6_port);
   pg_inst_7 : pg_generator_26 port map( A => A(7), B => B(7), P => 
                           pSignal_7_7_port, G => gSignal_7_7_port);
   pg_inst_8 : pg_generator_25 port map( A => A(8), B => B(8), P => 
                           pSignal_8_8_port, G => gSignal_8_8_port);
   pg_inst_9 : pg_generator_24 port map( A => A(9), B => B(9), P => 
                           pSignal_9_9_port, G => gSignal_9_9_port);
   pg_inst_10 : pg_generator_23 port map( A => A(10), B => B(10), P => 
                           pSignal_10_10_port, G => gSignal_10_10_port);
   pg_inst_11 : pg_generator_22 port map( A => A(11), B => B(11), P => 
                           pSignal_11_11_port, G => gSignal_11_11_port);
   pg_inst_12 : pg_generator_21 port map( A => A(12), B => B(12), P => 
                           pSignal_12_12_port, G => gSignal_12_12_port);
   pg_inst_13 : pg_generator_20 port map( A => A(13), B => B(13), P => 
                           pSignal_13_13_port, G => gSignal_13_13_port);
   pg_inst_14 : pg_generator_19 port map( A => A(14), B => B(14), P => 
                           pSignal_14_14_port, G => gSignal_14_14_port);
   pg_inst_15 : pg_generator_18 port map( A => A(15), B => B(15), P => 
                           pSignal_15_15_port, G => gSignal_15_15_port);
   pg_inst_16 : pg_generator_17 port map( A => A(16), B => B(16), P => 
                           pSignal_16_16_port, G => gSignal_16_16_port);
   pg_inst_17 : pg_generator_16 port map( A => A(17), B => B(17), P => 
                           pSignal_17_17_port, G => gSignal_17_17_port);
   pg_inst_18 : pg_generator_15 port map( A => A(18), B => B(18), P => 
                           pSignal_18_18_port, G => gSignal_18_18_port);
   pg_inst_19 : pg_generator_14 port map( A => A(19), B => B(19), P => 
                           pSignal_19_19_port, G => gSignal_19_19_port);
   pg_inst_20 : pg_generator_13 port map( A => A(20), B => B(20), P => 
                           pSignal_20_20_port, G => gSignal_20_20_port);
   pg_inst_21 : pg_generator_12 port map( A => A(21), B => B(21), P => 
                           pSignal_21_21_port, G => gSignal_21_21_port);
   pg_inst_22 : pg_generator_11 port map( A => A(22), B => B(22), P => 
                           pSignal_22_22_port, G => gSignal_22_22_port);
   pg_inst_23 : pg_generator_10 port map( A => A(23), B => B(23), P => 
                           pSignal_23_23_port, G => gSignal_23_23_port);
   pg_inst_24 : pg_generator_9 port map( A => A(24), B => B(24), P => 
                           pSignal_24_24_port, G => gSignal_24_24_port);
   pg_inst_25 : pg_generator_8 port map( A => A(25), B => B(25), P => 
                           pSignal_25_25_port, G => gSignal_25_25_port);
   pg_inst_26 : pg_generator_7 port map( A => A(26), B => B(26), P => 
                           pSignal_26_26_port, G => gSignal_26_26_port);
   pg_inst_27 : pg_generator_6 port map( A => A(27), B => B(27), P => 
                           pSignal_27_27_port, G => gSignal_27_27_port);
   pg_inst_28 : pg_generator_5 port map( A => A(28), B => B(28), P => 
                           pSignal_28_28_port, G => gSignal_28_28_port);
   pg_inst_29 : pg_generator_4 port map( A => A(29), B => B(29), P => 
                           pSignal_29_29_port, G => gSignal_29_29_port);
   pg_inst_30 : pg_generator_3 port map( A => A(30), B => B(30), P => 
                           pSignal_30_30_port, G => gSignal_30_30_port);
   pg_inst_31 : pg_generator_2 port map( A => A(31), B => B(31), P => 
                           pSignal_31_31_port, G => gSignal_31_31_port);
   pg_inst_32 : pg_generator_1 port map( A => A(32), B => B(32), P => 
                           pSignal_32_32_port, G => gSignal_32_32_port);
   G1_1_2 : G_0 port map( p_ik => pSignal_2_2_port, g_ik => gSignal_2_2_port, 
                           g_k1j => n4, G_ij => gSignal_2_1_port);
   PG_inst1_1_4 : PG_0 port map( p_ik => pSignal_4_4_port, g_ik => 
                           gSignal_4_4_port, p_k1j => pSignal_3_3_port, g_k1j 
                           => gSignal_3_3_port, P_ij => pSignal_4_3_port, G_ij 
                           => gSignal_4_3_port);
   PG_inst1_1_6 : PG_26 port map( p_ik => pSignal_6_6_port, g_ik => 
                           gSignal_6_6_port, p_k1j => pSignal_5_5_port, g_k1j 
                           => gSignal_5_5_port, P_ij => pSignal_6_5_port, G_ij 
                           => gSignal_6_5_port);
   PG_inst1_1_8 : PG_25 port map( p_ik => pSignal_8_8_port, g_ik => 
                           gSignal_8_8_port, p_k1j => pSignal_7_7_port, g_k1j 
                           => gSignal_7_7_port, P_ij => pSignal_8_7_port, G_ij 
                           => gSignal_8_7_port);
   PG_inst1_1_10 : PG_24 port map( p_ik => pSignal_10_10_port, g_ik => 
                           gSignal_10_10_port, p_k1j => pSignal_9_9_port, g_k1j
                           => gSignal_9_9_port, P_ij => pSignal_10_9_port, G_ij
                           => gSignal_10_9_port);
   PG_inst1_1_12 : PG_23 port map( p_ik => pSignal_12_12_port, g_ik => 
                           gSignal_12_12_port, p_k1j => pSignal_11_11_port, 
                           g_k1j => gSignal_11_11_port, P_ij => 
                           pSignal_12_11_port, G_ij => gSignal_12_11_port);
   PG_inst1_1_14 : PG_22 port map( p_ik => pSignal_14_14_port, g_ik => 
                           gSignal_14_14_port, p_k1j => pSignal_13_13_port, 
                           g_k1j => gSignal_13_13_port, P_ij => 
                           pSignal_14_13_port, G_ij => gSignal_14_13_port);
   PG_inst1_1_16 : PG_21 port map( p_ik => pSignal_16_16_port, g_ik => 
                           gSignal_16_16_port, p_k1j => pSignal_15_15_port, 
                           g_k1j => gSignal_15_15_port, P_ij => 
                           pSignal_16_15_port, G_ij => gSignal_16_15_port);
   PG_inst1_1_18 : PG_20 port map( p_ik => pSignal_18_18_port, g_ik => 
                           gSignal_18_18_port, p_k1j => pSignal_17_17_port, 
                           g_k1j => gSignal_17_17_port, P_ij => 
                           pSignal_18_17_port, G_ij => gSignal_18_17_port);
   PG_inst1_1_20 : PG_19 port map( p_ik => pSignal_20_20_port, g_ik => 
                           gSignal_20_20_port, p_k1j => pSignal_19_19_port, 
                           g_k1j => gSignal_19_19_port, P_ij => 
                           pSignal_20_19_port, G_ij => gSignal_20_19_port);
   PG_inst1_1_22 : PG_18 port map( p_ik => pSignal_22_22_port, g_ik => 
                           gSignal_22_22_port, p_k1j => pSignal_21_21_port, 
                           g_k1j => gSignal_21_21_port, P_ij => 
                           pSignal_22_21_port, G_ij => gSignal_22_21_port);
   PG_inst1_1_24 : PG_17 port map( p_ik => pSignal_24_24_port, g_ik => 
                           gSignal_24_24_port, p_k1j => pSignal_23_23_port, 
                           g_k1j => gSignal_23_23_port, P_ij => 
                           pSignal_24_23_port, G_ij => gSignal_24_23_port);
   PG_inst1_1_26 : PG_16 port map( p_ik => pSignal_26_26_port, g_ik => 
                           gSignal_26_26_port, p_k1j => pSignal_25_25_port, 
                           g_k1j => gSignal_25_25_port, P_ij => 
                           pSignal_26_25_port, G_ij => gSignal_26_25_port);
   PG_inst1_1_28 : PG_15 port map( p_ik => pSignal_28_28_port, g_ik => 
                           gSignal_28_28_port, p_k1j => pSignal_27_27_port, 
                           g_k1j => gSignal_27_27_port, P_ij => 
                           pSignal_28_27_port, G_ij => gSignal_28_27_port);
   PG_inst1_1_30 : PG_14 port map( p_ik => pSignal_30_30_port, g_ik => 
                           gSignal_30_30_port, p_k1j => pSignal_29_29_port, 
                           g_k1j => gSignal_29_29_port, P_ij => 
                           pSignal_30_29_port, G_ij => gSignal_30_29_port);
   PG_inst1_1_32 : PG_13 port map( p_ik => pSignal_32_32_port, g_ik => 
                           gSignal_32_32_port, p_k1j => pSignal_31_31_port, 
                           g_k1j => gSignal_31_31_port, P_ij => 
                           pSignal_32_31_port, G_ij => gSignal_32_31_port);
   G1_2_4 : G_8 port map( p_ik => pSignal_4_3_port, g_ik => gSignal_4_3_port, 
                           g_k1j => gSignal_2_1_port, G_ij => COUT_1_port);
   PG_inst1_2_8 : PG_12 port map( p_ik => pSignal_8_7_port, g_ik => 
                           gSignal_8_7_port, p_k1j => pSignal_6_5_port, g_k1j 
                           => gSignal_6_5_port, P_ij => pSignal_8_5_port, G_ij 
                           => gSignal_8_5_port);
   PG_inst1_2_12 : PG_11 port map( p_ik => pSignal_12_11_port, g_ik => 
                           gSignal_12_11_port, p_k1j => pSignal_10_9_port, 
                           g_k1j => gSignal_10_9_port, P_ij => 
                           pSignal_12_9_port, G_ij => gSignal_12_9_port);
   PG_inst1_2_16 : PG_10 port map( p_ik => pSignal_16_15_port, g_ik => 
                           gSignal_16_15_port, p_k1j => pSignal_14_13_port, 
                           g_k1j => gSignal_14_13_port, P_ij => 
                           pSignal_16_13_port, G_ij => gSignal_16_13_port);
   PG_inst1_2_20 : PG_9 port map( p_ik => pSignal_20_19_port, g_ik => 
                           gSignal_20_19_port, p_k1j => pSignal_18_17_port, 
                           g_k1j => gSignal_18_17_port, P_ij => 
                           pSignal_20_17_port, G_ij => gSignal_20_17_port);
   PG_inst1_2_24 : PG_8 port map( p_ik => pSignal_24_23_port, g_ik => 
                           gSignal_24_23_port, p_k1j => pSignal_22_21_port, 
                           g_k1j => gSignal_22_21_port, P_ij => 
                           pSignal_24_21_port, G_ij => gSignal_24_21_port);
   PG_inst1_2_28 : PG_7 port map( p_ik => pSignal_28_27_port, g_ik => 
                           gSignal_28_27_port, p_k1j => pSignal_26_25_port, 
                           g_k1j => gSignal_26_25_port, P_ij => 
                           pSignal_28_25_port, G_ij => gSignal_28_25_port);
   PG_inst1_2_32 : PG_6 port map( p_ik => pSignal_32_31_port, g_ik => 
                           gSignal_32_31_port, p_k1j => pSignal_30_29_port, 
                           g_k1j => gSignal_30_29_port, P_ij => 
                           pSignal_32_29_port, G_ij => gSignal_32_29_port);
   G_INST2_0_4_8 : G_7 port map( p_ik => pSignal_8_5_port, g_ik => 
                           gSignal_8_5_port, g_k1j => COUT_1_port, G_ij => 
                           COUT_2_port);
   PG_INST2_0_12_16 : PG_5 port map( p_ik => pSignal_16_13_port, g_ik => 
                           gSignal_16_13_port, p_k1j => pSignal_12_9_port, 
                           g_k1j => gSignal_12_9_port, P_ij => 
                           pSignal_16_9_port, G_ij => gSignal_16_9_port);
   PG_INST2_0_20_24 : PG_4 port map( p_ik => pSignal_24_21_port, g_ik => 
                           gSignal_24_21_port, p_k1j => pSignal_20_17_port, 
                           g_k1j => gSignal_20_17_port, P_ij => 
                           pSignal_24_17_port, G_ij => gSignal_24_17_port);
   PG_INST2_0_28_32 : PG_3 port map( p_ik => pSignal_32_29_port, g_ik => 
                           gSignal_32_29_port, p_k1j => pSignal_28_25_port, 
                           g_k1j => gSignal_28_25_port, P_ij => 
                           pSignal_32_25_port, G_ij => gSignal_32_25_port);
   G_INST2_1_8_12 : G_6 port map( p_ik => pSignal_12_9_port, g_ik => 
                           gSignal_12_9_port, g_k1j => COUT_2_port, G_ij => 
                           COUT_3_port);
   G_INST2_1_8_16 : G_5 port map( p_ik => pSignal_16_9_port, g_ik => 
                           gSignal_16_9_port, g_k1j => COUT_2_port, G_ij => 
                           COUT_4_port);
   PG_INST2_1_24_28 : PG_2 port map( p_ik => pSignal_28_25_port, g_ik => 
                           gSignal_28_25_port, p_k1j => pSignal_24_17_port, 
                           g_k1j => gSignal_24_17_port, P_ij => 
                           pSignal_28_17_port, G_ij => gSignal_28_17_port);
   PG_INST2_1_24_32 : PG_1 port map( p_ik => pSignal_32_25_port, g_ik => 
                           gSignal_32_25_port, p_k1j => pSignal_24_17_port, 
                           g_k1j => gSignal_24_17_port, P_ij => 
                           pSignal_32_17_port, G_ij => gSignal_32_17_port);
   G_INST2_2_16_20 : G_4 port map( p_ik => pSignal_20_17_port, g_ik => 
                           gSignal_20_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_5_port);
   G_INST2_2_16_24 : G_3 port map( p_ik => pSignal_24_17_port, g_ik => 
                           gSignal_24_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_6_port);
   G_INST2_2_16_28 : G_2 port map( p_ik => pSignal_28_17_port, g_ik => 
                           gSignal_28_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_7_port);
   G_INST2_2_16_32 : G_1 port map( p_ik => pSignal_32_17_port, g_ik => 
                           gSignal_32_17_port, g_k1j => COUT_4_port, G_ij => 
                           COUT_8_port);
   U1 : INV_X1 port map( A => n3, ZN => n4);
   U2 : AOI21_X1 port map( B1 => pi_1_port, B2 => C0, A => gi_1_port, ZN => n3)
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (8
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8;

architecture SYN_STRUCTURAL of 
   SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8 is

   component CarrySelect_1
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_2
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_3
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_4
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_5
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_6
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_7
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CarrySelect_0
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   carrySel_0 : CarrySelect_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Cin => Ci(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   carrySel_1 : CarrySelect_7 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Cin => Ci(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   carrySel_2 : CarrySelect_6 port map( A(3) => A(11), A(2) => A(10), A(1) => 
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Cin => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   carrySel_3 : CarrySelect_5 port map( A(3) => A(15), A(2) => A(14), A(1) => 
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Cin => Ci(3), S(3) => 
                           S(15), S(2) => S(14), S(1) => S(13), S(0) => S(12));
   carrySel_4 : CarrySelect_4 port map( A(3) => A(19), A(2) => A(18), A(1) => 
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Cin => Ci(4), S(3) => 
                           S(19), S(2) => S(18), S(1) => S(17), S(0) => S(16));
   carrySel_5 : CarrySelect_3 port map( A(3) => A(23), A(2) => A(22), A(1) => 
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Cin => Ci(5), S(3) => 
                           S(23), S(2) => S(22), S(1) => S(21), S(0) => S(20));
   carrySel_6 : CarrySelect_2 port map( A(3) => A(27), A(2) => A(26), A(1) => 
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Cin => Ci(6), S(3) => 
                           S(27), S(2) => S(26), S(1) => S(25), S(0) => S(24));
   carrySel_7 : CarrySelect_1 port map( A(3) => A(31), A(2) => A(30), A(1) => 
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Cin => Ci(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_logic_nbits32 is

   port( Cin : in std_logic;  B0 : in std_logic_vector (31 downto 0);  B : out 
         std_logic_vector (31 downto 0));

end xor_logic_nbits32;

architecture SYN_BEHAVIORAL of xor_logic_nbits32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => Cin, B => B0(9), Z => B(9));
   U2 : XOR2_X1 port map( A => Cin, B => B0(8), Z => B(8));
   U3 : XOR2_X1 port map( A => Cin, B => B0(7), Z => B(7));
   U4 : XOR2_X1 port map( A => Cin, B => B0(6), Z => B(6));
   U5 : XOR2_X1 port map( A => Cin, B => B0(5), Z => B(5));
   U6 : XOR2_X1 port map( A => Cin, B => B0(4), Z => B(4));
   U7 : XOR2_X1 port map( A => Cin, B => B0(3), Z => B(3));
   U8 : XOR2_X1 port map( A => Cin, B => B0(31), Z => B(31));
   U9 : XOR2_X1 port map( A => Cin, B => B0(30), Z => B(30));
   U10 : XOR2_X1 port map( A => Cin, B => B0(2), Z => B(2));
   U11 : XOR2_X1 port map( A => Cin, B => B0(29), Z => B(29));
   U12 : XOR2_X1 port map( A => Cin, B => B0(28), Z => B(28));
   U13 : XOR2_X1 port map( A => Cin, B => B0(27), Z => B(27));
   U14 : XOR2_X1 port map( A => Cin, B => B0(26), Z => B(26));
   U15 : XOR2_X1 port map( A => Cin, B => B0(25), Z => B(25));
   U16 : XOR2_X1 port map( A => Cin, B => B0(24), Z => B(24));
   U17 : XOR2_X1 port map( A => Cin, B => B0(23), Z => B(23));
   U18 : XOR2_X1 port map( A => Cin, B => B0(22), Z => B(22));
   U19 : XOR2_X1 port map( A => Cin, B => B0(21), Z => B(21));
   U20 : XOR2_X1 port map( A => Cin, B => B0(20), Z => B(20));
   U21 : XOR2_X1 port map( A => Cin, B => B0(1), Z => B(1));
   U22 : XOR2_X1 port map( A => Cin, B => B0(19), Z => B(19));
   U23 : XOR2_X1 port map( A => Cin, B => B0(18), Z => B(18));
   U24 : XOR2_X1 port map( A => Cin, B => B0(17), Z => B(17));
   U25 : XOR2_X1 port map( A => Cin, B => B0(16), Z => B(16));
   U26 : XOR2_X1 port map( A => Cin, B => B0(15), Z => B(15));
   U27 : XOR2_X1 port map( A => Cin, B => B0(14), Z => B(14));
   U28 : XOR2_X1 port map( A => Cin, B => B0(13), Z => B(13));
   U29 : XOR2_X1 port map( A => Cin, B => B0(12), Z => B(12));
   U30 : XOR2_X1 port map( A => Cin, B => B0(11), Z => B(11));
   U31 : XOR2_X1 port map( A => Cin, B => B0(10), Z => B(10));
   U32 : XOR2_X1 port map( A => Cin, B => B0(0), Z => B(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity logic_and_shift_N32 is

   port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
         downto 0));

end logic_and_shift_N32;

architecture SYN_BEHAVIOR of logic_and_shift_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component logic_and_shift_N32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component logic_and_shift_N32_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (30 downto 0);  SH_TC : in std_logic;  B : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,
      N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57
      , N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, 
      N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86
      , N87, N88, N89, N90, N91, N92, N190, N191, N192, N193, N194, N195, N196,
      N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, 
      N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, 
      N221, n3, n4, n207_port, n208_port, n209_port, n210_port, n211_port, 
      n212_port, n213_port, n214_port, n215_port, n216_port, n217_port, 
      n218_port, n219_port, n220_port, n221_port, n222, n223, n224, n225, n226,
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
      n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
      n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, 
      n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, 
      n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, 
      n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, 
      n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, 
      n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, 
      n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, 
      n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, 
      n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
      n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
      n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
      n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, 
      n407, n408, n409, n410 : std_logic;

begin
   
   OUTALU_reg_31_inst : DLH_X1 port map( G => n208_port, D => N221, Q => 
                           OUTALU(31));
   OUTALU_reg_30_inst : DLH_X1 port map( G => n208_port, D => N220, Q => 
                           OUTALU(30));
   OUTALU_reg_29_inst : DLH_X1 port map( G => n208_port, D => N219, Q => 
                           OUTALU(29));
   OUTALU_reg_28_inst : DLH_X1 port map( G => n208_port, D => N218, Q => 
                           OUTALU(28));
   OUTALU_reg_27_inst : DLH_X1 port map( G => n208_port, D => N217, Q => 
                           OUTALU(27));
   OUTALU_reg_26_inst : DLH_X1 port map( G => n208_port, D => N216, Q => 
                           OUTALU(26));
   OUTALU_reg_25_inst : DLH_X1 port map( G => n208_port, D => N215, Q => 
                           OUTALU(25));
   OUTALU_reg_24_inst : DLH_X1 port map( G => n208_port, D => N214, Q => 
                           OUTALU(24));
   OUTALU_reg_23_inst : DLH_X1 port map( G => n208_port, D => N213, Q => 
                           OUTALU(23));
   OUTALU_reg_22_inst : DLH_X1 port map( G => n208_port, D => N212, Q => 
                           OUTALU(22));
   OUTALU_reg_21_inst : DLH_X1 port map( G => n208_port, D => N211, Q => 
                           OUTALU(21));
   OUTALU_reg_20_inst : DLH_X1 port map( G => n208_port, D => N210, Q => 
                           OUTALU(20));
   OUTALU_reg_19_inst : DLH_X1 port map( G => n208_port, D => N209, Q => 
                           OUTALU(19));
   OUTALU_reg_18_inst : DLH_X1 port map( G => n208_port, D => N208, Q => 
                           OUTALU(18));
   OUTALU_reg_17_inst : DLH_X1 port map( G => n208_port, D => N207, Q => 
                           OUTALU(17));
   OUTALU_reg_16_inst : DLH_X1 port map( G => n208_port, D => N206, Q => 
                           OUTALU(16));
   OUTALU_reg_15_inst : DLH_X1 port map( G => n208_port, D => N205, Q => 
                           OUTALU(15));
   OUTALU_reg_14_inst : DLH_X1 port map( G => n208_port, D => N204, Q => 
                           OUTALU(14));
   OUTALU_reg_13_inst : DLH_X1 port map( G => n208_port, D => N203, Q => 
                           OUTALU(13));
   OUTALU_reg_12_inst : DLH_X1 port map( G => n208_port, D => N202, Q => 
                           OUTALU(12));
   OUTALU_reg_11_inst : DLH_X1 port map( G => n208_port, D => N201, Q => 
                           OUTALU(11));
   OUTALU_reg_10_inst : DLH_X1 port map( G => n208_port, D => N200, Q => 
                           OUTALU(10));
   OUTALU_reg_9_inst : DLH_X1 port map( G => n208_port, D => N199, Q => 
                           OUTALU(9));
   OUTALU_reg_8_inst : DLH_X1 port map( G => n208_port, D => N198, Q => 
                           OUTALU(8));
   OUTALU_reg_7_inst : DLH_X1 port map( G => n208_port, D => N197, Q => 
                           OUTALU(7));
   OUTALU_reg_6_inst : DLH_X1 port map( G => n208_port, D => N196, Q => 
                           OUTALU(6));
   OUTALU_reg_5_inst : DLH_X1 port map( G => n208_port, D => N195, Q => 
                           OUTALU(5));
   OUTALU_reg_4_inst : DLH_X1 port map( G => n208_port, D => N194, Q => 
                           OUTALU(4));
   OUTALU_reg_3_inst : DLH_X1 port map( G => n208_port, D => N193, Q => 
                           OUTALU(3));
   OUTALU_reg_2_inst : DLH_X1 port map( G => n208_port, D => N192, Q => 
                           OUTALU(2));
   OUTALU_reg_1_inst : DLH_X1 port map( G => n208_port, D => N191, Q => 
                           OUTALU(1));
   OUTALU_reg_0_inst : DLH_X1 port map( G => n208_port, D => N190, Q => 
                           OUTALU(0));
   n3 <= '0';
   n4 <= '0';
   srl_39 : logic_and_shift_N32_DW_rash_0 port map( A(31) => DATA1(31), A(30) 
                           => DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28)
                           , A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), DATA_TC => n3,
                           SH(30) => DATA2(30), SH(29) => DATA2(29), SH(28) => 
                           DATA2(28), SH(27) => DATA2(27), SH(26) => DATA2(26),
                           SH(25) => DATA2(25), SH(24) => DATA2(24), SH(23) => 
                           DATA2(23), SH(22) => DATA2(22), SH(21) => DATA2(21),
                           SH(20) => DATA2(20), SH(19) => DATA2(19), SH(18) => 
                           DATA2(18), SH(17) => DATA2(17), SH(16) => DATA2(16),
                           SH(15) => DATA2(15), SH(14) => DATA2(14), SH(13) => 
                           DATA2(13), SH(12) => DATA2(12), SH(11) => DATA2(11),
                           SH(10) => DATA2(10), SH(9) => DATA2(9), SH(8) => 
                           DATA2(8), SH(7) => DATA2(7), SH(6) => DATA2(6), 
                           SH(5) => DATA2(5), SH(4) => DATA2(4), SH(3) => 
                           DATA2(3), SH(2) => DATA2(2), SH(1) => DATA2(1), 
                           SH(0) => DATA2(0), SH_TC => n3, B(31) => N92, B(30) 
                           => N91, B(29) => N90, B(28) => N89, B(27) => N88, 
                           B(26) => N87, B(25) => N86, B(24) => N85, B(23) => 
                           N84, B(22) => N83, B(21) => N82, B(20) => N81, B(19)
                           => N80, B(18) => N79, B(17) => N78, B(16) => N77, 
                           B(15) => N76, B(14) => N75, B(13) => N74, B(12) => 
                           N73, B(11) => N72, B(10) => N71, B(9) => N70, B(8) 
                           => N69, B(7) => N68, B(6) => N67, B(5) => N66, B(4) 
                           => N65, B(3) => N64, B(2) => N63, B(1) => N62, B(0) 
                           => N61);
   sll_37 : logic_and_shift_N32_DW01_ash_0 port map( A(31) => DATA1(31), A(30) 
                           => DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28)
                           , A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), DATA_TC => n4,
                           SH(30) => DATA2(30), SH(29) => DATA2(29), SH(28) => 
                           DATA2(28), SH(27) => DATA2(27), SH(26) => DATA2(26),
                           SH(25) => DATA2(25), SH(24) => DATA2(24), SH(23) => 
                           DATA2(23), SH(22) => DATA2(22), SH(21) => DATA2(21),
                           SH(20) => DATA2(20), SH(19) => DATA2(19), SH(18) => 
                           DATA2(18), SH(17) => DATA2(17), SH(16) => DATA2(16),
                           SH(15) => DATA2(15), SH(14) => DATA2(14), SH(13) => 
                           DATA2(13), SH(12) => DATA2(12), SH(11) => DATA2(11),
                           SH(10) => DATA2(10), SH(9) => DATA2(9), SH(8) => 
                           DATA2(8), SH(7) => DATA2(7), SH(6) => DATA2(6), 
                           SH(5) => DATA2(5), SH(4) => DATA2(4), SH(3) => 
                           DATA2(3), SH(2) => DATA2(2), SH(1) => DATA2(1), 
                           SH(0) => DATA2(0), SH_TC => n4, B(31) => N60, B(30) 
                           => N59, B(29) => N58, B(28) => N57, B(27) => N56, 
                           B(26) => N55, B(25) => N54, B(24) => N53, B(23) => 
                           N52, B(22) => N51, B(21) => N50, B(20) => N49, B(19)
                           => N48, B(18) => N47, B(17) => N46, B(16) => N45, 
                           B(15) => N44, B(14) => N43, B(13) => N42, B(12) => 
                           N41, B(11) => N40, B(10) => N39, B(9) => N38, B(8) 
                           => N37, B(7) => N36, B(6) => N35, B(5) => N34, B(4) 
                           => N33, B(3) => N32, B(2) => N31, B(1) => N30, B(0) 
                           => N29);
   U5 : OR2_X1 port map( A1 => FUNC(0), A2 => n211_port, ZN => n207_port);
   U6 : INV_X1 port map( A => n207_port, ZN => n208_port);
   U7 : AND2_X4 port map( A1 => n213_port, A2 => FUNC(3), ZN => n220_port);
   U8 : AND3_X4 port map( A1 => FUNC(2), A2 => n407, A3 => FUNC(1), ZN => 
                           n212_port);
   U9 : NOR2_X4 port map( A1 => n410, A2 => FUNC(2), ZN => n213_port);
   U10 : OR3_X1 port map( A1 => FUNC(2), A2 => FUNC(1), A3 => n407, ZN => 
                           n214_port);
   U11 : INV_X2 port map( A => n214_port, ZN => n209_port);
   U12 : OR3_X1 port map( A1 => FUNC(2), A2 => FUNC(1), A3 => FUNC(3), ZN => 
                           n215_port);
   U13 : INV_X2 port map( A => n215_port, ZN => n210_port);
   U14 : NOR4_X1 port map( A1 => n212_port, A2 => n213_port, A3 => n209_port, 
                           A4 => n210_port, ZN => n211_port);
   U15 : OAI211_X1 port map( C1 => n216_port, C2 => n217_port, A => n218_port, 
                           B => n219_port, ZN => N221);
   U16 : AOI22_X1 port map( A1 => N60, A2 => n210_port, B1 => N92, B2 => 
                           n209_port, ZN => n219_port);
   U17 : OAI21_X1 port map( B1 => n220_port, B2 => n221_port, A => DATA2(31), 
                           ZN => n218_port);
   U18 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(31), Z =>
                           n221_port);
   U19 : INV_X1 port map( A => DATA1(31), ZN => n217_port);
   U20 : AOI21_X1 port map( B1 => n212_port, B2 => n222, A => n220_port, ZN => 
                           n216_port);
   U21 : INV_X1 port map( A => DATA2(31), ZN => n222);
   U22 : OAI211_X1 port map( C1 => n223, C2 => n224, A => n225, B => n226, ZN 
                           => N220);
   U23 : AOI22_X1 port map( A1 => N59, A2 => n210_port, B1 => N91, B2 => 
                           n209_port, ZN => n226);
   U24 : OAI21_X1 port map( B1 => n220_port, B2 => n227, A => DATA2(30), ZN => 
                           n225);
   U25 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(30), Z =>
                           n227);
   U26 : INV_X1 port map( A => DATA1(30), ZN => n224);
   U27 : AOI21_X1 port map( B1 => n212_port, B2 => n228, A => n220_port, ZN => 
                           n223);
   U28 : INV_X1 port map( A => DATA2(30), ZN => n228);
   U29 : OAI211_X1 port map( C1 => n229, C2 => n230, A => n231, B => n232, ZN 
                           => N219);
   U30 : AOI22_X1 port map( A1 => N58, A2 => n210_port, B1 => N90, B2 => 
                           n209_port, ZN => n232);
   U31 : OAI21_X1 port map( B1 => n220_port, B2 => n233, A => DATA2(29), ZN => 
                           n231);
   U32 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(29), Z =>
                           n233);
   U33 : INV_X1 port map( A => DATA1(29), ZN => n230);
   U34 : AOI21_X1 port map( B1 => n212_port, B2 => n234, A => n220_port, ZN => 
                           n229);
   U35 : INV_X1 port map( A => DATA2(29), ZN => n234);
   U36 : OAI211_X1 port map( C1 => n235, C2 => n236, A => n237, B => n238, ZN 
                           => N218);
   U37 : AOI22_X1 port map( A1 => N57, A2 => n210_port, B1 => N89, B2 => 
                           n209_port, ZN => n238);
   U38 : OAI21_X1 port map( B1 => n220_port, B2 => n239, A => DATA2(28), ZN => 
                           n237);
   U39 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(28), Z =>
                           n239);
   U40 : INV_X1 port map( A => DATA1(28), ZN => n236);
   U41 : AOI21_X1 port map( B1 => n212_port, B2 => n240, A => n220_port, ZN => 
                           n235);
   U42 : INV_X1 port map( A => DATA2(28), ZN => n240);
   U43 : OAI211_X1 port map( C1 => n241, C2 => n242, A => n243, B => n244, ZN 
                           => N217);
   U44 : AOI22_X1 port map( A1 => N56, A2 => n210_port, B1 => N88, B2 => 
                           n209_port, ZN => n244);
   U45 : OAI21_X1 port map( B1 => n220_port, B2 => n245, A => DATA2(27), ZN => 
                           n243);
   U46 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(27), Z =>
                           n245);
   U47 : INV_X1 port map( A => DATA1(27), ZN => n242);
   U48 : AOI21_X1 port map( B1 => n212_port, B2 => n246, A => n220_port, ZN => 
                           n241);
   U49 : INV_X1 port map( A => DATA2(27), ZN => n246);
   U50 : OAI211_X1 port map( C1 => n247, C2 => n248, A => n249, B => n250, ZN 
                           => N216);
   U51 : AOI22_X1 port map( A1 => N55, A2 => n210_port, B1 => N87, B2 => 
                           n209_port, ZN => n250);
   U52 : OAI21_X1 port map( B1 => n220_port, B2 => n251, A => DATA2(26), ZN => 
                           n249);
   U53 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(26), Z =>
                           n251);
   U54 : INV_X1 port map( A => DATA1(26), ZN => n248);
   U55 : AOI21_X1 port map( B1 => n212_port, B2 => n252, A => n220_port, ZN => 
                           n247);
   U56 : INV_X1 port map( A => DATA2(26), ZN => n252);
   U57 : OAI211_X1 port map( C1 => n253, C2 => n254, A => n255, B => n256, ZN 
                           => N215);
   U58 : AOI22_X1 port map( A1 => N54, A2 => n210_port, B1 => N86, B2 => 
                           n209_port, ZN => n256);
   U59 : OAI21_X1 port map( B1 => n220_port, B2 => n257, A => DATA2(25), ZN => 
                           n255);
   U60 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(25), Z =>
                           n257);
   U61 : INV_X1 port map( A => DATA1(25), ZN => n254);
   U62 : AOI21_X1 port map( B1 => n212_port, B2 => n258, A => n220_port, ZN => 
                           n253);
   U63 : INV_X1 port map( A => DATA2(25), ZN => n258);
   U64 : OAI211_X1 port map( C1 => n259, C2 => n260, A => n261, B => n262, ZN 
                           => N214);
   U65 : AOI22_X1 port map( A1 => N53, A2 => n210_port, B1 => N85, B2 => 
                           n209_port, ZN => n262);
   U66 : OAI21_X1 port map( B1 => n220_port, B2 => n263, A => DATA2(24), ZN => 
                           n261);
   U67 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(24), Z =>
                           n263);
   U68 : INV_X1 port map( A => DATA1(24), ZN => n260);
   U69 : AOI21_X1 port map( B1 => n212_port, B2 => n264, A => n220_port, ZN => 
                           n259);
   U70 : INV_X1 port map( A => DATA2(24), ZN => n264);
   U71 : OAI211_X1 port map( C1 => n265, C2 => n266, A => n267, B => n268, ZN 
                           => N213);
   U72 : AOI22_X1 port map( A1 => N52, A2 => n210_port, B1 => N84, B2 => 
                           n209_port, ZN => n268);
   U73 : OAI21_X1 port map( B1 => n220_port, B2 => n269, A => DATA2(23), ZN => 
                           n267);
   U74 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(23), Z =>
                           n269);
   U75 : INV_X1 port map( A => DATA1(23), ZN => n266);
   U76 : AOI21_X1 port map( B1 => n212_port, B2 => n270, A => n220_port, ZN => 
                           n265);
   U77 : INV_X1 port map( A => DATA2(23), ZN => n270);
   U78 : OAI211_X1 port map( C1 => n271, C2 => n272, A => n273, B => n274, ZN 
                           => N212);
   U79 : AOI22_X1 port map( A1 => N51, A2 => n210_port, B1 => N83, B2 => 
                           n209_port, ZN => n274);
   U80 : OAI21_X1 port map( B1 => n220_port, B2 => n275, A => DATA2(22), ZN => 
                           n273);
   U81 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(22), Z =>
                           n275);
   U82 : INV_X1 port map( A => DATA1(22), ZN => n272);
   U83 : AOI21_X1 port map( B1 => n212_port, B2 => n276, A => n220_port, ZN => 
                           n271);
   U84 : INV_X1 port map( A => DATA2(22), ZN => n276);
   U85 : OAI211_X1 port map( C1 => n277, C2 => n278, A => n279, B => n280, ZN 
                           => N211);
   U86 : AOI22_X1 port map( A1 => N50, A2 => n210_port, B1 => N82, B2 => 
                           n209_port, ZN => n280);
   U87 : OAI21_X1 port map( B1 => n220_port, B2 => n281, A => DATA2(21), ZN => 
                           n279);
   U88 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(21), Z =>
                           n281);
   U89 : INV_X1 port map( A => DATA1(21), ZN => n278);
   U90 : AOI21_X1 port map( B1 => n212_port, B2 => n282, A => n220_port, ZN => 
                           n277);
   U91 : INV_X1 port map( A => DATA2(21), ZN => n282);
   U92 : OAI211_X1 port map( C1 => n283, C2 => n284, A => n285, B => n286, ZN 
                           => N210);
   U93 : AOI22_X1 port map( A1 => N49, A2 => n210_port, B1 => N81, B2 => 
                           n209_port, ZN => n286);
   U94 : OAI21_X1 port map( B1 => n220_port, B2 => n287, A => DATA2(20), ZN => 
                           n285);
   U95 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(20), Z =>
                           n287);
   U96 : INV_X1 port map( A => DATA1(20), ZN => n284);
   U97 : AOI21_X1 port map( B1 => n212_port, B2 => n288, A => n220_port, ZN => 
                           n283);
   U98 : INV_X1 port map( A => DATA2(20), ZN => n288);
   U99 : OAI211_X1 port map( C1 => n289, C2 => n290, A => n291, B => n292, ZN 
                           => N209);
   U100 : AOI22_X1 port map( A1 => N48, A2 => n210_port, B1 => N80, B2 => 
                           n209_port, ZN => n292);
   U101 : OAI21_X1 port map( B1 => n220_port, B2 => n293, A => DATA2(19), ZN =>
                           n291);
   U102 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(19), Z 
                           => n293);
   U103 : INV_X1 port map( A => DATA1(19), ZN => n290);
   U104 : AOI21_X1 port map( B1 => n212_port, B2 => n294, A => n220_port, ZN =>
                           n289);
   U105 : INV_X1 port map( A => DATA2(19), ZN => n294);
   U106 : OAI211_X1 port map( C1 => n295, C2 => n296, A => n297, B => n298, ZN 
                           => N208);
   U107 : AOI22_X1 port map( A1 => N47, A2 => n210_port, B1 => N79, B2 => 
                           n209_port, ZN => n298);
   U108 : OAI21_X1 port map( B1 => n220_port, B2 => n299, A => DATA2(18), ZN =>
                           n297);
   U109 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(18), Z 
                           => n299);
   U110 : INV_X1 port map( A => DATA1(18), ZN => n296);
   U111 : AOI21_X1 port map( B1 => n212_port, B2 => n300, A => n220_port, ZN =>
                           n295);
   U112 : INV_X1 port map( A => DATA2(18), ZN => n300);
   U113 : OAI211_X1 port map( C1 => n301, C2 => n302, A => n303, B => n304, ZN 
                           => N207);
   U114 : AOI22_X1 port map( A1 => N46, A2 => n210_port, B1 => N78, B2 => 
                           n209_port, ZN => n304);
   U115 : OAI21_X1 port map( B1 => n220_port, B2 => n305, A => DATA2(17), ZN =>
                           n303);
   U116 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(17), Z 
                           => n305);
   U117 : INV_X1 port map( A => DATA1(17), ZN => n302);
   U118 : AOI21_X1 port map( B1 => n212_port, B2 => n306, A => n220_port, ZN =>
                           n301);
   U119 : INV_X1 port map( A => DATA2(17), ZN => n306);
   U120 : OAI211_X1 port map( C1 => n307, C2 => n308, A => n309, B => n310, ZN 
                           => N206);
   U121 : AOI22_X1 port map( A1 => N45, A2 => n210_port, B1 => N77, B2 => 
                           n209_port, ZN => n310);
   U122 : OAI21_X1 port map( B1 => n220_port, B2 => n311, A => DATA2(16), ZN =>
                           n309);
   U123 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(16), Z 
                           => n311);
   U124 : INV_X1 port map( A => DATA1(16), ZN => n308);
   U125 : AOI21_X1 port map( B1 => n212_port, B2 => n312, A => n220_port, ZN =>
                           n307);
   U126 : INV_X1 port map( A => DATA2(16), ZN => n312);
   U127 : OAI211_X1 port map( C1 => n313, C2 => n314, A => n315, B => n316, ZN 
                           => N205);
   U128 : AOI22_X1 port map( A1 => N44, A2 => n210_port, B1 => N76, B2 => 
                           n209_port, ZN => n316);
   U129 : OAI21_X1 port map( B1 => n220_port, B2 => n317, A => DATA2(15), ZN =>
                           n315);
   U130 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(15), Z 
                           => n317);
   U131 : INV_X1 port map( A => DATA1(15), ZN => n314);
   U132 : AOI21_X1 port map( B1 => n212_port, B2 => n318, A => n220_port, ZN =>
                           n313);
   U133 : INV_X1 port map( A => DATA2(15), ZN => n318);
   U134 : OAI211_X1 port map( C1 => n319, C2 => n320, A => n321, B => n322, ZN 
                           => N204);
   U135 : AOI22_X1 port map( A1 => N43, A2 => n210_port, B1 => N75, B2 => 
                           n209_port, ZN => n322);
   U136 : OAI21_X1 port map( B1 => n220_port, B2 => n323, A => DATA2(14), ZN =>
                           n321);
   U137 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(14), Z 
                           => n323);
   U138 : INV_X1 port map( A => DATA1(14), ZN => n320);
   U139 : AOI21_X1 port map( B1 => n212_port, B2 => n324, A => n220_port, ZN =>
                           n319);
   U140 : INV_X1 port map( A => DATA2(14), ZN => n324);
   U141 : OAI211_X1 port map( C1 => n325, C2 => n326, A => n327, B => n328, ZN 
                           => N203);
   U142 : AOI22_X1 port map( A1 => N42, A2 => n210_port, B1 => N74, B2 => 
                           n209_port, ZN => n328);
   U143 : OAI21_X1 port map( B1 => n220_port, B2 => n329, A => DATA2(13), ZN =>
                           n327);
   U144 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(13), Z 
                           => n329);
   U145 : INV_X1 port map( A => DATA1(13), ZN => n326);
   U146 : AOI21_X1 port map( B1 => n212_port, B2 => n330, A => n220_port, ZN =>
                           n325);
   U147 : INV_X1 port map( A => DATA2(13), ZN => n330);
   U148 : OAI211_X1 port map( C1 => n331, C2 => n332, A => n333, B => n334, ZN 
                           => N202);
   U149 : AOI22_X1 port map( A1 => N41, A2 => n210_port, B1 => N73, B2 => 
                           n209_port, ZN => n334);
   U150 : OAI21_X1 port map( B1 => n220_port, B2 => n335, A => DATA2(12), ZN =>
                           n333);
   U151 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(12), Z 
                           => n335);
   U152 : INV_X1 port map( A => DATA1(12), ZN => n332);
   U153 : AOI21_X1 port map( B1 => n212_port, B2 => n336, A => n220_port, ZN =>
                           n331);
   U154 : INV_X1 port map( A => DATA2(12), ZN => n336);
   U155 : OAI211_X1 port map( C1 => n337, C2 => n338, A => n339, B => n340, ZN 
                           => N201);
   U156 : AOI22_X1 port map( A1 => N40, A2 => n210_port, B1 => N72, B2 => 
                           n209_port, ZN => n340);
   U157 : OAI21_X1 port map( B1 => n220_port, B2 => n341, A => DATA2(11), ZN =>
                           n339);
   U158 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(11), Z 
                           => n341);
   U159 : INV_X1 port map( A => DATA1(11), ZN => n338);
   U160 : AOI21_X1 port map( B1 => n212_port, B2 => n342, A => n220_port, ZN =>
                           n337);
   U161 : INV_X1 port map( A => DATA2(11), ZN => n342);
   U162 : OAI211_X1 port map( C1 => n343, C2 => n344, A => n345, B => n346, ZN 
                           => N200);
   U163 : AOI22_X1 port map( A1 => N39, A2 => n210_port, B1 => N71, B2 => 
                           n209_port, ZN => n346);
   U164 : OAI21_X1 port map( B1 => n220_port, B2 => n347, A => DATA2(10), ZN =>
                           n345);
   U165 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(10), Z 
                           => n347);
   U166 : INV_X1 port map( A => DATA1(10), ZN => n344);
   U167 : AOI21_X1 port map( B1 => n212_port, B2 => n348, A => n220_port, ZN =>
                           n343);
   U168 : INV_X1 port map( A => DATA2(10), ZN => n348);
   U169 : OAI211_X1 port map( C1 => n349, C2 => n350, A => n351, B => n352, ZN 
                           => N199);
   U170 : AOI22_X1 port map( A1 => N38, A2 => n210_port, B1 => N70, B2 => 
                           n209_port, ZN => n352);
   U171 : OAI21_X1 port map( B1 => n220_port, B2 => n353, A => DATA2(9), ZN => 
                           n351);
   U172 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(9), Z =>
                           n353);
   U173 : INV_X1 port map( A => DATA1(9), ZN => n350);
   U174 : AOI21_X1 port map( B1 => n212_port, B2 => n354, A => n220_port, ZN =>
                           n349);
   U175 : INV_X1 port map( A => DATA2(9), ZN => n354);
   U176 : OAI211_X1 port map( C1 => n355, C2 => n356, A => n357, B => n358, ZN 
                           => N198);
   U177 : AOI22_X1 port map( A1 => N37, A2 => n210_port, B1 => N69, B2 => 
                           n209_port, ZN => n358);
   U178 : OAI21_X1 port map( B1 => n220_port, B2 => n359, A => DATA2(8), ZN => 
                           n357);
   U179 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(8), Z =>
                           n359);
   U180 : INV_X1 port map( A => DATA1(8), ZN => n356);
   U181 : AOI21_X1 port map( B1 => n212_port, B2 => n360, A => n220_port, ZN =>
                           n355);
   U182 : INV_X1 port map( A => DATA2(8), ZN => n360);
   U183 : OAI211_X1 port map( C1 => n361, C2 => n362, A => n363, B => n364, ZN 
                           => N197);
   U184 : AOI22_X1 port map( A1 => N36, A2 => n210_port, B1 => N68, B2 => 
                           n209_port, ZN => n364);
   U185 : OAI21_X1 port map( B1 => n220_port, B2 => n365, A => DATA2(7), ZN => 
                           n363);
   U186 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(7), Z =>
                           n365);
   U187 : INV_X1 port map( A => DATA1(7), ZN => n362);
   U188 : AOI21_X1 port map( B1 => n212_port, B2 => n366, A => n220_port, ZN =>
                           n361);
   U189 : INV_X1 port map( A => DATA2(7), ZN => n366);
   U190 : OAI211_X1 port map( C1 => n367, C2 => n368, A => n369, B => n370, ZN 
                           => N196);
   U191 : AOI22_X1 port map( A1 => N35, A2 => n210_port, B1 => N67, B2 => 
                           n209_port, ZN => n370);
   U192 : OAI21_X1 port map( B1 => n220_port, B2 => n371, A => DATA2(6), ZN => 
                           n369);
   U193 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(6), Z =>
                           n371);
   U194 : INV_X1 port map( A => DATA1(6), ZN => n368);
   U195 : AOI21_X1 port map( B1 => n212_port, B2 => n372, A => n220_port, ZN =>
                           n367);
   U196 : INV_X1 port map( A => DATA2(6), ZN => n372);
   U197 : OAI211_X1 port map( C1 => n373, C2 => n374, A => n375, B => n376, ZN 
                           => N195);
   U198 : AOI22_X1 port map( A1 => N34, A2 => n210_port, B1 => N66, B2 => 
                           n209_port, ZN => n376);
   U199 : OAI21_X1 port map( B1 => n220_port, B2 => n377, A => DATA2(5), ZN => 
                           n375);
   U200 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(5), Z =>
                           n377);
   U201 : INV_X1 port map( A => DATA1(5), ZN => n374);
   U202 : AOI21_X1 port map( B1 => n212_port, B2 => n378, A => n220_port, ZN =>
                           n373);
   U203 : INV_X1 port map( A => DATA2(5), ZN => n378);
   U204 : OAI211_X1 port map( C1 => n379, C2 => n380, A => n381, B => n382, ZN 
                           => N194);
   U205 : AOI22_X1 port map( A1 => N33, A2 => n210_port, B1 => N65, B2 => 
                           n209_port, ZN => n382);
   U206 : OAI21_X1 port map( B1 => n220_port, B2 => n383, A => DATA2(4), ZN => 
                           n381);
   U207 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(4), Z =>
                           n383);
   U208 : INV_X1 port map( A => DATA1(4), ZN => n380);
   U209 : AOI21_X1 port map( B1 => n212_port, B2 => n384, A => n220_port, ZN =>
                           n379);
   U210 : INV_X1 port map( A => DATA2(4), ZN => n384);
   U211 : OAI211_X1 port map( C1 => n385, C2 => n386, A => n387, B => n388, ZN 
                           => N193);
   U212 : AOI22_X1 port map( A1 => N32, A2 => n210_port, B1 => N64, B2 => 
                           n209_port, ZN => n388);
   U213 : OAI21_X1 port map( B1 => n220_port, B2 => n389, A => DATA2(3), ZN => 
                           n387);
   U214 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(3), Z =>
                           n389);
   U215 : INV_X1 port map( A => DATA1(3), ZN => n386);
   U216 : AOI21_X1 port map( B1 => n212_port, B2 => n390, A => n220_port, ZN =>
                           n385);
   U217 : INV_X1 port map( A => DATA2(3), ZN => n390);
   U218 : OAI211_X1 port map( C1 => n391, C2 => n392, A => n393, B => n394, ZN 
                           => N192);
   U219 : AOI22_X1 port map( A1 => N31, A2 => n210_port, B1 => N63, B2 => 
                           n209_port, ZN => n394);
   U220 : OAI21_X1 port map( B1 => n220_port, B2 => n395, A => DATA2(2), ZN => 
                           n393);
   U221 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(2), Z =>
                           n395);
   U222 : INV_X1 port map( A => DATA1(2), ZN => n392);
   U223 : AOI21_X1 port map( B1 => n212_port, B2 => n396, A => n220_port, ZN =>
                           n391);
   U224 : INV_X1 port map( A => DATA2(2), ZN => n396);
   U225 : OAI211_X1 port map( C1 => n397, C2 => n398, A => n399, B => n400, ZN 
                           => N191);
   U226 : AOI22_X1 port map( A1 => N30, A2 => n210_port, B1 => N62, B2 => 
                           n209_port, ZN => n400);
   U227 : OAI21_X1 port map( B1 => n220_port, B2 => n401, A => DATA2(1), ZN => 
                           n399);
   U228 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(1), Z =>
                           n401);
   U229 : INV_X1 port map( A => DATA1(1), ZN => n398);
   U230 : AOI21_X1 port map( B1 => n212_port, B2 => n402, A => n220_port, ZN =>
                           n397);
   U231 : INV_X1 port map( A => DATA2(1), ZN => n402);
   U232 : OAI211_X1 port map( C1 => n403, C2 => n404, A => n405, B => n406, ZN 
                           => N190);
   U233 : AOI22_X1 port map( A1 => N29, A2 => n210_port, B1 => N61, B2 => 
                           n209_port, ZN => n406);
   U234 : OAI21_X1 port map( B1 => n220_port, B2 => n408, A => DATA2(0), ZN => 
                           n405);
   U235 : MUX2_X1 port map( A => n212_port, B => n213_port, S => DATA1(0), Z =>
                           n408);
   U236 : INV_X1 port map( A => DATA1(0), ZN => n404);
   U237 : AOI21_X1 port map( B1 => n212_port, B2 => n409, A => n220_port, ZN =>
                           n403);
   U238 : INV_X1 port map( A => FUNC(1), ZN => n410);
   U239 : INV_X1 port map( A => DATA2(0), ZN => n409);
   U240 : INV_X1 port map( A => FUNC(3), ZN => n407);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity P4_ADDER_NBITS32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end P4_ADDER_NBITS32;

architecture SYN_STRUCTURAL of P4_ADDER_NBITS32 is

   component CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4
      port( A, B : in std_logic_vector (32 downto 1);  C0 : in std_logic;  COUT
            : out std_logic_vector (8 downto 0));
   end component;
   
   component SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (8 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component xor_logic_nbits32
      port( Cin : in std_logic;  B0 : in std_logic_vector (31 downto 0);  B : 
            out std_logic_vector (31 downto 0));
   end component;
   
   signal Co_port, B_diff_31_port, B_diff_30_port, B_diff_29_port, 
      B_diff_28_port, B_diff_27_port, B_diff_26_port, B_diff_25_port, 
      B_diff_24_port, B_diff_23_port, B_diff_22_port, B_diff_21_port, 
      B_diff_20_port, B_diff_19_port, B_diff_18_port, B_diff_17_port, 
      B_diff_16_port, B_diff_15_port, B_diff_14_port, B_diff_13_port, 
      B_diff_12_port, B_diff_11_port, B_diff_10_port, B_diff_9_port, 
      B_diff_8_port, B_diff_7_port, B_diff_6_port, B_diff_5_port, B_diff_4_port
      , B_diff_3_port, B_diff_2_port, B_diff_1_port, B_diff_0_port, 
      fromCarry_to_adder_7_port, fromCarry_to_adder_6_port, 
      fromCarry_to_adder_5_port, fromCarry_to_adder_4_port, 
      fromCarry_to_adder_3_port, fromCarry_to_adder_2_port, 
      fromCarry_to_adder_1_port, fromCarry_to_adder_0_port : std_logic;

begin
   Co <= Co_port;
   
   xor_gate : xor_logic_nbits32 port map( Cin => Ci, B0(31) => B(31), B0(30) =>
                           B(30), B0(29) => B(29), B0(28) => B(28), B0(27) => 
                           B(27), B0(26) => B(26), B0(25) => B(25), B0(24) => 
                           B(24), B0(23) => B(23), B0(22) => B(22), B0(21) => 
                           B(21), B0(20) => B(20), B0(19) => B(19), B0(18) => 
                           B(18), B0(17) => B(17), B0(16) => B(16), B0(15) => 
                           B(15), B0(14) => B(14), B0(13) => B(13), B0(12) => 
                           B(12), B0(11) => B(11), B0(10) => B(10), B0(9) => 
                           B(9), B0(8) => B(8), B0(7) => B(7), B0(6) => B(6), 
                           B0(5) => B(5), B0(4) => B(4), B0(3) => B(3), B0(2) 
                           => B(2), B0(1) => B(1), B0(0) => B(0), B(31) => 
                           B_diff_31_port, B(30) => B_diff_30_port, B(29) => 
                           B_diff_29_port, B(28) => B_diff_28_port, B(27) => 
                           B_diff_27_port, B(26) => B_diff_26_port, B(25) => 
                           B_diff_25_port, B(24) => B_diff_24_port, B(23) => 
                           B_diff_23_port, B(22) => B_diff_22_port, B(21) => 
                           B_diff_21_port, B(20) => B_diff_20_port, B(19) => 
                           B_diff_19_port, B(18) => B_diff_18_port, B(17) => 
                           B_diff_17_port, B(16) => B_diff_16_port, B(15) => 
                           B_diff_15_port, B(14) => B_diff_14_port, B(13) => 
                           B_diff_13_port, B(12) => B_diff_12_port, B(11) => 
                           B_diff_11_port, B(10) => B_diff_10_port, B(9) => 
                           B_diff_9_port, B(8) => B_diff_8_port, B(7) => 
                           B_diff_7_port, B(6) => B_diff_6_port, B(5) => 
                           B_diff_5_port, B(4) => B_diff_4_port, B(3) => 
                           B_diff_3_port, B(2) => B_diff_2_port, B(1) => 
                           B_diff_1_port, B(0) => B_diff_0_port);
   SUM_GEN : SUMGENERATOR_NBITS32_BITS_PER_MODULE4_NUM_MODULES8 port map( A(31)
                           => A(31), A(30) => A(30), A(29) => A(29), A(28) => 
                           A(28), A(27) => A(27), A(26) => A(26), A(25) => 
                           A(25), A(24) => A(24), A(23) => A(23), A(22) => 
                           A(22), A(21) => A(21), A(20) => A(20), A(19) => 
                           A(19), A(18) => A(18), A(17) => A(17), A(16) => 
                           A(16), A(15) => A(15), A(14) => A(14), A(13) => 
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => B_diff_31_port, B(30) => B_diff_30_port, 
                           B(29) => B_diff_29_port, B(28) => B_diff_28_port, 
                           B(27) => B_diff_27_port, B(26) => B_diff_26_port, 
                           B(25) => B_diff_25_port, B(24) => B_diff_24_port, 
                           B(23) => B_diff_23_port, B(22) => B_diff_22_port, 
                           B(21) => B_diff_21_port, B(20) => B_diff_20_port, 
                           B(19) => B_diff_19_port, B(18) => B_diff_18_port, 
                           B(17) => B_diff_17_port, B(16) => B_diff_16_port, 
                           B(15) => B_diff_15_port, B(14) => B_diff_14_port, 
                           B(13) => B_diff_13_port, B(12) => B_diff_12_port, 
                           B(11) => B_diff_11_port, B(10) => B_diff_10_port, 
                           B(9) => B_diff_9_port, B(8) => B_diff_8_port, B(7) 
                           => B_diff_7_port, B(6) => B_diff_6_port, B(5) => 
                           B_diff_5_port, B(4) => B_diff_4_port, B(3) => 
                           B_diff_3_port, B(2) => B_diff_2_port, B(1) => 
                           B_diff_1_port, B(0) => B_diff_0_port, Ci(8) => 
                           Co_port, Ci(7) => fromCarry_to_adder_7_port, Ci(6) 
                           => fromCarry_to_adder_6_port, Ci(5) => 
                           fromCarry_to_adder_5_port, Ci(4) => 
                           fromCarry_to_adder_4_port, Ci(3) => 
                           fromCarry_to_adder_3_port, Ci(2) => 
                           fromCarry_to_adder_2_port, Ci(1) => 
                           fromCarry_to_adder_1_port, Ci(0) => 
                           fromCarry_to_adder_0_port, S(31) => S(31), S(30) => 
                           S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));
   CLA : CLA_SPARSE_TREE_NBITS32_NBITS_CARRIES4 port map( A(32) => A(31), A(31)
                           => A(30), A(30) => A(29), A(29) => A(28), A(28) => 
                           A(27), A(27) => A(26), A(26) => A(25), A(25) => 
                           A(24), A(24) => A(23), A(23) => A(22), A(22) => 
                           A(21), A(21) => A(20), A(20) => A(19), A(19) => 
                           A(18), A(18) => A(17), A(17) => A(16), A(16) => 
                           A(15), A(15) => A(14), A(14) => A(13), A(13) => 
                           A(12), A(12) => A(11), A(11) => A(10), A(10) => A(9)
                           , A(9) => A(8), A(8) => A(7), A(7) => A(6), A(6) => 
                           A(5), A(5) => A(4), A(4) => A(3), A(3) => A(2), A(2)
                           => A(1), A(1) => A(0), B(32) => B_diff_31_port, 
                           B(31) => B_diff_30_port, B(30) => B_diff_29_port, 
                           B(29) => B_diff_28_port, B(28) => B_diff_27_port, 
                           B(27) => B_diff_26_port, B(26) => B_diff_25_port, 
                           B(25) => B_diff_24_port, B(24) => B_diff_23_port, 
                           B(23) => B_diff_22_port, B(22) => B_diff_21_port, 
                           B(21) => B_diff_20_port, B(20) => B_diff_19_port, 
                           B(19) => B_diff_18_port, B(18) => B_diff_17_port, 
                           B(17) => B_diff_16_port, B(16) => B_diff_15_port, 
                           B(15) => B_diff_14_port, B(14) => B_diff_13_port, 
                           B(13) => B_diff_12_port, B(12) => B_diff_11_port, 
                           B(11) => B_diff_10_port, B(10) => B_diff_9_port, 
                           B(9) => B_diff_8_port, B(8) => B_diff_7_port, B(7) 
                           => B_diff_6_port, B(6) => B_diff_5_port, B(5) => 
                           B_diff_4_port, B(4) => B_diff_3_port, B(3) => 
                           B_diff_2_port, B(2) => B_diff_1_port, B(1) => 
                           B_diff_0_port, C0 => Ci, COUT(8) => Co_port, COUT(7)
                           => fromCarry_to_adder_7_port, COUT(6) => 
                           fromCarry_to_adder_6_port, COUT(5) => 
                           fromCarry_to_adder_5_port, COUT(4) => 
                           fromCarry_to_adder_4_port, COUT(3) => 
                           fromCarry_to_adder_3_port, COUT(2) => 
                           fromCarry_to_adder_2_port, COUT(1) => 
                           fromCarry_to_adder_1_port, COUT(0) => 
                           fromCarry_to_adder_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ctrl_alu_NBITS32 is

   port( A, B : in std_logic_vector (31 downto 0);  FUNC : in std_logic_vector 
         (0 to 3);  Ap4, Bp4 : out std_logic_vector (31 downto 0);  Cin : out 
         std_logic;  Als, Bls : out std_logic_vector (31 downto 0);  enableComp
         : out std_logic);

end ctrl_alu_NBITS32;

architecture SYN_BEHAVIORAL of ctrl_alu_NBITS32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
      n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104
      , n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152 : 
      std_logic;

begin
   
   U3 : INV_X1 port map( A => n76, ZN => n77);
   U4 : INV_X2 port map( A => n77, ZN => Cin);
   U5 : AND2_X4 port map( A1 => n81, A2 => n79, ZN => n82);
   U6 : NAND2_X4 port map( A1 => n151, A2 => n152, ZN => n115);
   U7 : INV_X1 port map( A => n79, ZN => enableComp);
   U8 : OAI21_X1 port map( B1 => n80, B2 => n81, A => n79, ZN => n76);
   U9 : NOR2_X1 port map( A1 => n82, A2 => n83, ZN => Bp4(9));
   U10 : NOR2_X1 port map( A1 => n82, A2 => n84, ZN => Bp4(8));
   U11 : NOR2_X1 port map( A1 => n82, A2 => n85, ZN => Bp4(7));
   U12 : NOR2_X1 port map( A1 => n82, A2 => n86, ZN => Bp4(6));
   U13 : NOR2_X1 port map( A1 => n82, A2 => n87, ZN => Bp4(5));
   U14 : NOR2_X1 port map( A1 => n82, A2 => n88, ZN => Bp4(4));
   U15 : NOR2_X1 port map( A1 => n82, A2 => n89, ZN => Bp4(3));
   U16 : NOR2_X1 port map( A1 => n82, A2 => n90, ZN => Bp4(31));
   U17 : NOR2_X1 port map( A1 => n82, A2 => n91, ZN => Bp4(30));
   U18 : NOR2_X1 port map( A1 => n82, A2 => n92, ZN => Bp4(2));
   U19 : NOR2_X1 port map( A1 => n82, A2 => n93, ZN => Bp4(29));
   U20 : NOR2_X1 port map( A1 => n82, A2 => n94, ZN => Bp4(28));
   U21 : NOR2_X1 port map( A1 => n82, A2 => n95, ZN => Bp4(27));
   U22 : NOR2_X1 port map( A1 => n82, A2 => n96, ZN => Bp4(26));
   U23 : NOR2_X1 port map( A1 => n82, A2 => n97, ZN => Bp4(25));
   U24 : NOR2_X1 port map( A1 => n82, A2 => n98, ZN => Bp4(24));
   U25 : NOR2_X1 port map( A1 => n82, A2 => n99, ZN => Bp4(23));
   U26 : NOR2_X1 port map( A1 => n82, A2 => n100, ZN => Bp4(22));
   U27 : NOR2_X1 port map( A1 => n82, A2 => n101, ZN => Bp4(21));
   U28 : NOR2_X1 port map( A1 => n82, A2 => n102, ZN => Bp4(20));
   U29 : NOR2_X1 port map( A1 => n82, A2 => n103, ZN => Bp4(1));
   U30 : NOR2_X1 port map( A1 => n82, A2 => n104, ZN => Bp4(19));
   U31 : NOR2_X1 port map( A1 => n82, A2 => n105, ZN => Bp4(18));
   U32 : NOR2_X1 port map( A1 => n82, A2 => n106, ZN => Bp4(17));
   U33 : NOR2_X1 port map( A1 => n82, A2 => n107, ZN => Bp4(16));
   U34 : NOR2_X1 port map( A1 => n82, A2 => n108, ZN => Bp4(15));
   U35 : NOR2_X1 port map( A1 => n82, A2 => n109, ZN => Bp4(14));
   U36 : NOR2_X1 port map( A1 => n82, A2 => n110, ZN => Bp4(13));
   U37 : NOR2_X1 port map( A1 => n82, A2 => n111, ZN => Bp4(12));
   U38 : NOR2_X1 port map( A1 => n82, A2 => n112, ZN => Bp4(11));
   U39 : NOR2_X1 port map( A1 => n82, A2 => n113, ZN => Bp4(10));
   U40 : NOR2_X1 port map( A1 => n82, A2 => n114, ZN => Bp4(0));
   U41 : NOR2_X1 port map( A1 => n83, A2 => n115, ZN => Bls(9));
   U42 : INV_X1 port map( A => B(9), ZN => n83);
   U43 : NOR2_X1 port map( A1 => n84, A2 => n115, ZN => Bls(8));
   U44 : INV_X1 port map( A => B(8), ZN => n84);
   U45 : NOR2_X1 port map( A1 => n85, A2 => n115, ZN => Bls(7));
   U46 : INV_X1 port map( A => B(7), ZN => n85);
   U47 : NOR2_X1 port map( A1 => n86, A2 => n115, ZN => Bls(6));
   U48 : INV_X1 port map( A => B(6), ZN => n86);
   U49 : NOR2_X1 port map( A1 => n87, A2 => n115, ZN => Bls(5));
   U50 : INV_X1 port map( A => B(5), ZN => n87);
   U51 : NOR2_X1 port map( A1 => n88, A2 => n115, ZN => Bls(4));
   U52 : INV_X1 port map( A => B(4), ZN => n88);
   U53 : NOR2_X1 port map( A1 => n89, A2 => n115, ZN => Bls(3));
   U54 : INV_X1 port map( A => B(3), ZN => n89);
   U55 : NOR2_X1 port map( A1 => n90, A2 => n115, ZN => Bls(31));
   U56 : INV_X1 port map( A => B(31), ZN => n90);
   U57 : NOR2_X1 port map( A1 => n91, A2 => n115, ZN => Bls(30));
   U58 : INV_X1 port map( A => B(30), ZN => n91);
   U59 : NOR2_X1 port map( A1 => n92, A2 => n115, ZN => Bls(2));
   U60 : INV_X1 port map( A => B(2), ZN => n92);
   U61 : NOR2_X1 port map( A1 => n93, A2 => n115, ZN => Bls(29));
   U62 : INV_X1 port map( A => B(29), ZN => n93);
   U63 : NOR2_X1 port map( A1 => n94, A2 => n115, ZN => Bls(28));
   U64 : INV_X1 port map( A => B(28), ZN => n94);
   U65 : NOR2_X1 port map( A1 => n95, A2 => n115, ZN => Bls(27));
   U66 : INV_X1 port map( A => B(27), ZN => n95);
   U67 : NOR2_X1 port map( A1 => n96, A2 => n115, ZN => Bls(26));
   U68 : INV_X1 port map( A => B(26), ZN => n96);
   U69 : NOR2_X1 port map( A1 => n97, A2 => n115, ZN => Bls(25));
   U70 : INV_X1 port map( A => B(25), ZN => n97);
   U71 : NOR2_X1 port map( A1 => n98, A2 => n115, ZN => Bls(24));
   U72 : INV_X1 port map( A => B(24), ZN => n98);
   U73 : NOR2_X1 port map( A1 => n99, A2 => n115, ZN => Bls(23));
   U74 : INV_X1 port map( A => B(23), ZN => n99);
   U75 : NOR2_X1 port map( A1 => n100, A2 => n115, ZN => Bls(22));
   U76 : INV_X1 port map( A => B(22), ZN => n100);
   U77 : NOR2_X1 port map( A1 => n101, A2 => n115, ZN => Bls(21));
   U78 : INV_X1 port map( A => B(21), ZN => n101);
   U79 : NOR2_X1 port map( A1 => n102, A2 => n115, ZN => Bls(20));
   U80 : INV_X1 port map( A => B(20), ZN => n102);
   U81 : NOR2_X1 port map( A1 => n103, A2 => n115, ZN => Bls(1));
   U82 : INV_X1 port map( A => B(1), ZN => n103);
   U83 : NOR2_X1 port map( A1 => n104, A2 => n115, ZN => Bls(19));
   U84 : INV_X1 port map( A => B(19), ZN => n104);
   U85 : NOR2_X1 port map( A1 => n105, A2 => n115, ZN => Bls(18));
   U86 : INV_X1 port map( A => B(18), ZN => n105);
   U87 : NOR2_X1 port map( A1 => n106, A2 => n115, ZN => Bls(17));
   U88 : INV_X1 port map( A => B(17), ZN => n106);
   U89 : NOR2_X1 port map( A1 => n107, A2 => n115, ZN => Bls(16));
   U90 : INV_X1 port map( A => B(16), ZN => n107);
   U91 : NOR2_X1 port map( A1 => n108, A2 => n115, ZN => Bls(15));
   U92 : INV_X1 port map( A => B(15), ZN => n108);
   U93 : NOR2_X1 port map( A1 => n109, A2 => n115, ZN => Bls(14));
   U94 : INV_X1 port map( A => B(14), ZN => n109);
   U95 : NOR2_X1 port map( A1 => n110, A2 => n115, ZN => Bls(13));
   U96 : INV_X1 port map( A => B(13), ZN => n110);
   U97 : NOR2_X1 port map( A1 => n111, A2 => n115, ZN => Bls(12));
   U98 : INV_X1 port map( A => B(12), ZN => n111);
   U99 : NOR2_X1 port map( A1 => n112, A2 => n115, ZN => Bls(11));
   U100 : INV_X1 port map( A => B(11), ZN => n112);
   U101 : NOR2_X1 port map( A1 => n113, A2 => n115, ZN => Bls(10));
   U102 : INV_X1 port map( A => B(10), ZN => n113);
   U103 : NOR2_X1 port map( A1 => n114, A2 => n115, ZN => Bls(0));
   U104 : INV_X1 port map( A => B(0), ZN => n114);
   U105 : NOR2_X1 port map( A1 => n82, A2 => n116, ZN => Ap4(9));
   U106 : NOR2_X1 port map( A1 => n82, A2 => n117, ZN => Ap4(8));
   U107 : NOR2_X1 port map( A1 => n82, A2 => n118, ZN => Ap4(7));
   U108 : NOR2_X1 port map( A1 => n82, A2 => n119, ZN => Ap4(6));
   U109 : NOR2_X1 port map( A1 => n82, A2 => n120, ZN => Ap4(5));
   U110 : NOR2_X1 port map( A1 => n82, A2 => n121, ZN => Ap4(4));
   U111 : NOR2_X1 port map( A1 => n82, A2 => n122, ZN => Ap4(3));
   U112 : NOR2_X1 port map( A1 => n82, A2 => n123, ZN => Ap4(31));
   U113 : NOR2_X1 port map( A1 => n82, A2 => n124, ZN => Ap4(30));
   U114 : NOR2_X1 port map( A1 => n82, A2 => n125, ZN => Ap4(2));
   U115 : NOR2_X1 port map( A1 => n82, A2 => n126, ZN => Ap4(29));
   U116 : NOR2_X1 port map( A1 => n82, A2 => n127, ZN => Ap4(28));
   U117 : NOR2_X1 port map( A1 => n82, A2 => n128, ZN => Ap4(27));
   U118 : NOR2_X1 port map( A1 => n82, A2 => n129, ZN => Ap4(26));
   U119 : NOR2_X1 port map( A1 => n82, A2 => n130, ZN => Ap4(25));
   U120 : NOR2_X1 port map( A1 => n82, A2 => n131, ZN => Ap4(24));
   U121 : NOR2_X1 port map( A1 => n82, A2 => n132, ZN => Ap4(23));
   U122 : NOR2_X1 port map( A1 => n82, A2 => n133, ZN => Ap4(22));
   U123 : NOR2_X1 port map( A1 => n82, A2 => n134, ZN => Ap4(21));
   U124 : NOR2_X1 port map( A1 => n82, A2 => n135, ZN => Ap4(20));
   U125 : NOR2_X1 port map( A1 => n82, A2 => n136, ZN => Ap4(1));
   U126 : NOR2_X1 port map( A1 => n82, A2 => n137, ZN => Ap4(19));
   U127 : NOR2_X1 port map( A1 => n82, A2 => n138, ZN => Ap4(18));
   U128 : NOR2_X1 port map( A1 => n82, A2 => n139, ZN => Ap4(17));
   U129 : NOR2_X1 port map( A1 => n82, A2 => n140, ZN => Ap4(16));
   U130 : NOR2_X1 port map( A1 => n82, A2 => n141, ZN => Ap4(15));
   U131 : NOR2_X1 port map( A1 => n82, A2 => n142, ZN => Ap4(14));
   U132 : NOR2_X1 port map( A1 => n82, A2 => n143, ZN => Ap4(13));
   U133 : NOR2_X1 port map( A1 => n82, A2 => n144, ZN => Ap4(12));
   U134 : NOR2_X1 port map( A1 => n82, A2 => n145, ZN => Ap4(11));
   U135 : NOR2_X1 port map( A1 => n82, A2 => n146, ZN => Ap4(10));
   U136 : NOR2_X1 port map( A1 => n82, A2 => n147, ZN => Ap4(0));
   U137 : NAND2_X1 port map( A1 => n148, A2 => n149, ZN => n79);
   U138 : OAI21_X1 port map( B1 => FUNC(0), B2 => n80, A => FUNC(1), ZN => n149
                           );
   U139 : INV_X1 port map( A => FUNC(3), ZN => n80);
   U140 : MUX2_X1 port map( A => FUNC(0), B => FUNC(1), S => FUNC(2), Z => n148
                           );
   U141 : NAND3_X1 port map( A1 => n150, A2 => n151, A3 => FUNC(2), ZN => n81);
   U142 : NOR2_X1 port map( A1 => n115, A2 => n116, ZN => Als(9));
   U143 : INV_X1 port map( A => A(9), ZN => n116);
   U144 : NOR2_X1 port map( A1 => n115, A2 => n117, ZN => Als(8));
   U145 : INV_X1 port map( A => A(8), ZN => n117);
   U146 : NOR2_X1 port map( A1 => n115, A2 => n118, ZN => Als(7));
   U147 : INV_X1 port map( A => A(7), ZN => n118);
   U148 : NOR2_X1 port map( A1 => n115, A2 => n119, ZN => Als(6));
   U149 : INV_X1 port map( A => A(6), ZN => n119);
   U150 : NOR2_X1 port map( A1 => n115, A2 => n120, ZN => Als(5));
   U151 : INV_X1 port map( A => A(5), ZN => n120);
   U152 : NOR2_X1 port map( A1 => n115, A2 => n121, ZN => Als(4));
   U153 : INV_X1 port map( A => A(4), ZN => n121);
   U154 : NOR2_X1 port map( A1 => n115, A2 => n122, ZN => Als(3));
   U155 : INV_X1 port map( A => A(3), ZN => n122);
   U156 : NOR2_X1 port map( A1 => n115, A2 => n123, ZN => Als(31));
   U157 : INV_X1 port map( A => A(31), ZN => n123);
   U158 : NOR2_X1 port map( A1 => n115, A2 => n124, ZN => Als(30));
   U159 : INV_X1 port map( A => A(30), ZN => n124);
   U160 : NOR2_X1 port map( A1 => n115, A2 => n125, ZN => Als(2));
   U161 : INV_X1 port map( A => A(2), ZN => n125);
   U162 : NOR2_X1 port map( A1 => n115, A2 => n126, ZN => Als(29));
   U163 : INV_X1 port map( A => A(29), ZN => n126);
   U164 : NOR2_X1 port map( A1 => n115, A2 => n127, ZN => Als(28));
   U165 : INV_X1 port map( A => A(28), ZN => n127);
   U166 : NOR2_X1 port map( A1 => n115, A2 => n128, ZN => Als(27));
   U167 : INV_X1 port map( A => A(27), ZN => n128);
   U168 : NOR2_X1 port map( A1 => n115, A2 => n129, ZN => Als(26));
   U169 : INV_X1 port map( A => A(26), ZN => n129);
   U170 : NOR2_X1 port map( A1 => n115, A2 => n130, ZN => Als(25));
   U171 : INV_X1 port map( A => A(25), ZN => n130);
   U172 : NOR2_X1 port map( A1 => n115, A2 => n131, ZN => Als(24));
   U173 : INV_X1 port map( A => A(24), ZN => n131);
   U174 : NOR2_X1 port map( A1 => n115, A2 => n132, ZN => Als(23));
   U175 : INV_X1 port map( A => A(23), ZN => n132);
   U176 : NOR2_X1 port map( A1 => n115, A2 => n133, ZN => Als(22));
   U177 : INV_X1 port map( A => A(22), ZN => n133);
   U178 : NOR2_X1 port map( A1 => n115, A2 => n134, ZN => Als(21));
   U179 : INV_X1 port map( A => A(21), ZN => n134);
   U180 : NOR2_X1 port map( A1 => n115, A2 => n135, ZN => Als(20));
   U181 : INV_X1 port map( A => A(20), ZN => n135);
   U182 : NOR2_X1 port map( A1 => n115, A2 => n136, ZN => Als(1));
   U183 : INV_X1 port map( A => A(1), ZN => n136);
   U184 : NOR2_X1 port map( A1 => n115, A2 => n137, ZN => Als(19));
   U185 : INV_X1 port map( A => A(19), ZN => n137);
   U186 : NOR2_X1 port map( A1 => n115, A2 => n138, ZN => Als(18));
   U187 : INV_X1 port map( A => A(18), ZN => n138);
   U188 : NOR2_X1 port map( A1 => n115, A2 => n139, ZN => Als(17));
   U189 : INV_X1 port map( A => A(17), ZN => n139);
   U190 : NOR2_X1 port map( A1 => n115, A2 => n140, ZN => Als(16));
   U191 : INV_X1 port map( A => A(16), ZN => n140);
   U192 : NOR2_X1 port map( A1 => n115, A2 => n141, ZN => Als(15));
   U193 : INV_X1 port map( A => A(15), ZN => n141);
   U194 : NOR2_X1 port map( A1 => n115, A2 => n142, ZN => Als(14));
   U195 : INV_X1 port map( A => A(14), ZN => n142);
   U196 : NOR2_X1 port map( A1 => n115, A2 => n143, ZN => Als(13));
   U197 : INV_X1 port map( A => A(13), ZN => n143);
   U198 : NOR2_X1 port map( A1 => n115, A2 => n144, ZN => Als(12));
   U199 : INV_X1 port map( A => A(12), ZN => n144);
   U200 : NOR2_X1 port map( A1 => n115, A2 => n145, ZN => Als(11));
   U201 : INV_X1 port map( A => A(11), ZN => n145);
   U202 : NOR2_X1 port map( A1 => n115, A2 => n146, ZN => Als(10));
   U203 : INV_X1 port map( A => A(10), ZN => n146);
   U204 : NOR2_X1 port map( A1 => n115, A2 => n147, ZN => Als(0));
   U205 : INV_X1 port map( A => A(0), ZN => n147);
   U206 : OAI21_X1 port map( B1 => FUNC(3), B2 => n150, A => FUNC(2), ZN => 
                           n152);
   U207 : INV_X1 port map( A => FUNC(1), ZN => n150);
   U208 : INV_X1 port map( A => FUNC(0), ZN => n151);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity comparator_bits32 is

   port( Cout, EN : in std_logic;  func : in std_logic_vector (0 to 3);  sum : 
         in std_logic_vector (31 downto 0);  set : out std_logic_vector (31 
         downto 0));

end comparator_bits32;

architecture SYN_BEHAVIORAL of comparator_bits32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, set_0_port, n19, n20, n21, n22, n23, n24, n25, n26, 
      n27, n28, n29, n30, n31, n32, n33, n34, n35, n36 : std_logic;

begin
   set <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, set_0_port 
      );
   
   X_Logic0_port <= '0';
   U2 : AND2_X1 port map( A1 => n19, A2 => EN, ZN => set_0_port);
   U3 : MUX2_X1 port map( A => n20, B => n21, S => func(1), Z => n19);
   U4 : AND4_X1 port map( A1 => n22, A2 => n23, A3 => func(3), A4 => func(2), 
                           ZN => n21);
   U5 : INV_X1 port map( A => n24, ZN => n23);
   U6 : NOR3_X1 port map( A1 => n22, A2 => func(2), A3 => n25, ZN => n20);
   U7 : XOR2_X1 port map( A => n26, B => Cout, Z => n25);
   U8 : OR2_X1 port map( A1 => func(3), A2 => n24, ZN => n26);
   U9 : NOR2_X1 port map( A1 => n27, A2 => n28, ZN => n24);
   U10 : NAND4_X1 port map( A1 => n29, A2 => n30, A3 => n31, A4 => n32, ZN => 
                           n28);
   U11 : NOR4_X1 port map( A1 => sum(23), A2 => sum(22), A3 => sum(21), A4 => 
                           sum(20), ZN => n32);
   U12 : NOR4_X1 port map( A1 => sum(1), A2 => sum(19), A3 => sum(18), A4 => 
                           sum(17), ZN => n31);
   U13 : NOR4_X1 port map( A1 => sum(16), A2 => sum(15), A3 => sum(14), A4 => 
                           sum(13), ZN => n30);
   U14 : NOR4_X1 port map( A1 => sum(12), A2 => sum(11), A3 => sum(10), A4 => 
                           sum(0), ZN => n29);
   U15 : NAND4_X1 port map( A1 => n33, A2 => n34, A3 => n35, A4 => n36, ZN => 
                           n27);
   U16 : NOR4_X1 port map( A1 => sum(9), A2 => sum(8), A3 => sum(7), A4 => 
                           sum(6), ZN => n36);
   U17 : NOR4_X1 port map( A1 => sum(5), A2 => sum(4), A3 => sum(3), A4 => 
                           sum(31), ZN => n35);
   U18 : NOR4_X1 port map( A1 => sum(30), A2 => sum(2), A3 => sum(29), A4 => 
                           sum(28), ZN => n34);
   U19 : NOR4_X1 port map( A1 => sum(27), A2 => sum(26), A3 => sum(25), A4 => 
                           sum(24), ZN => n33);
   U20 : INV_X1 port map( A => func(0), ZN => n22);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity outputSelect_nbits32 is

   port( FUNC : in std_logic_vector (0 to 3);  p4_out, LS_OUT, comp_out : in 
         std_logic_vector (31 downto 0);  outputSel : out std_logic_vector (31 
         downto 0));

end outputSelect_nbits32;

architecture SYN_BEHAVIORAL of outputSelect_nbits32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118 : std_logic;

begin
   
   U2 : INV_X2 port map( A => n112, ZN => n80);
   U3 : AND2_X2 port map( A1 => n118, A2 => n117, ZN => n79);
   U4 : OR3_X1 port map( A1 => FUNC(1), A2 => FUNC(0), A3 => n116, ZN => n78);
   U5 : INV_X2 port map( A => n78, ZN => n76);
   U6 : INV_X1 port map( A => n77, ZN => outputSel(0));
   U7 : AOI222_X1 port map( A1 => p4_out(0), A2 => n76, B1 => LS_OUT(0), B2 => 
                           n79, C1 => comp_out(0), C2 => n80, ZN => n77);
   U8 : INV_X1 port map( A => n81, ZN => outputSel(11));
   U9 : AOI222_X1 port map( A1 => p4_out(11), A2 => n76, B1 => LS_OUT(11), B2 
                           => n79, C1 => comp_out(11), C2 => n80, ZN => n81);
   U10 : INV_X1 port map( A => n82, ZN => outputSel(10));
   U11 : AOI222_X1 port map( A1 => p4_out(10), A2 => n76, B1 => LS_OUT(10), B2 
                           => n79, C1 => comp_out(10), C2 => n80, ZN => n82);
   U12 : INV_X1 port map( A => n83, ZN => outputSel(9));
   U13 : AOI222_X1 port map( A1 => p4_out(9), A2 => n76, B1 => LS_OUT(9), B2 =>
                           n79, C1 => comp_out(9), C2 => n80, ZN => n83);
   U14 : INV_X1 port map( A => n84, ZN => outputSel(8));
   U15 : AOI222_X1 port map( A1 => p4_out(8), A2 => n76, B1 => LS_OUT(8), B2 =>
                           n79, C1 => comp_out(8), C2 => n80, ZN => n84);
   U16 : INV_X1 port map( A => n85, ZN => outputSel(15));
   U17 : AOI222_X1 port map( A1 => p4_out(15), A2 => n76, B1 => LS_OUT(15), B2 
                           => n79, C1 => comp_out(15), C2 => n80, ZN => n85);
   U18 : INV_X1 port map( A => n86, ZN => outputSel(14));
   U19 : AOI222_X1 port map( A1 => p4_out(14), A2 => n76, B1 => LS_OUT(14), B2 
                           => n79, C1 => comp_out(14), C2 => n80, ZN => n86);
   U20 : INV_X1 port map( A => n87, ZN => outputSel(13));
   U21 : AOI222_X1 port map( A1 => p4_out(13), A2 => n76, B1 => LS_OUT(13), B2 
                           => n79, C1 => comp_out(13), C2 => n80, ZN => n87);
   U22 : INV_X1 port map( A => n88, ZN => outputSel(12));
   U23 : AOI222_X1 port map( A1 => p4_out(12), A2 => n76, B1 => LS_OUT(12), B2 
                           => n79, C1 => comp_out(12), C2 => n80, ZN => n88);
   U24 : INV_X1 port map( A => n89, ZN => outputSel(19));
   U25 : AOI222_X1 port map( A1 => p4_out(19), A2 => n76, B1 => LS_OUT(19), B2 
                           => n79, C1 => comp_out(19), C2 => n80, ZN => n89);
   U26 : INV_X1 port map( A => n90, ZN => outputSel(18));
   U27 : AOI222_X1 port map( A1 => p4_out(18), A2 => n76, B1 => LS_OUT(18), B2 
                           => n79, C1 => comp_out(18), C2 => n80, ZN => n90);
   U28 : INV_X1 port map( A => n91, ZN => outputSel(17));
   U29 : AOI222_X1 port map( A1 => p4_out(17), A2 => n76, B1 => LS_OUT(17), B2 
                           => n79, C1 => comp_out(17), C2 => n80, ZN => n91);
   U30 : INV_X1 port map( A => n92, ZN => outputSel(16));
   U31 : AOI222_X1 port map( A1 => p4_out(16), A2 => n76, B1 => LS_OUT(16), B2 
                           => n79, C1 => comp_out(16), C2 => n80, ZN => n92);
   U32 : INV_X1 port map( A => n93, ZN => outputSel(23));
   U33 : AOI222_X1 port map( A1 => p4_out(23), A2 => n76, B1 => LS_OUT(23), B2 
                           => n79, C1 => comp_out(23), C2 => n80, ZN => n93);
   U34 : INV_X1 port map( A => n94, ZN => outputSel(22));
   U35 : AOI222_X1 port map( A1 => p4_out(22), A2 => n76, B1 => LS_OUT(22), B2 
                           => n79, C1 => comp_out(22), C2 => n80, ZN => n94);
   U36 : INV_X1 port map( A => n95, ZN => outputSel(21));
   U37 : AOI222_X1 port map( A1 => p4_out(21), A2 => n76, B1 => LS_OUT(21), B2 
                           => n79, C1 => comp_out(21), C2 => n80, ZN => n95);
   U38 : INV_X1 port map( A => n96, ZN => outputSel(20));
   U39 : AOI222_X1 port map( A1 => p4_out(20), A2 => n76, B1 => LS_OUT(20), B2 
                           => n79, C1 => comp_out(20), C2 => n80, ZN => n96);
   U40 : INV_X1 port map( A => n97, ZN => outputSel(27));
   U41 : AOI222_X1 port map( A1 => p4_out(27), A2 => n76, B1 => LS_OUT(27), B2 
                           => n79, C1 => comp_out(27), C2 => n80, ZN => n97);
   U42 : INV_X1 port map( A => n98, ZN => outputSel(26));
   U43 : AOI222_X1 port map( A1 => p4_out(26), A2 => n76, B1 => LS_OUT(26), B2 
                           => n79, C1 => comp_out(26), C2 => n80, ZN => n98);
   U44 : INV_X1 port map( A => n99, ZN => outputSel(25));
   U45 : AOI222_X1 port map( A1 => p4_out(25), A2 => n76, B1 => LS_OUT(25), B2 
                           => n79, C1 => comp_out(25), C2 => n80, ZN => n99);
   U46 : INV_X1 port map( A => n100, ZN => outputSel(24));
   U47 : AOI222_X1 port map( A1 => p4_out(24), A2 => n76, B1 => LS_OUT(24), B2 
                           => n79, C1 => comp_out(24), C2 => n80, ZN => n100);
   U48 : INV_X1 port map( A => n101, ZN => outputSel(31));
   U49 : AOI222_X1 port map( A1 => p4_out(31), A2 => n76, B1 => LS_OUT(31), B2 
                           => n79, C1 => comp_out(31), C2 => n80, ZN => n101);
   U50 : INV_X1 port map( A => n102, ZN => outputSel(30));
   U51 : AOI222_X1 port map( A1 => p4_out(30), A2 => n76, B1 => LS_OUT(30), B2 
                           => n79, C1 => comp_out(30), C2 => n80, ZN => n102);
   U52 : INV_X1 port map( A => n103, ZN => outputSel(29));
   U53 : AOI222_X1 port map( A1 => p4_out(29), A2 => n76, B1 => LS_OUT(29), B2 
                           => n79, C1 => comp_out(29), C2 => n80, ZN => n103);
   U54 : INV_X1 port map( A => n104, ZN => outputSel(28));
   U55 : AOI222_X1 port map( A1 => p4_out(28), A2 => n76, B1 => LS_OUT(28), B2 
                           => n79, C1 => comp_out(28), C2 => n80, ZN => n104);
   U56 : INV_X1 port map( A => n105, ZN => outputSel(7));
   U57 : AOI222_X1 port map( A1 => p4_out(7), A2 => n76, B1 => LS_OUT(7), B2 =>
                           n79, C1 => comp_out(7), C2 => n80, ZN => n105);
   U58 : INV_X1 port map( A => n106, ZN => outputSel(6));
   U59 : AOI222_X1 port map( A1 => p4_out(6), A2 => n76, B1 => LS_OUT(6), B2 =>
                           n79, C1 => comp_out(6), C2 => n80, ZN => n106);
   U60 : INV_X1 port map( A => n107, ZN => outputSel(5));
   U61 : AOI222_X1 port map( A1 => p4_out(5), A2 => n76, B1 => LS_OUT(5), B2 =>
                           n79, C1 => comp_out(5), C2 => n80, ZN => n107);
   U62 : INV_X1 port map( A => n108, ZN => outputSel(4));
   U63 : AOI222_X1 port map( A1 => p4_out(4), A2 => n76, B1 => LS_OUT(4), B2 =>
                           n79, C1 => comp_out(4), C2 => n80, ZN => n108);
   U64 : INV_X1 port map( A => n109, ZN => outputSel(3));
   U65 : AOI222_X1 port map( A1 => p4_out(3), A2 => n76, B1 => LS_OUT(3), B2 =>
                           n79, C1 => comp_out(3), C2 => n80, ZN => n109);
   U66 : INV_X1 port map( A => n110, ZN => outputSel(2));
   U67 : AOI222_X1 port map( A1 => p4_out(2), A2 => n76, B1 => LS_OUT(2), B2 =>
                           n79, C1 => comp_out(2), C2 => n80, ZN => n110);
   U68 : INV_X1 port map( A => n111, ZN => outputSel(1));
   U69 : AOI222_X1 port map( A1 => p4_out(1), A2 => n76, B1 => LS_OUT(1), B2 =>
                           n79, C1 => comp_out(1), C2 => n80, ZN => n111);
   U70 : MUX2_X1 port map( A => n113, B => n114, S => n115, Z => n112);
   U71 : NAND2_X1 port map( A1 => FUNC(0), A2 => n116, ZN => n114);
   U72 : NAND3_X1 port map( A1 => FUNC(2), A2 => n117, A3 => FUNC(3), ZN => 
                           n113);
   U73 : INV_X1 port map( A => FUNC(0), ZN => n117);
   U74 : OAI21_X1 port map( B1 => FUNC(3), B2 => n115, A => FUNC(2), ZN => n118
                           );
   U75 : INV_X1 port map( A => FUNC(1), ZN => n115);
   U76 : INV_X1 port map( A => FUNC(2), ZN => n116);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21;

architecture SYN_BEHAVIORAL of MUX21 is

   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X2 port map( A => B, B => A, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity XNOR_logic is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR_logic;

architecture SYN_BEHAVIORAL of XNOR_logic is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity alu_nbits32 is

   port( FUNC : in std_logic_vector (0 to 3);  A, B : in std_logic_vector (31 
         downto 0);  OUTALU : out std_logic_vector (31 downto 0));

end alu_nbits32;

architecture SYN_STRUCTURAL of alu_nbits32 is

   component logic_and_shift_N32
      port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4_ADDER_NBITS32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component ctrl_alu_NBITS32
      port( A, B : in std_logic_vector (31 downto 0);  FUNC : in 
            std_logic_vector (0 to 3);  Ap4, Bp4 : out std_logic_vector (31 
            downto 0);  Cin : out std_logic;  Als, Bls : out std_logic_vector 
            (31 downto 0);  enableComp : out std_logic);
   end component;
   
   component comparator_bits32
      port( Cout, EN : in std_logic;  func : in std_logic_vector (0 to 3);  sum
            : in std_logic_vector (31 downto 0);  set : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component outputSelect_nbits32
      port( FUNC : in std_logic_vector (0 to 3);  p4_out, LS_OUT, comp_out : in
            std_logic_vector (31 downto 0);  outputSel : out std_logic_vector 
            (31 downto 0));
   end component;
   
   signal p4_outsig_31_port, p4_outsig_30_port, p4_outsig_29_port, 
      p4_outsig_28_port, p4_outsig_27_port, p4_outsig_26_port, 
      p4_outsig_25_port, p4_outsig_24_port, p4_outsig_23_port, 
      p4_outsig_22_port, p4_outsig_21_port, p4_outsig_20_port, 
      p4_outsig_19_port, p4_outsig_18_port, p4_outsig_17_port, 
      p4_outsig_16_port, p4_outsig_15_port, p4_outsig_14_port, 
      p4_outsig_13_port, p4_outsig_12_port, p4_outsig_11_port, 
      p4_outsig_10_port, p4_outsig_9_port, p4_outsig_8_port, p4_outsig_7_port, 
      p4_outsig_6_port, p4_outsig_5_port, p4_outsig_4_port, p4_outsig_3_port, 
      p4_outsig_2_port, p4_outsig_1_port, p4_outsig_0_port, LS_OUTsig_31_port, 
      LS_OUTsig_30_port, LS_OUTsig_29_port, LS_OUTsig_28_port, 
      LS_OUTsig_27_port, LS_OUTsig_26_port, LS_OUTsig_25_port, 
      LS_OUTsig_24_port, LS_OUTsig_23_port, LS_OUTsig_22_port, 
      LS_OUTsig_21_port, LS_OUTsig_20_port, LS_OUTsig_19_port, 
      LS_OUTsig_18_port, LS_OUTsig_17_port, LS_OUTsig_16_port, 
      LS_OUTsig_15_port, LS_OUTsig_14_port, LS_OUTsig_13_port, 
      LS_OUTsig_12_port, LS_OUTsig_11_port, LS_OUTsig_10_port, LS_OUTsig_9_port
      , LS_OUTsig_8_port, LS_OUTsig_7_port, LS_OUTsig_6_port, LS_OUTsig_5_port,
      LS_OUTsig_4_port, LS_OUTsig_3_port, LS_OUTsig_2_port, LS_OUTsig_1_port, 
      LS_OUTsig_0_port, comp_outsig_31_port, comp_outsig_30_port, 
      comp_outsig_29_port, comp_outsig_28_port, comp_outsig_27_port, 
      comp_outsig_26_port, comp_outsig_25_port, comp_outsig_24_port, 
      comp_outsig_23_port, comp_outsig_22_port, comp_outsig_21_port, 
      comp_outsig_20_port, comp_outsig_19_port, comp_outsig_18_port, 
      comp_outsig_17_port, comp_outsig_16_port, comp_outsig_15_port, 
      comp_outsig_14_port, comp_outsig_13_port, comp_outsig_12_port, 
      comp_outsig_11_port, comp_outsig_10_port, comp_outsig_9_port, 
      comp_outsig_8_port, comp_outsig_7_port, comp_outsig_6_port, 
      comp_outsig_5_port, comp_outsig_4_port, comp_outsig_3_port, 
      comp_outsig_2_port, comp_outsig_1_port, comp_outsig_0_port, p4_comp_Co, 
      enable_Comp, p4_ctrl_A_31_port, p4_ctrl_A_30_port, p4_ctrl_A_29_port, 
      p4_ctrl_A_28_port, p4_ctrl_A_27_port, p4_ctrl_A_26_port, 
      p4_ctrl_A_25_port, p4_ctrl_A_24_port, p4_ctrl_A_23_port, 
      p4_ctrl_A_22_port, p4_ctrl_A_21_port, p4_ctrl_A_20_port, 
      p4_ctrl_A_19_port, p4_ctrl_A_18_port, p4_ctrl_A_17_port, 
      p4_ctrl_A_16_port, p4_ctrl_A_15_port, p4_ctrl_A_14_port, 
      p4_ctrl_A_13_port, p4_ctrl_A_12_port, p4_ctrl_A_11_port, 
      p4_ctrl_A_10_port, p4_ctrl_A_9_port, p4_ctrl_A_8_port, p4_ctrl_A_7_port, 
      p4_ctrl_A_6_port, p4_ctrl_A_5_port, p4_ctrl_A_4_port, p4_ctrl_A_3_port, 
      p4_ctrl_A_2_port, p4_ctrl_A_1_port, p4_ctrl_A_0_port, p4_ctrl_B_31_port, 
      p4_ctrl_B_30_port, p4_ctrl_B_29_port, p4_ctrl_B_28_port, 
      p4_ctrl_B_27_port, p4_ctrl_B_26_port, p4_ctrl_B_25_port, 
      p4_ctrl_B_24_port, p4_ctrl_B_23_port, p4_ctrl_B_22_port, 
      p4_ctrl_B_21_port, p4_ctrl_B_20_port, p4_ctrl_B_19_port, 
      p4_ctrl_B_18_port, p4_ctrl_B_17_port, p4_ctrl_B_16_port, 
      p4_ctrl_B_15_port, p4_ctrl_B_14_port, p4_ctrl_B_13_port, 
      p4_ctrl_B_12_port, p4_ctrl_B_11_port, p4_ctrl_B_10_port, p4_ctrl_B_9_port
      , p4_ctrl_B_8_port, p4_ctrl_B_7_port, p4_ctrl_B_6_port, p4_ctrl_B_5_port,
      p4_ctrl_B_4_port, p4_ctrl_B_3_port, p4_ctrl_B_2_port, p4_ctrl_B_1_port, 
      p4_ctrl_B_0_port, p4_ctrl_Cin, ctrl_LS_A_31_port, ctrl_LS_A_30_port, 
      ctrl_LS_A_29_port, ctrl_LS_A_28_port, ctrl_LS_A_27_port, 
      ctrl_LS_A_26_port, ctrl_LS_A_25_port, ctrl_LS_A_24_port, 
      ctrl_LS_A_23_port, ctrl_LS_A_22_port, ctrl_LS_A_21_port, 
      ctrl_LS_A_20_port, ctrl_LS_A_19_port, ctrl_LS_A_18_port, 
      ctrl_LS_A_17_port, ctrl_LS_A_16_port, ctrl_LS_A_15_port, 
      ctrl_LS_A_14_port, ctrl_LS_A_13_port, ctrl_LS_A_12_port, 
      ctrl_LS_A_11_port, ctrl_LS_A_10_port, ctrl_LS_A_9_port, ctrl_LS_A_8_port,
      ctrl_LS_A_7_port, ctrl_LS_A_6_port, ctrl_LS_A_5_port, ctrl_LS_A_4_port, 
      ctrl_LS_A_3_port, ctrl_LS_A_2_port, ctrl_LS_A_1_port, ctrl_LS_A_0_port, 
      ctrl_LS_B_31_port, ctrl_LS_B_30_port, ctrl_LS_B_29_port, 
      ctrl_LS_B_28_port, ctrl_LS_B_27_port, ctrl_LS_B_26_port, 
      ctrl_LS_B_25_port, ctrl_LS_B_24_port, ctrl_LS_B_23_port, 
      ctrl_LS_B_22_port, ctrl_LS_B_21_port, ctrl_LS_B_20_port, 
      ctrl_LS_B_19_port, ctrl_LS_B_18_port, ctrl_LS_B_17_port, 
      ctrl_LS_B_16_port, ctrl_LS_B_15_port, ctrl_LS_B_14_port, 
      ctrl_LS_B_13_port, ctrl_LS_B_12_port, ctrl_LS_B_11_port, 
      ctrl_LS_B_10_port, ctrl_LS_B_9_port, ctrl_LS_B_8_port, ctrl_LS_B_7_port, 
      ctrl_LS_B_6_port, ctrl_LS_B_5_port, ctrl_LS_B_4_port, ctrl_LS_B_3_port, 
      ctrl_LS_B_2_port, ctrl_LS_B_1_port, ctrl_LS_B_0_port, n_1373, n_1374, 
      n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, 
      n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, 
      n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, 
      n_1402, n_1403 : std_logic;

begin
   
   comp_outsig_1_port <= '0';
   comp_outsig_2_port <= '0';
   comp_outsig_3_port <= '0';
   comp_outsig_4_port <= '0';
   comp_outsig_5_port <= '0';
   comp_outsig_6_port <= '0';
   comp_outsig_7_port <= '0';
   comp_outsig_8_port <= '0';
   comp_outsig_9_port <= '0';
   comp_outsig_10_port <= '0';
   comp_outsig_11_port <= '0';
   comp_outsig_12_port <= '0';
   comp_outsig_13_port <= '0';
   comp_outsig_14_port <= '0';
   comp_outsig_15_port <= '0';
   comp_outsig_16_port <= '0';
   comp_outsig_17_port <= '0';
   comp_outsig_18_port <= '0';
   comp_outsig_19_port <= '0';
   comp_outsig_20_port <= '0';
   comp_outsig_21_port <= '0';
   comp_outsig_22_port <= '0';
   comp_outsig_23_port <= '0';
   comp_outsig_24_port <= '0';
   comp_outsig_25_port <= '0';
   comp_outsig_26_port <= '0';
   comp_outsig_27_port <= '0';
   comp_outsig_28_port <= '0';
   comp_outsig_29_port <= '0';
   comp_outsig_30_port <= '0';
   comp_outsig_31_port <= '0';
   SELOUT : outputSelect_nbits32 port map( FUNC(0) => FUNC(0), FUNC(1) => 
                           FUNC(1), FUNC(2) => FUNC(2), FUNC(3) => FUNC(3), 
                           p4_out(31) => p4_outsig_31_port, p4_out(30) => 
                           p4_outsig_30_port, p4_out(29) => p4_outsig_29_port, 
                           p4_out(28) => p4_outsig_28_port, p4_out(27) => 
                           p4_outsig_27_port, p4_out(26) => p4_outsig_26_port, 
                           p4_out(25) => p4_outsig_25_port, p4_out(24) => 
                           p4_outsig_24_port, p4_out(23) => p4_outsig_23_port, 
                           p4_out(22) => p4_outsig_22_port, p4_out(21) => 
                           p4_outsig_21_port, p4_out(20) => p4_outsig_20_port, 
                           p4_out(19) => p4_outsig_19_port, p4_out(18) => 
                           p4_outsig_18_port, p4_out(17) => p4_outsig_17_port, 
                           p4_out(16) => p4_outsig_16_port, p4_out(15) => 
                           p4_outsig_15_port, p4_out(14) => p4_outsig_14_port, 
                           p4_out(13) => p4_outsig_13_port, p4_out(12) => 
                           p4_outsig_12_port, p4_out(11) => p4_outsig_11_port, 
                           p4_out(10) => p4_outsig_10_port, p4_out(9) => 
                           p4_outsig_9_port, p4_out(8) => p4_outsig_8_port, 
                           p4_out(7) => p4_outsig_7_port, p4_out(6) => 
                           p4_outsig_6_port, p4_out(5) => p4_outsig_5_port, 
                           p4_out(4) => p4_outsig_4_port, p4_out(3) => 
                           p4_outsig_3_port, p4_out(2) => p4_outsig_2_port, 
                           p4_out(1) => p4_outsig_1_port, p4_out(0) => 
                           p4_outsig_0_port, LS_OUT(31) => LS_OUTsig_31_port, 
                           LS_OUT(30) => LS_OUTsig_30_port, LS_OUT(29) => 
                           LS_OUTsig_29_port, LS_OUT(28) => LS_OUTsig_28_port, 
                           LS_OUT(27) => LS_OUTsig_27_port, LS_OUT(26) => 
                           LS_OUTsig_26_port, LS_OUT(25) => LS_OUTsig_25_port, 
                           LS_OUT(24) => LS_OUTsig_24_port, LS_OUT(23) => 
                           LS_OUTsig_23_port, LS_OUT(22) => LS_OUTsig_22_port, 
                           LS_OUT(21) => LS_OUTsig_21_port, LS_OUT(20) => 
                           LS_OUTsig_20_port, LS_OUT(19) => LS_OUTsig_19_port, 
                           LS_OUT(18) => LS_OUTsig_18_port, LS_OUT(17) => 
                           LS_OUTsig_17_port, LS_OUT(16) => LS_OUTsig_16_port, 
                           LS_OUT(15) => LS_OUTsig_15_port, LS_OUT(14) => 
                           LS_OUTsig_14_port, LS_OUT(13) => LS_OUTsig_13_port, 
                           LS_OUT(12) => LS_OUTsig_12_port, LS_OUT(11) => 
                           LS_OUTsig_11_port, LS_OUT(10) => LS_OUTsig_10_port, 
                           LS_OUT(9) => LS_OUTsig_9_port, LS_OUT(8) => 
                           LS_OUTsig_8_port, LS_OUT(7) => LS_OUTsig_7_port, 
                           LS_OUT(6) => LS_OUTsig_6_port, LS_OUT(5) => 
                           LS_OUTsig_5_port, LS_OUT(4) => LS_OUTsig_4_port, 
                           LS_OUT(3) => LS_OUTsig_3_port, LS_OUT(2) => 
                           LS_OUTsig_2_port, LS_OUT(1) => LS_OUTsig_1_port, 
                           LS_OUT(0) => LS_OUTsig_0_port, comp_out(31) => 
                           comp_outsig_31_port, comp_out(30) => 
                           comp_outsig_30_port, comp_out(29) => 
                           comp_outsig_29_port, comp_out(28) => 
                           comp_outsig_28_port, comp_out(27) => 
                           comp_outsig_27_port, comp_out(26) => 
                           comp_outsig_26_port, comp_out(25) => 
                           comp_outsig_25_port, comp_out(24) => 
                           comp_outsig_24_port, comp_out(23) => 
                           comp_outsig_23_port, comp_out(22) => 
                           comp_outsig_22_port, comp_out(21) => 
                           comp_outsig_21_port, comp_out(20) => 
                           comp_outsig_20_port, comp_out(19) => 
                           comp_outsig_19_port, comp_out(18) => 
                           comp_outsig_18_port, comp_out(17) => 
                           comp_outsig_17_port, comp_out(16) => 
                           comp_outsig_16_port, comp_out(15) => 
                           comp_outsig_15_port, comp_out(14) => 
                           comp_outsig_14_port, comp_out(13) => 
                           comp_outsig_13_port, comp_out(12) => 
                           comp_outsig_12_port, comp_out(11) => 
                           comp_outsig_11_port, comp_out(10) => 
                           comp_outsig_10_port, comp_out(9) => 
                           comp_outsig_9_port, comp_out(8) => 
                           comp_outsig_8_port, comp_out(7) => 
                           comp_outsig_7_port, comp_out(6) => 
                           comp_outsig_6_port, comp_out(5) => 
                           comp_outsig_5_port, comp_out(4) => 
                           comp_outsig_4_port, comp_out(3) => 
                           comp_outsig_3_port, comp_out(2) => 
                           comp_outsig_2_port, comp_out(1) => 
                           comp_outsig_1_port, comp_out(0) => 
                           comp_outsig_0_port, outputSel(31) => OUTALU(31), 
                           outputSel(30) => OUTALU(30), outputSel(29) => 
                           OUTALU(29), outputSel(28) => OUTALU(28), 
                           outputSel(27) => OUTALU(27), outputSel(26) => 
                           OUTALU(26), outputSel(25) => OUTALU(25), 
                           outputSel(24) => OUTALU(24), outputSel(23) => 
                           OUTALU(23), outputSel(22) => OUTALU(22), 
                           outputSel(21) => OUTALU(21), outputSel(20) => 
                           OUTALU(20), outputSel(19) => OUTALU(19), 
                           outputSel(18) => OUTALU(18), outputSel(17) => 
                           OUTALU(17), outputSel(16) => OUTALU(16), 
                           outputSel(15) => OUTALU(15), outputSel(14) => 
                           OUTALU(14), outputSel(13) => OUTALU(13), 
                           outputSel(12) => OUTALU(12), outputSel(11) => 
                           OUTALU(11), outputSel(10) => OUTALU(10), 
                           outputSel(9) => OUTALU(9), outputSel(8) => OUTALU(8)
                           , outputSel(7) => OUTALU(7), outputSel(6) => 
                           OUTALU(6), outputSel(5) => OUTALU(5), outputSel(4) 
                           => OUTALU(4), outputSel(3) => OUTALU(3), 
                           outputSel(2) => OUTALU(2), outputSel(1) => OUTALU(1)
                           , outputSel(0) => OUTALU(0));
   COMP : comparator_bits32 port map( Cout => p4_comp_Co, EN => enable_Comp, 
                           func(0) => FUNC(0), func(1) => FUNC(1), func(2) => 
                           FUNC(2), func(3) => FUNC(3), sum(31) => 
                           p4_outsig_31_port, sum(30) => p4_outsig_30_port, 
                           sum(29) => p4_outsig_29_port, sum(28) => 
                           p4_outsig_28_port, sum(27) => p4_outsig_27_port, 
                           sum(26) => p4_outsig_26_port, sum(25) => 
                           p4_outsig_25_port, sum(24) => p4_outsig_24_port, 
                           sum(23) => p4_outsig_23_port, sum(22) => 
                           p4_outsig_22_port, sum(21) => p4_outsig_21_port, 
                           sum(20) => p4_outsig_20_port, sum(19) => 
                           p4_outsig_19_port, sum(18) => p4_outsig_18_port, 
                           sum(17) => p4_outsig_17_port, sum(16) => 
                           p4_outsig_16_port, sum(15) => p4_outsig_15_port, 
                           sum(14) => p4_outsig_14_port, sum(13) => 
                           p4_outsig_13_port, sum(12) => p4_outsig_12_port, 
                           sum(11) => p4_outsig_11_port, sum(10) => 
                           p4_outsig_10_port, sum(9) => p4_outsig_9_port, 
                           sum(8) => p4_outsig_8_port, sum(7) => 
                           p4_outsig_7_port, sum(6) => p4_outsig_6_port, sum(5)
                           => p4_outsig_5_port, sum(4) => p4_outsig_4_port, 
                           sum(3) => p4_outsig_3_port, sum(2) => 
                           p4_outsig_2_port, sum(1) => p4_outsig_1_port, sum(0)
                           => p4_outsig_0_port, set(31) => n_1373, set(30) => 
                           n_1374, set(29) => n_1375, set(28) => n_1376, 
                           set(27) => n_1377, set(26) => n_1378, set(25) => 
                           n_1379, set(24) => n_1380, set(23) => n_1381, 
                           set(22) => n_1382, set(21) => n_1383, set(20) => 
                           n_1384, set(19) => n_1385, set(18) => n_1386, 
                           set(17) => n_1387, set(16) => n_1388, set(15) => 
                           n_1389, set(14) => n_1390, set(13) => n_1391, 
                           set(12) => n_1392, set(11) => n_1393, set(10) => 
                           n_1394, set(9) => n_1395, set(8) => n_1396, set(7) 
                           => n_1397, set(6) => n_1398, set(5) => n_1399, 
                           set(4) => n_1400, set(3) => n_1401, set(2) => n_1402
                           , set(1) => n_1403, set(0) => comp_outsig_0_port);
   CTRLALU : ctrl_alu_NBITS32 port map( A(31) => A(31), A(30) => A(30), A(29) 
                           => A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), FUNC(0) => FUNC(0), FUNC(1) => FUNC(1), 
                           FUNC(2) => FUNC(2), FUNC(3) => FUNC(3), Ap4(31) => 
                           p4_ctrl_A_31_port, Ap4(30) => p4_ctrl_A_30_port, 
                           Ap4(29) => p4_ctrl_A_29_port, Ap4(28) => 
                           p4_ctrl_A_28_port, Ap4(27) => p4_ctrl_A_27_port, 
                           Ap4(26) => p4_ctrl_A_26_port, Ap4(25) => 
                           p4_ctrl_A_25_port, Ap4(24) => p4_ctrl_A_24_port, 
                           Ap4(23) => p4_ctrl_A_23_port, Ap4(22) => 
                           p4_ctrl_A_22_port, Ap4(21) => p4_ctrl_A_21_port, 
                           Ap4(20) => p4_ctrl_A_20_port, Ap4(19) => 
                           p4_ctrl_A_19_port, Ap4(18) => p4_ctrl_A_18_port, 
                           Ap4(17) => p4_ctrl_A_17_port, Ap4(16) => 
                           p4_ctrl_A_16_port, Ap4(15) => p4_ctrl_A_15_port, 
                           Ap4(14) => p4_ctrl_A_14_port, Ap4(13) => 
                           p4_ctrl_A_13_port, Ap4(12) => p4_ctrl_A_12_port, 
                           Ap4(11) => p4_ctrl_A_11_port, Ap4(10) => 
                           p4_ctrl_A_10_port, Ap4(9) => p4_ctrl_A_9_port, 
                           Ap4(8) => p4_ctrl_A_8_port, Ap4(7) => 
                           p4_ctrl_A_7_port, Ap4(6) => p4_ctrl_A_6_port, Ap4(5)
                           => p4_ctrl_A_5_port, Ap4(4) => p4_ctrl_A_4_port, 
                           Ap4(3) => p4_ctrl_A_3_port, Ap4(2) => 
                           p4_ctrl_A_2_port, Ap4(1) => p4_ctrl_A_1_port, Ap4(0)
                           => p4_ctrl_A_0_port, Bp4(31) => p4_ctrl_B_31_port, 
                           Bp4(30) => p4_ctrl_B_30_port, Bp4(29) => 
                           p4_ctrl_B_29_port, Bp4(28) => p4_ctrl_B_28_port, 
                           Bp4(27) => p4_ctrl_B_27_port, Bp4(26) => 
                           p4_ctrl_B_26_port, Bp4(25) => p4_ctrl_B_25_port, 
                           Bp4(24) => p4_ctrl_B_24_port, Bp4(23) => 
                           p4_ctrl_B_23_port, Bp4(22) => p4_ctrl_B_22_port, 
                           Bp4(21) => p4_ctrl_B_21_port, Bp4(20) => 
                           p4_ctrl_B_20_port, Bp4(19) => p4_ctrl_B_19_port, 
                           Bp4(18) => p4_ctrl_B_18_port, Bp4(17) => 
                           p4_ctrl_B_17_port, Bp4(16) => p4_ctrl_B_16_port, 
                           Bp4(15) => p4_ctrl_B_15_port, Bp4(14) => 
                           p4_ctrl_B_14_port, Bp4(13) => p4_ctrl_B_13_port, 
                           Bp4(12) => p4_ctrl_B_12_port, Bp4(11) => 
                           p4_ctrl_B_11_port, Bp4(10) => p4_ctrl_B_10_port, 
                           Bp4(9) => p4_ctrl_B_9_port, Bp4(8) => 
                           p4_ctrl_B_8_port, Bp4(7) => p4_ctrl_B_7_port, Bp4(6)
                           => p4_ctrl_B_6_port, Bp4(5) => p4_ctrl_B_5_port, 
                           Bp4(4) => p4_ctrl_B_4_port, Bp4(3) => 
                           p4_ctrl_B_3_port, Bp4(2) => p4_ctrl_B_2_port, Bp4(1)
                           => p4_ctrl_B_1_port, Bp4(0) => p4_ctrl_B_0_port, Cin
                           => p4_ctrl_Cin, Als(31) => ctrl_LS_A_31_port, 
                           Als(30) => ctrl_LS_A_30_port, Als(29) => 
                           ctrl_LS_A_29_port, Als(28) => ctrl_LS_A_28_port, 
                           Als(27) => ctrl_LS_A_27_port, Als(26) => 
                           ctrl_LS_A_26_port, Als(25) => ctrl_LS_A_25_port, 
                           Als(24) => ctrl_LS_A_24_port, Als(23) => 
                           ctrl_LS_A_23_port, Als(22) => ctrl_LS_A_22_port, 
                           Als(21) => ctrl_LS_A_21_port, Als(20) => 
                           ctrl_LS_A_20_port, Als(19) => ctrl_LS_A_19_port, 
                           Als(18) => ctrl_LS_A_18_port, Als(17) => 
                           ctrl_LS_A_17_port, Als(16) => ctrl_LS_A_16_port, 
                           Als(15) => ctrl_LS_A_15_port, Als(14) => 
                           ctrl_LS_A_14_port, Als(13) => ctrl_LS_A_13_port, 
                           Als(12) => ctrl_LS_A_12_port, Als(11) => 
                           ctrl_LS_A_11_port, Als(10) => ctrl_LS_A_10_port, 
                           Als(9) => ctrl_LS_A_9_port, Als(8) => 
                           ctrl_LS_A_8_port, Als(7) => ctrl_LS_A_7_port, Als(6)
                           => ctrl_LS_A_6_port, Als(5) => ctrl_LS_A_5_port, 
                           Als(4) => ctrl_LS_A_4_port, Als(3) => 
                           ctrl_LS_A_3_port, Als(2) => ctrl_LS_A_2_port, Als(1)
                           => ctrl_LS_A_1_port, Als(0) => ctrl_LS_A_0_port, 
                           Bls(31) => ctrl_LS_B_31_port, Bls(30) => 
                           ctrl_LS_B_30_port, Bls(29) => ctrl_LS_B_29_port, 
                           Bls(28) => ctrl_LS_B_28_port, Bls(27) => 
                           ctrl_LS_B_27_port, Bls(26) => ctrl_LS_B_26_port, 
                           Bls(25) => ctrl_LS_B_25_port, Bls(24) => 
                           ctrl_LS_B_24_port, Bls(23) => ctrl_LS_B_23_port, 
                           Bls(22) => ctrl_LS_B_22_port, Bls(21) => 
                           ctrl_LS_B_21_port, Bls(20) => ctrl_LS_B_20_port, 
                           Bls(19) => ctrl_LS_B_19_port, Bls(18) => 
                           ctrl_LS_B_18_port, Bls(17) => ctrl_LS_B_17_port, 
                           Bls(16) => ctrl_LS_B_16_port, Bls(15) => 
                           ctrl_LS_B_15_port, Bls(14) => ctrl_LS_B_14_port, 
                           Bls(13) => ctrl_LS_B_13_port, Bls(12) => 
                           ctrl_LS_B_12_port, Bls(11) => ctrl_LS_B_11_port, 
                           Bls(10) => ctrl_LS_B_10_port, Bls(9) => 
                           ctrl_LS_B_9_port, Bls(8) => ctrl_LS_B_8_port, Bls(7)
                           => ctrl_LS_B_7_port, Bls(6) => ctrl_LS_B_6_port, 
                           Bls(5) => ctrl_LS_B_5_port, Bls(4) => 
                           ctrl_LS_B_4_port, Bls(3) => ctrl_LS_B_3_port, Bls(2)
                           => ctrl_LS_B_2_port, Bls(1) => ctrl_LS_B_1_port, 
                           Bls(0) => ctrl_LS_B_0_port, enableComp => 
                           enable_Comp);
   ADDER_SUB : P4_ADDER_NBITS32 port map( A(31) => p4_ctrl_A_31_port, A(30) => 
                           p4_ctrl_A_30_port, A(29) => p4_ctrl_A_29_port, A(28)
                           => p4_ctrl_A_28_port, A(27) => p4_ctrl_A_27_port, 
                           A(26) => p4_ctrl_A_26_port, A(25) => 
                           p4_ctrl_A_25_port, A(24) => p4_ctrl_A_24_port, A(23)
                           => p4_ctrl_A_23_port, A(22) => p4_ctrl_A_22_port, 
                           A(21) => p4_ctrl_A_21_port, A(20) => 
                           p4_ctrl_A_20_port, A(19) => p4_ctrl_A_19_port, A(18)
                           => p4_ctrl_A_18_port, A(17) => p4_ctrl_A_17_port, 
                           A(16) => p4_ctrl_A_16_port, A(15) => 
                           p4_ctrl_A_15_port, A(14) => p4_ctrl_A_14_port, A(13)
                           => p4_ctrl_A_13_port, A(12) => p4_ctrl_A_12_port, 
                           A(11) => p4_ctrl_A_11_port, A(10) => 
                           p4_ctrl_A_10_port, A(9) => p4_ctrl_A_9_port, A(8) =>
                           p4_ctrl_A_8_port, A(7) => p4_ctrl_A_7_port, A(6) => 
                           p4_ctrl_A_6_port, A(5) => p4_ctrl_A_5_port, A(4) => 
                           p4_ctrl_A_4_port, A(3) => p4_ctrl_A_3_port, A(2) => 
                           p4_ctrl_A_2_port, A(1) => p4_ctrl_A_1_port, A(0) => 
                           p4_ctrl_A_0_port, B(31) => p4_ctrl_B_31_port, B(30) 
                           => p4_ctrl_B_30_port, B(29) => p4_ctrl_B_29_port, 
                           B(28) => p4_ctrl_B_28_port, B(27) => 
                           p4_ctrl_B_27_port, B(26) => p4_ctrl_B_26_port, B(25)
                           => p4_ctrl_B_25_port, B(24) => p4_ctrl_B_24_port, 
                           B(23) => p4_ctrl_B_23_port, B(22) => 
                           p4_ctrl_B_22_port, B(21) => p4_ctrl_B_21_port, B(20)
                           => p4_ctrl_B_20_port, B(19) => p4_ctrl_B_19_port, 
                           B(18) => p4_ctrl_B_18_port, B(17) => 
                           p4_ctrl_B_17_port, B(16) => p4_ctrl_B_16_port, B(15)
                           => p4_ctrl_B_15_port, B(14) => p4_ctrl_B_14_port, 
                           B(13) => p4_ctrl_B_13_port, B(12) => 
                           p4_ctrl_B_12_port, B(11) => p4_ctrl_B_11_port, B(10)
                           => p4_ctrl_B_10_port, B(9) => p4_ctrl_B_9_port, B(8)
                           => p4_ctrl_B_8_port, B(7) => p4_ctrl_B_7_port, B(6) 
                           => p4_ctrl_B_6_port, B(5) => p4_ctrl_B_5_port, B(4) 
                           => p4_ctrl_B_4_port, B(3) => p4_ctrl_B_3_port, B(2) 
                           => p4_ctrl_B_2_port, B(1) => p4_ctrl_B_1_port, B(0) 
                           => p4_ctrl_B_0_port, Ci => p4_ctrl_Cin, S(31) => 
                           p4_outsig_31_port, S(30) => p4_outsig_30_port, S(29)
                           => p4_outsig_29_port, S(28) => p4_outsig_28_port, 
                           S(27) => p4_outsig_27_port, S(26) => 
                           p4_outsig_26_port, S(25) => p4_outsig_25_port, S(24)
                           => p4_outsig_24_port, S(23) => p4_outsig_23_port, 
                           S(22) => p4_outsig_22_port, S(21) => 
                           p4_outsig_21_port, S(20) => p4_outsig_20_port, S(19)
                           => p4_outsig_19_port, S(18) => p4_outsig_18_port, 
                           S(17) => p4_outsig_17_port, S(16) => 
                           p4_outsig_16_port, S(15) => p4_outsig_15_port, S(14)
                           => p4_outsig_14_port, S(13) => p4_outsig_13_port, 
                           S(12) => p4_outsig_12_port, S(11) => 
                           p4_outsig_11_port, S(10) => p4_outsig_10_port, S(9) 
                           => p4_outsig_9_port, S(8) => p4_outsig_8_port, S(7) 
                           => p4_outsig_7_port, S(6) => p4_outsig_6_port, S(5) 
                           => p4_outsig_5_port, S(4) => p4_outsig_4_port, S(3) 
                           => p4_outsig_3_port, S(2) => p4_outsig_2_port, S(1) 
                           => p4_outsig_1_port, S(0) => p4_outsig_0_port, Co =>
                           p4_comp_Co);
   LOGIC_SHIFT : logic_and_shift_N32 port map( FUNC(0) => FUNC(0), FUNC(1) => 
                           FUNC(1), FUNC(2) => FUNC(2), FUNC(3) => FUNC(3), 
                           DATA1(31) => ctrl_LS_A_31_port, DATA1(30) => 
                           ctrl_LS_A_30_port, DATA1(29) => ctrl_LS_A_29_port, 
                           DATA1(28) => ctrl_LS_A_28_port, DATA1(27) => 
                           ctrl_LS_A_27_port, DATA1(26) => ctrl_LS_A_26_port, 
                           DATA1(25) => ctrl_LS_A_25_port, DATA1(24) => 
                           ctrl_LS_A_24_port, DATA1(23) => ctrl_LS_A_23_port, 
                           DATA1(22) => ctrl_LS_A_22_port, DATA1(21) => 
                           ctrl_LS_A_21_port, DATA1(20) => ctrl_LS_A_20_port, 
                           DATA1(19) => ctrl_LS_A_19_port, DATA1(18) => 
                           ctrl_LS_A_18_port, DATA1(17) => ctrl_LS_A_17_port, 
                           DATA1(16) => ctrl_LS_A_16_port, DATA1(15) => 
                           ctrl_LS_A_15_port, DATA1(14) => ctrl_LS_A_14_port, 
                           DATA1(13) => ctrl_LS_A_13_port, DATA1(12) => 
                           ctrl_LS_A_12_port, DATA1(11) => ctrl_LS_A_11_port, 
                           DATA1(10) => ctrl_LS_A_10_port, DATA1(9) => 
                           ctrl_LS_A_9_port, DATA1(8) => ctrl_LS_A_8_port, 
                           DATA1(7) => ctrl_LS_A_7_port, DATA1(6) => 
                           ctrl_LS_A_6_port, DATA1(5) => ctrl_LS_A_5_port, 
                           DATA1(4) => ctrl_LS_A_4_port, DATA1(3) => 
                           ctrl_LS_A_3_port, DATA1(2) => ctrl_LS_A_2_port, 
                           DATA1(1) => ctrl_LS_A_1_port, DATA1(0) => 
                           ctrl_LS_A_0_port, DATA2(31) => ctrl_LS_B_31_port, 
                           DATA2(30) => ctrl_LS_B_30_port, DATA2(29) => 
                           ctrl_LS_B_29_port, DATA2(28) => ctrl_LS_B_28_port, 
                           DATA2(27) => ctrl_LS_B_27_port, DATA2(26) => 
                           ctrl_LS_B_26_port, DATA2(25) => ctrl_LS_B_25_port, 
                           DATA2(24) => ctrl_LS_B_24_port, DATA2(23) => 
                           ctrl_LS_B_23_port, DATA2(22) => ctrl_LS_B_22_port, 
                           DATA2(21) => ctrl_LS_B_21_port, DATA2(20) => 
                           ctrl_LS_B_20_port, DATA2(19) => ctrl_LS_B_19_port, 
                           DATA2(18) => ctrl_LS_B_18_port, DATA2(17) => 
                           ctrl_LS_B_17_port, DATA2(16) => ctrl_LS_B_16_port, 
                           DATA2(15) => ctrl_LS_B_15_port, DATA2(14) => 
                           ctrl_LS_B_14_port, DATA2(13) => ctrl_LS_B_13_port, 
                           DATA2(12) => ctrl_LS_B_12_port, DATA2(11) => 
                           ctrl_LS_B_11_port, DATA2(10) => ctrl_LS_B_10_port, 
                           DATA2(9) => ctrl_LS_B_9_port, DATA2(8) => 
                           ctrl_LS_B_8_port, DATA2(7) => ctrl_LS_B_7_port, 
                           DATA2(6) => ctrl_LS_B_6_port, DATA2(5) => 
                           ctrl_LS_B_5_port, DATA2(4) => ctrl_LS_B_4_port, 
                           DATA2(3) => ctrl_LS_B_3_port, DATA2(2) => 
                           ctrl_LS_B_2_port, DATA2(1) => ctrl_LS_B_1_port, 
                           DATA2(0) => ctrl_LS_B_0_port, OUTALU(31) => 
                           LS_OUTsig_31_port, OUTALU(30) => LS_OUTsig_30_port, 
                           OUTALU(29) => LS_OUTsig_29_port, OUTALU(28) => 
                           LS_OUTsig_28_port, OUTALU(27) => LS_OUTsig_27_port, 
                           OUTALU(26) => LS_OUTsig_26_port, OUTALU(25) => 
                           LS_OUTsig_25_port, OUTALU(24) => LS_OUTsig_24_port, 
                           OUTALU(23) => LS_OUTsig_23_port, OUTALU(22) => 
                           LS_OUTsig_22_port, OUTALU(21) => LS_OUTsig_21_port, 
                           OUTALU(20) => LS_OUTsig_20_port, OUTALU(19) => 
                           LS_OUTsig_19_port, OUTALU(18) => LS_OUTsig_18_port, 
                           OUTALU(17) => LS_OUTsig_17_port, OUTALU(16) => 
                           LS_OUTsig_16_port, OUTALU(15) => LS_OUTsig_15_port, 
                           OUTALU(14) => LS_OUTsig_14_port, OUTALU(13) => 
                           LS_OUTsig_13_port, OUTALU(12) => LS_OUTsig_12_port, 
                           OUTALU(11) => LS_OUTsig_11_port, OUTALU(10) => 
                           LS_OUTsig_10_port, OUTALU(9) => LS_OUTsig_9_port, 
                           OUTALU(8) => LS_OUTsig_8_port, OUTALU(7) => 
                           LS_OUTsig_7_port, OUTALU(6) => LS_OUTsig_6_port, 
                           OUTALU(5) => LS_OUTsig_5_port, OUTALU(4) => 
                           LS_OUTsig_4_port, OUTALU(3) => LS_OUTsig_3_port, 
                           OUTALU(2) => LS_OUTsig_2_port, OUTALU(1) => 
                           LS_OUTsig_1_port, OUTALU(0) => LS_OUTsig_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ZERO_DEC_bits32 is

   port( data : in std_logic_vector (31 downto 0);  zero_detect : out std_logic
         );

end ZERO_DEC_bits32;

architecture SYN_BEHAVIORAL of ZERO_DEC_bits32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n11, n12, n13, n14, n15, n16, n17, n18, n19, n20 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n11, A2 => n12, ZN => zero_detect);
   U2 : NAND4_X1 port map( A1 => n13, A2 => n14, A3 => n15, A4 => n16, ZN => 
                           n12);
   U3 : NOR4_X1 port map( A1 => data(23), A2 => data(22), A3 => data(21), A4 =>
                           data(20), ZN => n16);
   U4 : NOR4_X1 port map( A1 => data(1), A2 => data(19), A3 => data(18), A4 => 
                           data(17), ZN => n15);
   U5 : NOR4_X1 port map( A1 => data(16), A2 => data(15), A3 => data(14), A4 =>
                           data(13), ZN => n14);
   U6 : NOR4_X1 port map( A1 => data(12), A2 => data(11), A3 => data(10), A4 =>
                           data(0), ZN => n13);
   U7 : NAND4_X1 port map( A1 => n17, A2 => n18, A3 => n19, A4 => n20, ZN => 
                           n11);
   U8 : NOR4_X1 port map( A1 => data(9), A2 => data(8), A3 => data(7), A4 => 
                           data(6), ZN => n20);
   U9 : NOR4_X1 port map( A1 => data(5), A2 => data(4), A3 => data(3), A4 => 
                           data(31), ZN => n19);
   U10 : NOR4_X1 port map( A1 => data(30), A2 => data(2), A3 => data(29), A4 =>
                           data(28), ZN => n18);
   U11 : NOR4_X1 port map( A1 => data(27), A2 => data(26), A3 => data(25), A4 
                           => data(24), ZN => n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity REGISTER_FILE_NBITS32_NREGISTERS32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end REGISTER_FILE_NBITS32_NREGISTERS32;

architecture SYN_BEHAVIORAL of REGISTER_FILE_NBITS32_NREGISTERS32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, OUT1_27_port,
      OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, 
      OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, 
      OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, OUT1_12_port, 
      OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, OUT1_7_port, 
      OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, OUT1_2_port, 
      OUT1_1_port, OUT1_0_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, 
      OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, 
      OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, 
      OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, 
      OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, 
      OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, 
      OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port, n1303, n1304, n1305, 
      n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, 
      n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, 
      n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, 
      n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, 
      n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, 
      n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, 
      n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, 
      n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, 
      n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, 
      n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, 
      n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, 
      n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, 
      n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, 
      n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, 
      n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, 
      n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, 
      n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, 
      n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, 
      n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, 
      n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, 
      n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, 
      n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, 
      n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, 
      n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, 
      n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, 
      n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, 
      n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, 
      n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, 
      n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, 
      n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, 
      n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, 
      n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, 
      n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, 
      n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, 
      n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, 
      n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, 
      n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, 
      n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, 
      n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, 
      n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, 
      n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, 
      n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, 
      n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, 
      n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, 
      n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, 
      n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, 
      n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, 
      n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, 
      n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, 
      n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, 
      n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, 
      n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, 
      n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, 
      n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, 
      n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, 
      n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, 
      n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, 
      n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, 
      n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, 
      n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, 
      n2326, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, 
      n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
      n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, 
      n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, 
      n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, 
      n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, 
      n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, 
      n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, 
      n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, 
      n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, 
      n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, 
      n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, 
      n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, 
      n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, 
      n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, 
      n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, 
      n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, 
      n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, 
      n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, 
      n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, 
      n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, 
      n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, 
      n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, 
      n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, 
      n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, 
      n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, 
      n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, 
      n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, 
      n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, 
      n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, 
      n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, 
      n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, 
      n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, 
      n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, 
      n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, 
      n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, 
      n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, 
      n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, 
      n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, 
      n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, 
      n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, 
      n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, 
      n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, 
      n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, 
      n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, 
      n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, 
      n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, 
      n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, 
      n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, 
      n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, 
      n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, 
      n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, 
      n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, 
      n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, 
      n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, 
      n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, 
      n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, 
      n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, 
      n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, 
      n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, 
      n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, 
      n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, 
      n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, 
      n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, 
      n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, 
      n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, 
      n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, 
      n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, 
      n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, 
      n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, 
      n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, 
      n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, 
      n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, 
      n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, 
      n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, 
      n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, 
      n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, 
      n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, 
      n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, 
      n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, 
      n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, 
      n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, 
      n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, 
      n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, 
      n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, 
      n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, 
      n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, 
      n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, 
      n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, 
      n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, 
      n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, 
      n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, 
      n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, 
      n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, 
      n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, 
      n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, 
      n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, 
      n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, 
      n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, 
      n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, 
      n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, 
      n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, 
      n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, 
      n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, 
      n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, 
      n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, 
      n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, 
      n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, 
      n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, 
      n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, 
      n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, 
      n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, 
      n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, 
      n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, 
      n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, 
      n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, 
      n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, 
      n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, 
      n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, 
      n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, 
      n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, 
      n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, 
      n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, 
      n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, 
      n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, 
      n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, 
      n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, 
      n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, 
      n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, 
      n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, 
      n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, 
      n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, 
      n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, 
      n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, 
      n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, 
      n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, 
      n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, 
      n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, 
      n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, 
      n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, 
      n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, 
      n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, 
      n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, 
      n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, 
      n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, 
      n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, 
      n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, 
      n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, 
      n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, 
      n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, 
      n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, 
      n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, 
      n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, 
      n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, 
      n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, 
      n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, 
      n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, 
      n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, 
      n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, 
      n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, 
      n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, 
      n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, 
      n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, 
      n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, 
      n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, 
      n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, 
      n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, 
      n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, 
      n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, 
      n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, 
      n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, 
      n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, 
      n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, 
      n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, 
      n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, 
      n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, 
      n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, 
      n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, 
      n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, 
      n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, 
      n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, 
      n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, 
      n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, 
      n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, 
      n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, 
      n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, 
      n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, 
      n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, 
      n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, 
      n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, 
      n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, 
      n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, 
      n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, 
      n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, 
      n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, 
      n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, 
      n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, 
      n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, 
      n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, 
      n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, 
      n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, 
      n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, 
      n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, 
      n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, 
      n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, 
      n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, 
      n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, 
      n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, 
      n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, 
      n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, 
      n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, 
      n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, 
      n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, 
      n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, 
      n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, 
      n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, 
      n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, 
      n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, 
      n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, 
      n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, 
      n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, 
      n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, 
      n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, 
      n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, 
      n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, 
      n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, 
      n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, 
      n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, 
      n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, 
      n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, 
      n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, 
      n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, 
      n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, 
      n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, 
      n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, 
      n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, 
      n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, 
      n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, 
      n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, 
      n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, 
      n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, 
      n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, 
      n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, 
      n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, 
      n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, 
      n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, 
      n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, 
      n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, 
      n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, 
      n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, 
      n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, 
      n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, 
      n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, 
      n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, 
      n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, 
      n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, 
      n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, 
      n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, 
      n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, 
      n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, 
      n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, 
      n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, 
      n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, 
      n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, 
      n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, 
      n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, 
      n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, 
      n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, 
      n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, 
      n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, 
      n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, 
      n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, 
      n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, 
      n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, 
      n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, 
      n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, 
      n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, 
      n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, 
      n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, 
      n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, 
      n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, 
      n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, 
      n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, 
      n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, 
      n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, 
      n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, 
      n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, 
      n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, 
      n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, 
      n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, 
      n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, 
      n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, 
      n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, 
      n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, 
      n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, 
      n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, 
      n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, 
      n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, 
      n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, 
      n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, 
      n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, 
      n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, 
      n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, 
      n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, 
      n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, 
      n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, 
      n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, 
      n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, 
      n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, 
      n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, 
      n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, 
      n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, 
      n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, 
      n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, 
      n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, 
      n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, 
      n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, 
      n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, 
      n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, 
      n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, 
      n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, 
      n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, 
      n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, 
      n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, 
      n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, 
      n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, 
      n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, 
      n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, 
      n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, 
      n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, 
      n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, 
      n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, 
      n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, 
      n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, 
      n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, 
      n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, 
      n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, 
      n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, 
      n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, 
      n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, 
      n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, 
      n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, 
      n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, 
      n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, 
      n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, 
      n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, 
      n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, 
      n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, 
      n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, 
      n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, 
      n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, 
      n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, 
      n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, 
      n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, 
      n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, 
      n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, 
      n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, 
      n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, 
      n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, 
      n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, 
      n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, 
      n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, 
      n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, 
      n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, 
      n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, 
      n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, 
      n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, 
      n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, 
      n_2043 : std_logic;

begin
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   OUT2_reg_31_inst : DFF_X1 port map( D => n4130, CK => n5285, Q => 
                           OUT2_31_port, QN => n_1404);
   OUT2_reg_30_inst : DFF_X1 port map( D => n4129, CK => n5223, Q => 
                           OUT2_30_port, QN => n_1405);
   OUT2_reg_29_inst : DFF_X1 port map( D => n4128, CK => n5227, Q => 
                           OUT2_29_port, QN => n_1406);
   OUT2_reg_28_inst : DFF_X1 port map( D => n4127, CK => n5230, Q => 
                           OUT2_28_port, QN => n_1407);
   OUT2_reg_27_inst : DFF_X1 port map( D => n4126, CK => n5233, Q => 
                           OUT2_27_port, QN => n_1408);
   OUT2_reg_26_inst : DFF_X1 port map( D => n4125, CK => n5236, Q => 
                           OUT2_26_port, QN => n_1409);
   OUT2_reg_25_inst : DFF_X1 port map( D => n4124, CK => n5239, Q => 
                           OUT2_25_port, QN => n_1410);
   OUT2_reg_24_inst : DFF_X1 port map( D => n4123, CK => n5242, Q => 
                           OUT2_24_port, QN => n_1411);
   OUT2_reg_23_inst : DFF_X1 port map( D => n4122, CK => n5245, Q => 
                           OUT2_23_port, QN => n_1412);
   OUT2_reg_22_inst : DFF_X1 port map( D => n4121, CK => n5248, Q => 
                           OUT2_22_port, QN => n_1413);
   OUT2_reg_21_inst : DFF_X1 port map( D => n4120, CK => n5251, Q => 
                           OUT2_21_port, QN => n_1414);
   OUT2_reg_20_inst : DFF_X1 port map( D => n4119, CK => n5254, Q => 
                           OUT2_20_port, QN => n_1415);
   OUT2_reg_19_inst : DFF_X1 port map( D => n4118, CK => n5257, Q => 
                           OUT2_19_port, QN => n_1416);
   OUT2_reg_18_inst : DFF_X1 port map( D => n4117, CK => n5261, Q => 
                           OUT2_18_port, QN => n_1417);
   OUT2_reg_17_inst : DFF_X1 port map( D => n4116, CK => n5264, Q => 
                           OUT2_17_port, QN => n_1418);
   OUT2_reg_16_inst : DFF_X1 port map( D => n4115, CK => n5267, Q => 
                           OUT2_16_port, QN => n_1419);
   OUT2_reg_15_inst : DFF_X1 port map( D => n4114, CK => n5270, Q => 
                           OUT2_15_port, QN => n_1420);
   OUT2_reg_14_inst : DFF_X1 port map( D => n4113, CK => n5273, Q => 
                           OUT2_14_port, QN => n_1421);
   OUT2_reg_13_inst : DFF_X1 port map( D => n4112, CK => n5276, Q => 
                           OUT2_13_port, QN => n_1422);
   OUT2_reg_12_inst : DFF_X1 port map( D => n4111, CK => n5279, Q => 
                           OUT2_12_port, QN => n_1423);
   OUT2_reg_11_inst : DFF_X1 port map( D => n4110, CK => n5282, Q => 
                           OUT2_11_port, QN => n_1424);
   OUT2_reg_10_inst : DFF_X1 port map( D => n4109, CK => n5202, Q => 
                           OUT2_10_port, QN => n_1425);
   OUT2_reg_9_inst : DFF_X1 port map( D => n4108, CK => n5205, Q => OUT2_9_port
                           , QN => n_1426);
   OUT2_reg_8_inst : DFF_X1 port map( D => n4107, CK => n5208, Q => OUT2_8_port
                           , QN => n_1427);
   OUT2_reg_7_inst : DFF_X1 port map( D => n4106, CK => n5211, Q => OUT2_7_port
                           , QN => n_1428);
   OUT2_reg_6_inst : DFF_X1 port map( D => n4105, CK => n5214, Q => OUT2_6_port
                           , QN => n_1429);
   OUT2_reg_5_inst : DFF_X1 port map( D => n4104, CK => n5217, Q => OUT2_5_port
                           , QN => n_1430);
   OUT2_reg_4_inst : DFF_X1 port map( D => n4103, CK => n5220, Q => OUT2_4_port
                           , QN => n_1431);
   OUT2_reg_3_inst : DFF_X1 port map( D => n4102, CK => n5196, Q => OUT2_3_port
                           , QN => n_1432);
   OUT2_reg_2_inst : DFF_X1 port map( D => n4101, CK => n5199, Q => OUT2_2_port
                           , QN => n_1433);
   OUT2_reg_1_inst : DFF_X1 port map( D => n4100, CK => n5288, Q => OUT2_1_port
                           , QN => n_1434);
   OUT2_reg_0_inst : DFF_X1 port map( D => n4099, CK => n5291, Q => OUT2_0_port
                           , QN => n_1435);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2326, CK => n5285, Q => 
                           n_1436, QN => n4485);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2325, CK => n5224, Q => 
                           n_1437, QN => n4486);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2324, CK => n5227, Q => 
                           n_1438, QN => n4487);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2323, CK => n5230, Q => 
                           n_1439, QN => n4488);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2322, CK => n5233, Q => 
                           n_1440, QN => n4489);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2321, CK => n5236, Q => 
                           n_1441, QN => n4490);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2320, CK => n5239, Q => 
                           n_1442, QN => n4491);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2319, CK => n5242, Q => 
                           n_1443, QN => n4492);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2318, CK => n5245, Q => 
                           n_1444, QN => n4493);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2317, CK => n5248, Q => 
                           n_1445, QN => n4494);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2316, CK => n5251, Q => 
                           n_1446, QN => n4495);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2315, CK => n5254, Q => 
                           n_1447, QN => n4496);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2314, CK => n5258, Q => 
                           n_1448, QN => n4497);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2313, CK => n5261, Q => 
                           n_1449, QN => n4498);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2312, CK => n5264, Q => 
                           n_1450, QN => n4499);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2311, CK => n5267, Q => 
                           n_1451, QN => n4500);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2310, CK => n5270, Q => 
                           n_1452, QN => n4501);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2309, CK => n5273, Q => 
                           n_1453, QN => n4502);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2308, CK => n5276, Q => 
                           n_1454, QN => n4503);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2307, CK => n5279, Q => 
                           n_1455, QN => n4504);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2306, CK => n5282, Q => 
                           n_1456, QN => n4505);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2305, CK => n5202, Q => 
                           n_1457, QN => n4506);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2304, CK => n5205, Q => 
                           n_1458, QN => n4507);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2303, CK => n5208, Q => 
                           n_1459, QN => n4508);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2302, CK => n5211, Q => 
                           n_1460, QN => n4509);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2301, CK => n5214, Q => 
                           n_1461, QN => n4510);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2300, CK => n5217, Q => 
                           n_1462, QN => n4511);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2299, CK => n5220, Q => 
                           n_1463, QN => n4512);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2298, CK => n5196, Q => 
                           n_1464, QN => n4513);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2297, CK => n5199, Q => 
                           n_1465, QN => n4514);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2296, CK => n5288, Q => 
                           n_1466, QN => n4515);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2295, CK => n5292, Q => 
                           n_1467, QN => n4516);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2294, CK => n5285, Q => 
                           n6640, QN => n4965);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2293, CK => n5224, Q => 
                           n6641, QN => n4966);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2292, CK => n5227, Q => 
                           n6642, QN => n4967);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2291, CK => n5230, Q => 
                           n6643, QN => n4968);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2290, CK => n5233, Q => 
                           n6644, QN => n4969);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2289, CK => n5236, Q => 
                           n6645, QN => n4970);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2288, CK => n5239, Q => 
                           n6646, QN => n4971);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2287, CK => n5242, Q => 
                           n6647, QN => n4972);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2286, CK => n5245, Q => 
                           n6648, QN => n4973);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2285, CK => n5248, Q => 
                           n6649, QN => n4974);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2284, CK => n5251, Q => 
                           n6650, QN => n4975);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2283, CK => n5255, Q => 
                           n6651, QN => n4976);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2282, CK => n5258, Q => 
                           n6652, QN => n4977);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2281, CK => n5261, Q => 
                           n6653, QN => n4978);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2280, CK => n5264, Q => 
                           n6654, QN => n4979);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2279, CK => n5267, Q => 
                           n6655, QN => n4980);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2278, CK => n5270, Q => 
                           n6656, QN => n4981);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2277, CK => n5273, Q => 
                           n6657, QN => n4982);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2276, CK => n5276, Q => 
                           n6658, QN => n4983);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2275, CK => n5279, Q => 
                           n6659, QN => n4984);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2274, CK => n5282, Q => 
                           n6660, QN => n4985);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2273, CK => n5202, Q => 
                           n6661, QN => n4986);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2272, CK => n5205, Q => 
                           n6662, QN => n4987);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2271, CK => n5208, Q => 
                           n6663, QN => n4988);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2270, CK => n5211, Q => 
                           n6664, QN => n4989);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2269, CK => n5214, Q => 
                           n6665, QN => n4990);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2268, CK => n5217, Q => 
                           n6666, QN => n4991);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2267, CK => n5221, Q => 
                           n6667, QN => n4992);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2266, CK => n5196, Q => 
                           n6668, QN => n4993);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2265, CK => n5199, Q => 
                           n6669, QN => n4994);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2264, CK => n5289, Q => 
                           n6670, QN => n4995);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2263, CK => n5292, Q => 
                           n6671, QN => n4996);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2262, CK => n5286, Q => 
                           n6672, QN => n4997);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2261, CK => n5224, Q => 
                           n6673, QN => n4998);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2260, CK => n5227, Q => 
                           n6674, QN => n4999);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2259, CK => n5230, Q => 
                           n6675, QN => n5000);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2258, CK => n5233, Q => 
                           n6676, QN => n5001);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2257, CK => n5236, Q => 
                           n6677, QN => n5002);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2256, CK => n5239, Q => 
                           n6678, QN => n5003);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2255, CK => n5242, Q => 
                           n6679, QN => n5004);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2254, CK => n5245, Q => 
                           n6680, QN => n5005);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2253, CK => n5248, Q => 
                           n6681, QN => n5006);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2252, CK => n5252, Q => 
                           n6682, QN => n5007);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2251, CK => n5255, Q => 
                           n6683, QN => n5008);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2250, CK => n5258, Q => 
                           n6684, QN => n5009);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2249, CK => n5261, Q => 
                           n6685, QN => n5010);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2248, CK => n5264, Q => 
                           n6686, QN => n5011);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2247, CK => n5267, Q => 
                           n6687, QN => n5012);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2246, CK => n5270, Q => 
                           n6688, QN => n5013);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2245, CK => n5273, Q => 
                           n6689, QN => n5014);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2244, CK => n5276, Q => 
                           n6690, QN => n5015);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2243, CK => n5279, Q => 
                           n6691, QN => n5016);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2242, CK => n5282, Q => 
                           n6692, QN => n5017);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2241, CK => n5202, Q => 
                           n6693, QN => n5018);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2240, CK => n5205, Q => 
                           n6694, QN => n5019);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2239, CK => n5208, Q => 
                           n6695, QN => n5020);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2238, CK => n5211, Q => 
                           n6696, QN => n5021);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2237, CK => n5214, Q => 
                           n6697, QN => n5022);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2236, CK => n5218, Q => 
                           n6698, QN => n5023);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2235, CK => n5221, Q => 
                           n6699, QN => n5024);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2234, CK => n5196, Q => 
                           n6700, QN => n5025);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2233, CK => n5199, Q => 
                           n6701, QN => n5026);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2232, CK => n5289, Q => 
                           n6702, QN => n5027);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2231, CK => n5292, Q => 
                           n6703, QN => n5028);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2230, CK => n5286, Q => 
                           n6704, QN => n4741);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2229, CK => n5224, Q => 
                           n6705, QN => n4742);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2228, CK => n5227, Q => 
                           n6706, QN => n4743);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2227, CK => n5230, Q => 
                           n6707, QN => n4744);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2226, CK => n5233, Q => 
                           n6708, QN => n4745);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2225, CK => n5236, Q => 
                           n6709, QN => n4746);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2224, CK => n5239, Q => 
                           n6710, QN => n4747);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2223, CK => n5242, Q => 
                           n6711, QN => n4748);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2222, CK => n5245, Q => 
                           n6712, QN => n4749);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2221, CK => n5249, Q => 
                           n6713, QN => n4750);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2220, CK => n5252, Q => 
                           n6714, QN => n4751);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2219, CK => n5255, Q => 
                           n6715, QN => n4752);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2218, CK => n5258, Q => 
                           n6716, QN => n4753);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2217, CK => n5261, Q => 
                           n6717, QN => n4754);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2216, CK => n5264, Q => 
                           n6718, QN => n4755);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2215, CK => n5267, Q => 
                           n6719, QN => n4756);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2214, CK => n5270, Q => 
                           n6720, QN => n4757);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2213, CK => n5273, Q => 
                           n6721, QN => n4758);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2212, CK => n5276, Q => 
                           n6722, QN => n4759);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2211, CK => n5279, Q => 
                           n6723, QN => n4760);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2210, CK => n5283, Q => 
                           n6724, QN => n4761);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2209, CK => n5202, Q => 
                           n6725, QN => n4762);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2208, CK => n5205, Q => 
                           n6726, QN => n4763);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2207, CK => n5208, Q => 
                           n6727, QN => n4764);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2206, CK => n5211, Q => 
                           n6728, QN => n4765);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2205, CK => n5215, Q => 
                           n6729, QN => n4766);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2204, CK => n5218, Q => 
                           n6730, QN => n4767);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2203, CK => n5221, Q => 
                           n6731, QN => n4768);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2202, CK => n5196, Q => 
                           n6732, QN => n4769);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2201, CK => n5199, Q => 
                           n6733, QN => n4770);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2200, CK => n5289, Q => 
                           n6734, QN => n4771);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2199, CK => n5292, Q => 
                           n6735, QN => n4772);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2198, CK => n5286, Q => 
                           n6736, QN => n4773);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2197, CK => n5224, Q => 
                           n6737, QN => n4774);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2196, CK => n5227, Q => 
                           n6738, QN => n4775);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2195, CK => n5230, Q => 
                           n6739, QN => n4776);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2194, CK => n5233, Q => 
                           n6740, QN => n4777);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2193, CK => n5236, Q => 
                           n6741, QN => n4778);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2192, CK => n5239, Q => 
                           n6742, QN => n4779);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2191, CK => n5242, Q => 
                           n6743, QN => n4780);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2190, CK => n5246, Q => 
                           n6744, QN => n4781);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2189, CK => n5249, Q => 
                           n6745, QN => n4782);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2188, CK => n5252, Q => 
                           n6746, QN => n4783);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2187, CK => n5255, Q => 
                           n6747, QN => n4784);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2186, CK => n5258, Q => 
                           n6748, QN => n4785);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2185, CK => n5261, Q => 
                           n6749, QN => n4786);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2184, CK => n5264, Q => 
                           n6750, QN => n4787);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2183, CK => n5267, Q => 
                           n6751, QN => n4788);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2182, CK => n5270, Q => 
                           n6752, QN => n4789);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2181, CK => n5273, Q => 
                           n6753, QN => n4790);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2180, CK => n5276, Q => 
                           n6754, QN => n4791);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2179, CK => n5280, Q => 
                           n6755, QN => n4792);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2178, CK => n5283, Q => 
                           n6756, QN => n4793);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2177, CK => n5202, Q => 
                           n6757, QN => n4794);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2176, CK => n5205, Q => 
                           n6758, QN => n4795);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2175, CK => n5208, Q => 
                           n6759, QN => n4796);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2174, CK => n5212, Q => 
                           n6760, QN => n4797);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2173, CK => n5215, Q => 
                           n6761, QN => n4798);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2172, CK => n5218, Q => 
                           n6762, QN => n4799);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2171, CK => n5221, Q => 
                           n6763, QN => n4800);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2170, CK => n5196, Q => 
                           n6764, QN => n4801);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2169, CK => n5199, Q => 
                           n6765, QN => n4802);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2168, CK => n5289, Q => 
                           n6766, QN => n4803);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2167, CK => n5292, Q => 
                           n6767, QN => n4804);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2166, CK => n5286, Q => 
                           n_1468, QN => n4163);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2165, CK => n5224, Q => 
                           n_1469, QN => n4164);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2164, CK => n5227, Q => 
                           n_1470, QN => n4165);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2163, CK => n5230, Q => 
                           n_1471, QN => n4166);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2162, CK => n5233, Q => 
                           n_1472, QN => n4167);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2161, CK => n5236, Q => 
                           n_1473, QN => n4168);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2160, CK => n5239, Q => 
                           n_1474, QN => n4169);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n2159, CK => n5243, Q => 
                           n_1475, QN => n4170);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n2158, CK => n5246, Q => 
                           n_1476, QN => n4171);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n2157, CK => n5249, Q => 
                           n_1477, QN => n4172);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n2156, CK => n5252, Q => 
                           n_1478, QN => n4173);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n2155, CK => n5255, Q => 
                           n_1479, QN => n4174);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n2154, CK => n5258, Q => 
                           n_1480, QN => n4175);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n2153, CK => n5261, Q => 
                           n_1481, QN => n4176);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n2152, CK => n5264, Q => 
                           n_1482, QN => n4177);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n2151, CK => n5267, Q => 
                           n_1483, QN => n4178);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n2150, CK => n5270, Q => 
                           n_1484, QN => n4179);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n2149, CK => n5273, Q => 
                           n_1485, QN => n4180);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n2148, CK => n5277, Q => 
                           n_1486, QN => n4181);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n2147, CK => n5280, Q => 
                           n_1487, QN => n4182);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n2146, CK => n5283, Q => 
                           n_1488, QN => n4183);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n2145, CK => n5202, Q => 
                           n_1489, QN => n4184);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n2144, CK => n5205, Q => 
                           n_1490, QN => n4185);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n2143, CK => n5209, Q => 
                           n_1491, QN => n4186);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n2142, CK => n5212, Q => 
                           n_1492, QN => n4187);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n2141, CK => n5215, Q => 
                           n_1493, QN => n4188);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n2140, CK => n5218, Q => 
                           n_1494, QN => n4189);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n2139, CK => n5221, Q => 
                           n_1495, QN => n4190);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n2138, CK => n5196, Q => 
                           n_1496, QN => n4191);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n2137, CK => n5199, Q => 
                           n_1497, QN => n4192);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n2136, CK => n5289, Q => 
                           n_1498, QN => n4193);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n2135, CK => n5292, Q => 
                           n_1499, QN => n4194);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n2134, CK => n5286, Q => 
                           n_1500, QN => n4677);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n2133, CK => n5224, Q => 
                           n_1501, QN => n4678);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n2132, CK => n5227, Q => 
                           n_1502, QN => n4679);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n2131, CK => n5230, Q => 
                           n_1503, QN => n4680);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n2130, CK => n5233, Q => 
                           n_1504, QN => n4681);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n2129, CK => n5236, Q => 
                           n_1505, QN => n4682);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n2128, CK => n5240, Q => 
                           n_1506, QN => n4683);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n2127, CK => n5243, Q => 
                           n_1507, QN => n4684);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n2126, CK => n5246, Q => 
                           n_1508, QN => n4685);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n2125, CK => n5249, Q => 
                           n_1509, QN => n4686);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n2124, CK => n5252, Q => 
                           n_1510, QN => n4687);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n2123, CK => n5255, Q => 
                           n_1511, QN => n4688);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n2122, CK => n5258, Q => 
                           n_1512, QN => n4689);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n2121, CK => n5261, Q => 
                           n_1513, QN => n4690);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n2120, CK => n5264, Q => 
                           n_1514, QN => n4691);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n2119, CK => n5267, Q => 
                           n_1515, QN => n4692);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n2118, CK => n5270, Q => 
                           n_1516, QN => n4693);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n2117, CK => n5274, Q => 
                           n_1517, QN => n4694);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n2116, CK => n5277, Q => 
                           n_1518, QN => n4695);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n2115, CK => n5280, Q => 
                           n_1519, QN => n4696);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n2114, CK => n5283, Q => 
                           n_1520, QN => n4697);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n2113, CK => n5202, Q => 
                           n_1521, QN => n4698);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n2112, CK => n5206, Q => 
                           n_1522, QN => n4699);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n2111, CK => n5209, Q => 
                           n_1523, QN => n4700);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n2110, CK => n5212, Q => 
                           n_1524, QN => n4701);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n2109, CK => n5215, Q => 
                           n_1525, QN => n4702);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n2108, CK => n5218, Q => 
                           n_1526, QN => n4703);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n2107, CK => n5221, Q => 
                           n_1527, QN => n4704);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n2106, CK => n5196, Q => 
                           n_1528, QN => n4705);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n2105, CK => n5199, Q => 
                           n_1529, QN => n4706);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n2104, CK => n5289, Q => 
                           n_1530, QN => n4707);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n2103, CK => n5292, Q => 
                           n_1531, QN => n4708);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n2102, CK => n5286, Q => 
                           n_1532, QN => n4419);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n2101, CK => n5224, Q => 
                           n_1533, QN => n4420);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n2100, CK => n5227, Q => 
                           n_1534, QN => n4421);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n2099, CK => n5230, Q => 
                           n_1535, QN => n4422);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n2098, CK => n5233, Q => 
                           n_1536, QN => n4423);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n2097, CK => n5237, Q => 
                           n_1537, QN => n4424);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n2096, CK => n5240, Q => 
                           n_1538, QN => n4425);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n2095, CK => n5243, Q => 
                           n_1539, QN => n4426);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n2094, CK => n5246, Q => 
                           n_1540, QN => n4427);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n2093, CK => n5249, Q => 
                           n_1541, QN => n4428);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n2092, CK => n5252, Q => 
                           n_1542, QN => n4429);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n2091, CK => n5255, Q => 
                           n_1543, QN => n4430);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n2090, CK => n5258, Q => 
                           n_1544, QN => n4431);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n2089, CK => n5261, Q => 
                           n_1545, QN => n4432);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n2088, CK => n5264, Q => 
                           n_1546, QN => n4433);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n2087, CK => n5267, Q => 
                           n_1547, QN => n4434);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n2086, CK => n5271, Q => 
                           n_1548, QN => n4435);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n2085, CK => n5274, Q => 
                           n_1549, QN => n4436);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n2084, CK => n5277, Q => 
                           n_1550, QN => n4437);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n2083, CK => n5280, Q => 
                           n_1551, QN => n4438);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n2082, CK => n5283, Q => 
                           n_1552, QN => n4439);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n2081, CK => n5203, Q => 
                           n_1553, QN => n4440);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n2080, CK => n5206, Q => 
                           n_1554, QN => n4441);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n2079, CK => n5209, Q => 
                           n_1555, QN => n4442);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n2078, CK => n5212, Q => 
                           n_1556, QN => n4443);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n2077, CK => n5215, Q => 
                           n_1557, QN => n4444);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n2076, CK => n5218, Q => 
                           n_1558, QN => n4445);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n2075, CK => n5221, Q => 
                           n_1559, QN => n4446);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n2074, CK => n5196, Q => 
                           n_1560, QN => n4447);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n2073, CK => n5200, Q => 
                           n_1561, QN => n4448);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n2072, CK => n5289, Q => 
                           n_1562, QN => n4449);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n2071, CK => n5292, Q => 
                           n_1563, QN => n4450);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n2070, CK => n5286, Q => 
                           n6768, QN => n4805);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n2069, CK => n5224, Q => 
                           n6769, QN => n4806);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n2068, CK => n5227, Q => 
                           n6770, QN => n4807);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n2067, CK => n5230, Q => 
                           n6771, QN => n4808);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n2066, CK => n5234, Q => 
                           n6772, QN => n4809);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n2065, CK => n5237, Q => 
                           n6773, QN => n4810);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n2064, CK => n5240, Q => 
                           n6774, QN => n4811);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n2063, CK => n5243, Q => 
                           n6775, QN => n4812);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n2062, CK => n5246, Q => 
                           n6776, QN => n4813);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n2061, CK => n5249, Q => 
                           n6777, QN => n4814);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n2060, CK => n5252, Q => 
                           n6778, QN => n4815);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n2059, CK => n5255, Q => 
                           n6779, QN => n4816);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n2058, CK => n5258, Q => 
                           n6780, QN => n4817);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n2057, CK => n5261, Q => 
                           n6781, QN => n4818);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n2056, CK => n5264, Q => 
                           n6782, QN => n4819);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n2055, CK => n5268, Q => 
                           n6783, QN => n4820);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n2054, CK => n5271, Q => 
                           n6784, QN => n4821);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n2053, CK => n5274, Q => 
                           n6785, QN => n4822);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n2052, CK => n5277, Q => 
                           n6786, QN => n4823);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n2051, CK => n5280, Q => 
                           n6787, QN => n4824);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n2050, CK => n5283, Q => 
                           n6788, QN => n4825);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n2049, CK => n5203, Q => 
                           n6789, QN => n4826);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n2048, CK => n5206, Q => 
                           n6790, QN => n4827);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n2047, CK => n5209, Q => 
                           n6791, QN => n4828);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n2046, CK => n5212, Q => 
                           n6792, QN => n4829);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n2045, CK => n5215, Q => 
                           n6793, QN => n4830);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n2044, CK => n5218, Q => 
                           n6794, QN => n4831);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n2043, CK => n5221, Q => 
                           n6795, QN => n4832);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n2042, CK => n5197, Q => 
                           n6796, QN => n4833);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n2041, CK => n5200, Q => 
                           n6797, QN => n4834);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n2040, CK => n5289, Q => 
                           n6798, QN => n4835);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n2039, CK => n5292, Q => 
                           n6799, QN => n4836);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n2038, CK => n5286, Q => 
                           n_1564, QN => n4227);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n2037, CK => n5224, Q => 
                           n_1565, QN => n4228);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n2036, CK => n5227, Q => 
                           n_1566, QN => n4229);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n2035, CK => n5231, Q => 
                           n_1567, QN => n4230);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n2034, CK => n5234, Q => 
                           n_1568, QN => n4231);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n2033, CK => n5237, Q => 
                           n_1569, QN => n4232);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n2032, CK => n5240, Q => 
                           n_1570, QN => n4233);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n2031, CK => n5243, Q => 
                           n_1571, QN => n4234);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n2030, CK => n5246, Q => 
                           n_1572, QN => n4235);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n2029, CK => n5249, Q => 
                           n_1573, QN => n4236);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n2028, CK => n5252, Q => 
                           n_1574, QN => n4237);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n2027, CK => n5255, Q => 
                           n_1575, QN => n4238);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n2026, CK => n5258, Q => 
                           n_1576, QN => n4239);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n2025, CK => n5261, Q => 
                           n_1577, QN => n4240);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n2024, CK => n5265, Q => 
                           n_1578, QN => n4241);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n2023, CK => n5268, Q => 
                           n_1579, QN => n4242);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n2022, CK => n5271, Q => 
                           n_1580, QN => n4243);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n2021, CK => n5274, Q => 
                           n_1581, QN => n4244);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n2020, CK => n5277, Q => 
                           n_1582, QN => n4245);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n2019, CK => n5280, Q => 
                           n_1583, QN => n4246);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n2018, CK => n5283, Q => 
                           n_1584, QN => n4247);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n2017, CK => n5203, Q => 
                           n_1585, QN => n4248);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n2016, CK => n5206, Q => 
                           n_1586, QN => n4249);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n2015, CK => n5209, Q => 
                           n_1587, QN => n4250);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n2014, CK => n5212, Q => 
                           n_1588, QN => n4251);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n2013, CK => n5215, Q => 
                           n_1589, QN => n4252);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n2012, CK => n5218, Q => 
                           n_1590, QN => n4253);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n2011, CK => n5221, Q => 
                           n_1591, QN => n4254);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n2010, CK => n5197, Q => 
                           n_1592, QN => n4255);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n2009, CK => n5200, Q => 
                           n_1593, QN => n4256);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n2008, CK => n5289, Q => 
                           n_1594, QN => n4257);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n2007, CK => n5292, Q => 
                           n_1595, QN => n4258);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n2006, CK => n5286, Q => 
                           n_1596, QN => n4195);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n2005, CK => n5224, Q => 
                           n_1597, QN => n4196);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n2004, CK => n5228, Q => 
                           n_1598, QN => n4197);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n2003, CK => n5231, Q => 
                           n_1599, QN => n4198);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n2002, CK => n5234, Q => 
                           n_1600, QN => n4199);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n2001, CK => n5237, Q => 
                           n_1601, QN => n4200);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n2000, CK => n5240, Q => 
                           n_1602, QN => n4201);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1999, CK => n5243, Q => 
                           n_1603, QN => n4202);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1998, CK => n5246, Q => 
                           n_1604, QN => n4203);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1997, CK => n5249, Q => 
                           n_1605, QN => n4204);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1996, CK => n5252, Q => 
                           n_1606, QN => n4205);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1995, CK => n5255, Q => 
                           n_1607, QN => n4206);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1994, CK => n5258, Q => 
                           n_1608, QN => n4207);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1993, CK => n5262, Q => 
                           n_1609, QN => n4208);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1992, CK => n5265, Q => 
                           n_1610, QN => n4209);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1991, CK => n5268, Q => 
                           n_1611, QN => n4210);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1990, CK => n5271, Q => 
                           n_1612, QN => n4211);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1989, CK => n5274, Q => 
                           n_1613, QN => n4212);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1988, CK => n5277, Q => 
                           n_1614, QN => n4213);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1987, CK => n5280, Q => 
                           n_1615, QN => n4214);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1986, CK => n5283, Q => 
                           n_1616, QN => n4215);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1985, CK => n5203, Q => 
                           n_1617, QN => n4216);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1984, CK => n5206, Q => 
                           n_1618, QN => n4217);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1983, CK => n5209, Q => 
                           n_1619, QN => n4218);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1982, CK => n5212, Q => 
                           n_1620, QN => n4219);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1981, CK => n5215, Q => 
                           n_1621, QN => n4220);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1980, CK => n5218, Q => 
                           n_1622, QN => n4221);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1979, CK => n5221, Q => 
                           n_1623, QN => n4222);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1978, CK => n5197, Q => 
                           n_1624, QN => n4223);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1977, CK => n5200, Q => 
                           n_1625, QN => n4224);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1976, CK => n5289, Q => 
                           n_1626, QN => n4225);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1975, CK => n5292, Q => 
                           n_1627, QN => n4226);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1974, CK => n5286, Q => 
                           n6800, QN => n5029);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1973, CK => n5225, Q => 
                           n6801, QN => n5030);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1972, CK => n5228, Q => 
                           n6802, QN => n5031);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1971, CK => n5231, Q => 
                           n6803, QN => n5032);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1970, CK => n5234, Q => 
                           n6804, QN => n5033);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1969, CK => n5237, Q => 
                           n6805, QN => n5034);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1968, CK => n5240, Q => 
                           n6806, QN => n5035);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1967, CK => n5243, Q => 
                           n6807, QN => n5036);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1966, CK => n5246, Q => 
                           n6808, QN => n5037);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1965, CK => n5249, Q => 
                           n6809, QN => n5038);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1964, CK => n5252, Q => 
                           n6810, QN => n5039);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1963, CK => n5255, Q => 
                           n6811, QN => n5040);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1962, CK => n5259, Q => 
                           n6812, QN => n5041);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1961, CK => n5262, Q => 
                           n6813, QN => n5042);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1960, CK => n5265, Q => 
                           n6814, QN => n5043);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1959, CK => n5268, Q => 
                           n6815, QN => n5044);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1958, CK => n5271, Q => 
                           n6816, QN => n5045);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1957, CK => n5274, Q => 
                           n6817, QN => n5046);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1956, CK => n5277, Q => 
                           n6818, QN => n5047);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1955, CK => n5280, Q => 
                           n6819, QN => n5048);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1954, CK => n5283, Q => 
                           n6820, QN => n5049);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1953, CK => n5203, Q => 
                           n6821, QN => n5050);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1952, CK => n5206, Q => 
                           n6822, QN => n5051);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1951, CK => n5209, Q => 
                           n6823, QN => n5052);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1950, CK => n5212, Q => 
                           n6824, QN => n5053);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1949, CK => n5215, Q => 
                           n6825, QN => n5054);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1948, CK => n5218, Q => 
                           n6826, QN => n5055);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1947, CK => n5221, Q => 
                           n6827, QN => n5056);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1946, CK => n5197, Q => 
                           n6828, QN => n5057);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1945, CK => n5200, Q => 
                           n6829, QN => n5058);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1944, CK => n5289, Q => 
                           n6830, QN => n5059);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1943, CK => n5293, Q => 
                           n6831, QN => n5060);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1942, CK => n5286, Q => 
                           n6832, QN => n5061);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1941, CK => n5225, Q => 
                           n6833, QN => n5062);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1940, CK => n5228, Q => 
                           n6834, QN => n5063);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1939, CK => n5231, Q => 
                           n6835, QN => n5064);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1938, CK => n5234, Q => 
                           n6836, QN => n5065);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1937, CK => n5237, Q => 
                           n6837, QN => n5066);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1936, CK => n5240, Q => 
                           n6838, QN => n5067);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1935, CK => n5243, Q => 
                           n6839, QN => n5068);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1934, CK => n5246, Q => 
                           n6840, QN => n5069);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1933, CK => n5249, Q => 
                           n6841, QN => n5070);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1932, CK => n5252, Q => 
                           n6842, QN => n5071);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1931, CK => n5256, Q => 
                           n6843, QN => n5072);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1930, CK => n5259, Q => 
                           n6844, QN => n5073);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1929, CK => n5262, Q => 
                           n6845, QN => n5074);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1928, CK => n5265, Q => 
                           n6846, QN => n5075);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1927, CK => n5268, Q => 
                           n6847, QN => n5076);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1926, CK => n5271, Q => 
                           n6848, QN => n5077);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1925, CK => n5274, Q => 
                           n6849, QN => n5078);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1924, CK => n5277, Q => 
                           n6850, QN => n5079);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1923, CK => n5280, Q => 
                           n6851, QN => n5080);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1922, CK => n5283, Q => 
                           n6852, QN => n5081);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1921, CK => n5203, Q => 
                           n6853, QN => n5082);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1920, CK => n5206, Q => 
                           n6854, QN => n5083);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1919, CK => n5209, Q => 
                           n6855, QN => n5084);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1918, CK => n5212, Q => 
                           n6856, QN => n5085);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1917, CK => n5215, Q => 
                           n6857, QN => n5086);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1916, CK => n5218, Q => 
                           n6858, QN => n5087);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1915, CK => n5222, Q => 
                           n6859, QN => n5088);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1914, CK => n5197, Q => 
                           n6860, QN => n5089);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1913, CK => n5200, Q => 
                           n6861, QN => n5090);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1912, CK => n5290, Q => 
                           n6862, QN => n5091);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1911, CK => n5293, Q => 
                           n6863, QN => n5092);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1910, CK => n5287, Q => 
                           n_1628, QN => n4709);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1909, CK => n5225, Q => 
                           n_1629, QN => n4710);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1908, CK => n5228, Q => 
                           n_1630, QN => n4711);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1907, CK => n5231, Q => 
                           n_1631, QN => n4712);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1906, CK => n5234, Q => 
                           n_1632, QN => n4713);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1905, CK => n5237, Q => 
                           n_1633, QN => n4714);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1904, CK => n5240, Q => 
                           n_1634, QN => n4715);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1903, CK => n5243, Q => 
                           n_1635, QN => n4716);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1902, CK => n5246, Q => 
                           n_1636, QN => n4717);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1901, CK => n5249, Q => 
                           n_1637, QN => n4718);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1900, CK => n5253, Q => 
                           n_1638, QN => n4719);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1899, CK => n5256, Q => 
                           n_1639, QN => n4720);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1898, CK => n5259, Q => 
                           n_1640, QN => n4721);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1897, CK => n5262, Q => 
                           n_1641, QN => n4722);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1896, CK => n5265, Q => 
                           n_1642, QN => n4723);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1895, CK => n5268, Q => 
                           n_1643, QN => n4724);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1894, CK => n5271, Q => 
                           n_1644, QN => n4725);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1893, CK => n5274, Q => 
                           n_1645, QN => n4726);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1892, CK => n5277, Q => 
                           n_1646, QN => n4727);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1891, CK => n5280, Q => 
                           n_1647, QN => n4728);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1890, CK => n5283, Q => 
                           n_1648, QN => n4729);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1889, CK => n5203, Q => 
                           n_1649, QN => n4730);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1888, CK => n5206, Q => 
                           n_1650, QN => n4731);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1887, CK => n5209, Q => 
                           n_1651, QN => n4732);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1886, CK => n5212, Q => 
                           n_1652, QN => n4733);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1885, CK => n5215, Q => 
                           n_1653, QN => n4734);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1884, CK => n5219, Q => 
                           n_1654, QN => n4735);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1883, CK => n5222, Q => 
                           n_1655, QN => n4736);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1882, CK => n5197, Q => 
                           n_1656, QN => n4737);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1881, CK => n5200, Q => 
                           n_1657, QN => n4738);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1880, CK => n5290, Q => 
                           n_1658, QN => n4739);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1879, CK => n5293, Q => 
                           n_1659, QN => n4740);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1878, CK => n5287, Q => 
                           n_1660, QN => n4451);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1877, CK => n5225, Q => 
                           n_1661, QN => n4452);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1876, CK => n5228, Q => 
                           n_1662, QN => n4453);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1875, CK => n5231, Q => 
                           n_1663, QN => n4454);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1874, CK => n5234, Q => 
                           n_1664, QN => n4455);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1873, CK => n5237, Q => 
                           n_1665, QN => n4456);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1872, CK => n5240, Q => 
                           n_1666, QN => n4457);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1871, CK => n5243, Q => 
                           n_1667, QN => n4458);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1870, CK => n5246, Q => 
                           n_1668, QN => n4459);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1869, CK => n5250, Q => 
                           n_1669, QN => n4460);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1868, CK => n5253, Q => 
                           n_1670, QN => n4461);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1867, CK => n5256, Q => 
                           n_1671, QN => n4462);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1866, CK => n5259, Q => 
                           n_1672, QN => n4463);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1865, CK => n5262, Q => 
                           n_1673, QN => n4464);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1864, CK => n5265, Q => 
                           n_1674, QN => n4465);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1863, CK => n5268, Q => 
                           n_1675, QN => n4466);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1862, CK => n5271, Q => 
                           n_1676, QN => n4467);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1861, CK => n5274, Q => 
                           n_1677, QN => n4468);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1860, CK => n5277, Q => 
                           n_1678, QN => n4469);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1859, CK => n5280, Q => 
                           n_1679, QN => n4470);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1858, CK => n5284, Q => 
                           n_1680, QN => n4471);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1857, CK => n5203, Q => 
                           n_1681, QN => n4472);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1856, CK => n5206, Q => 
                           n_1682, QN => n4473);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1855, CK => n5209, Q => 
                           n_1683, QN => n4474);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1854, CK => n5212, Q => 
                           n_1684, QN => n4475);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1853, CK => n5216, Q => 
                           n_1685, QN => n4476);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1852, CK => n5219, Q => 
                           n_1686, QN => n4477);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1851, CK => n5222, Q => 
                           n_1687, QN => n4478);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1850, CK => n5197, Q => 
                           n_1688, QN => n4479);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1849, CK => n5200, Q => 
                           n_1689, QN => n4480);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1848, CK => n5290, Q => 
                           n_1690, QN => n4481);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1847, CK => n5293, Q => 
                           n_1691, QN => n4482);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1846, CK => n5287, Q => 
                           n6864, QN => n4837);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1845, CK => n5225, Q => 
                           n6865, QN => n4838);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1844, CK => n5228, Q => 
                           n6866, QN => n4839);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1843, CK => n5231, Q => 
                           n6867, QN => n4840);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1842, CK => n5234, Q => 
                           n6868, QN => n4841);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1841, CK => n5237, Q => 
                           n6869, QN => n4842);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1840, CK => n5240, Q => 
                           n6870, QN => n4843);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1839, CK => n5243, Q => 
                           n6871, QN => n4844);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1838, CK => n5247, Q => 
                           n6872, QN => n4845);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1837, CK => n5250, Q => 
                           n6873, QN => n4846);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1836, CK => n5253, Q => 
                           n6874, QN => n4847);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1835, CK => n5256, Q => 
                           n6875, QN => n4848);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1834, CK => n5259, Q => 
                           n6876, QN => n4849);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1833, CK => n5262, Q => 
                           n6877, QN => n4850);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1832, CK => n5265, Q => 
                           n6878, QN => n4851);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1831, CK => n5268, Q => 
                           n6879, QN => n4852);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1830, CK => n5271, Q => 
                           n6880, QN => n4853);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1829, CK => n5274, Q => 
                           n6881, QN => n4854);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1828, CK => n5277, Q => 
                           n6882, QN => n4855);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1827, CK => n5281, Q => 
                           n6883, QN => n4856);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1826, CK => n5284, Q => 
                           n6884, QN => n4857);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1825, CK => n5203, Q => 
                           n6885, QN => n4858);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1824, CK => n5206, Q => 
                           n6886, QN => n4859);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1823, CK => n5209, Q => 
                           n6887, QN => n4860);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1822, CK => n5213, Q => 
                           n6888, QN => n4861);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1821, CK => n5216, Q => 
                           n6889, QN => n4862);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1820, CK => n5219, Q => 
                           n6890, QN => n4863);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1819, CK => n5222, Q => 
                           n6891, QN => n4864);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1818, CK => n5197, Q => 
                           n6892, QN => n4865);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1817, CK => n5200, Q => 
                           n6893, QN => n4866);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1816, CK => n5290, Q => 
                           n6894, QN => n4867);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1815, CK => n5293, Q => 
                           n6895, QN => n4868);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1814, CK => n5287, Q => 
                           n7087, QN => n5093);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1813, CK => n5225, Q => 
                           n7086, QN => n5094);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1812, CK => n5228, Q => 
                           n7085, QN => n5095);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1811, CK => n5231, Q => 
                           n7084, QN => n5096);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1810, CK => n5234, Q => 
                           n7083, QN => n5097);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1809, CK => n5237, Q => 
                           n7082, QN => n5098);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1808, CK => n5240, Q => 
                           n7081, QN => n5099);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1807, CK => n5244, Q => 
                           n7080, QN => n5100);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1806, CK => n5247, Q => 
                           n7079, QN => n5101);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1805, CK => n5250, Q => 
                           n7078, QN => n5102);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1804, CK => n5253, Q => 
                           n7077, QN => n5103);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1803, CK => n5256, Q => 
                           n7076, QN => n5104);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1802, CK => n5259, Q => 
                           n7075, QN => n5105);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1801, CK => n5262, Q => 
                           n7074, QN => n5106);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1800, CK => n5265, Q => 
                           n7073, QN => n5107);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1799, CK => n5268, Q => 
                           n7072, QN => n5108);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1798, CK => n5271, Q => 
                           n7071, QN => n5109);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1797, CK => n5274, Q => 
                           n7070, QN => n5110);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1796, CK => n5278, Q => 
                           n7069, QN => n5111);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1795, CK => n5281, Q => 
                           n7068, QN => n5112);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1794, CK => n5284, Q => 
                           n7067, QN => n5113);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1793, CK => n5203, Q => 
                           n7066, QN => n5114);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1792, CK => n5206, Q => 
                           n7065, QN => n5115);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1791, CK => n5210, Q => 
                           n7064, QN => n5116);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1790, CK => n5213, Q => 
                           n7063, QN => n5117);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1789, CK => n5216, Q => 
                           n7062, QN => n5118);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1788, CK => n5219, Q => 
                           n7061, QN => n5119);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1787, CK => n5222, Q => 
                           n7060, QN => n5120);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1786, CK => n5197, Q => 
                           n7059, QN => n5121);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1785, CK => n5200, Q => 
                           n7058, QN => n5122);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1784, CK => n5290, Q => 
                           n7057, QN => n5123);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1783, CK => n5293, Q => 
                           n7056, QN => n5124);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1782, CK => n5287, Q => 
                           n_1692, QN => n4517);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1781, CK => n5225, Q => 
                           n_1693, QN => n4518);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1780, CK => n5228, Q => 
                           n_1694, QN => n4519);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1779, CK => n5231, Q => 
                           n_1695, QN => n4520);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1778, CK => n5234, Q => 
                           n_1696, QN => n4521);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1777, CK => n5237, Q => 
                           n_1697, QN => n4522);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1776, CK => n5241, Q => 
                           n_1698, QN => n4523);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1775, CK => n5244, Q => 
                           n_1699, QN => n4524);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1774, CK => n5247, Q => 
                           n_1700, QN => n4525);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1773, CK => n5250, Q => 
                           n_1701, QN => n4526);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1772, CK => n5253, Q => 
                           n_1702, QN => n4527);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1771, CK => n5256, Q => 
                           n_1703, QN => n4528);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1770, CK => n5259, Q => 
                           n_1704, QN => n4529);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1769, CK => n5262, Q => 
                           n_1705, QN => n4530);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1768, CK => n5265, Q => 
                           n_1706, QN => n4531);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1767, CK => n5268, Q => 
                           n_1707, QN => n4532);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1766, CK => n5271, Q => 
                           n_1708, QN => n4533);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1765, CK => n5275, Q => 
                           n_1709, QN => n4534);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1764, CK => n5278, Q => 
                           n_1710, QN => n4535);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1763, CK => n5281, Q => 
                           n_1711, QN => n4536);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1762, CK => n5284, Q => 
                           n_1712, QN => n4537);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1761, CK => n5203, Q => 
                           n_1713, QN => n4538);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1760, CK => n5207, Q => 
                           n_1714, QN => n4539);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1759, CK => n5210, Q => 
                           n_1715, QN => n4540);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1758, CK => n5213, Q => 
                           n_1716, QN => n4541);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1757, CK => n5216, Q => 
                           n_1717, QN => n4542);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1756, CK => n5219, Q => 
                           n_1718, QN => n4543);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1755, CK => n5222, Q => 
                           n_1719, QN => n4544);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1754, CK => n5197, Q => 
                           n_1720, QN => n4545);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1753, CK => n5200, Q => 
                           n_1721, QN => n4546);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1752, CK => n5290, Q => 
                           n_1722, QN => n4547);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1751, CK => n5293, Q => 
                           n_1723, QN => n4548);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1750, CK => n5287, Q => 
                           n7055, QN => n5125);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1749, CK => n5225, Q => 
                           n7054, QN => n5126);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1748, CK => n5228, Q => 
                           n7053, QN => n5127);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1747, CK => n5231, Q => 
                           n7052, QN => n5128);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1746, CK => n5234, Q => 
                           n7051, QN => n5129);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1745, CK => n5238, Q => 
                           n7050, QN => n5130);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1744, CK => n5241, Q => 
                           n7049, QN => n5131);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1743, CK => n5244, Q => 
                           n7048, QN => n5132);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1742, CK => n5247, Q => 
                           n7047, QN => n5133);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1741, CK => n5250, Q => 
                           n7046, QN => n5134);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1740, CK => n5253, Q => 
                           n7045, QN => n5135);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1739, CK => n5256, Q => 
                           n7044, QN => n5136);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1738, CK => n5259, Q => 
                           n7043, QN => n5137);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1737, CK => n5262, Q => 
                           n7042, QN => n5138);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1736, CK => n5265, Q => 
                           n7041, QN => n5139);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1735, CK => n5268, Q => 
                           n7040, QN => n5140);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1734, CK => n5272, Q => 
                           n7039, QN => n5141);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1733, CK => n5275, Q => 
                           n7038, QN => n5142);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1732, CK => n5278, Q => 
                           n7037, QN => n5143);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1731, CK => n5281, Q => 
                           n7036, QN => n5144);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1730, CK => n5284, Q => 
                           n7035, QN => n5145);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1729, CK => n5204, Q => 
                           n7034, QN => n5146);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1728, CK => n5207, Q => 
                           n7033, QN => n5147);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1727, CK => n5210, Q => 
                           n7032, QN => n5148);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1726, CK => n5213, Q => 
                           n7031, QN => n5149);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1725, CK => n5216, Q => 
                           n7030, QN => n5150);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1724, CK => n5219, Q => 
                           n7029, QN => n5151);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1723, CK => n5222, Q => 
                           n7028, QN => n5152);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1722, CK => n5197, Q => 
                           n7027, QN => n5153);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1721, CK => n5201, Q => 
                           n7026, QN => n5154);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1720, CK => n5290, Q => 
                           n7025, QN => n5155);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1719, CK => n5293, Q => 
                           n7024, QN => n5156);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1718, CK => n5287, Q => 
                           n6896, QN => n4869);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1717, CK => n5225, Q => 
                           n6897, QN => n4870);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1716, CK => n5228, Q => 
                           n6898, QN => n4871);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1715, CK => n5231, Q => 
                           n6899, QN => n4872);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1714, CK => n5235, Q => 
                           n6900, QN => n4873);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1713, CK => n5238, Q => 
                           n6901, QN => n4874);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1712, CK => n5241, Q => 
                           n6902, QN => n4875);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1711, CK => n5244, Q => 
                           n6903, QN => n4876);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1710, CK => n5247, Q => 
                           n6904, QN => n4877);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1709, CK => n5250, Q => 
                           n6905, QN => n4878);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1708, CK => n5253, Q => 
                           n6906, QN => n4879);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1707, CK => n5256, Q => 
                           n6907, QN => n4880);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1706, CK => n5259, Q => 
                           n6908, QN => n4881);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1705, CK => n5262, Q => 
                           n6909, QN => n4882);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1704, CK => n5265, Q => 
                           n6910, QN => n4883);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1703, CK => n5269, Q => 
                           n6911, QN => n4884);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1702, CK => n5272, Q => 
                           n6912, QN => n4885);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1701, CK => n5275, Q => 
                           n6913, QN => n4886);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1700, CK => n5278, Q => 
                           n6914, QN => n4887);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1699, CK => n5281, Q => 
                           n6915, QN => n4888);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1698, CK => n5284, Q => 
                           n6916, QN => n4889);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1697, CK => n5204, Q => 
                           n6917, QN => n4890);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1696, CK => n5207, Q => 
                           n6918, QN => n4891);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1695, CK => n5210, Q => 
                           n6919, QN => n4892);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1694, CK => n5213, Q => 
                           n6920, QN => n4893);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1693, CK => n5216, Q => 
                           n6921, QN => n4894);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1692, CK => n5219, Q => 
                           n6922, QN => n4895);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1691, CK => n5222, Q => 
                           n6923, QN => n4896);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1690, CK => n5198, Q => 
                           n6924, QN => n4897);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1689, CK => n5201, Q => 
                           n6925, QN => n4898);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1688, CK => n5290, Q => 
                           n6926, QN => n4899);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1687, CK => n5293, Q => 
                           n6927, QN => n4900);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1686, CK => n5287, Q => 
                           n_1724, QN => n4259);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1685, CK => n5225, Q => 
                           n_1725, QN => n4260);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1684, CK => n5228, Q => 
                           n_1726, QN => n4261);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1683, CK => n5232, Q => 
                           n_1727, QN => n4262);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1682, CK => n5235, Q => 
                           n_1728, QN => n4263);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1681, CK => n5238, Q => 
                           n_1729, QN => n4264);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1680, CK => n5241, Q => 
                           n_1730, QN => n4265);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1679, CK => n5244, Q => 
                           n_1731, QN => n4266);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1678, CK => n5247, Q => 
                           n_1732, QN => n4267);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1677, CK => n5250, Q => 
                           n_1733, QN => n4268);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1676, CK => n5253, Q => 
                           n_1734, QN => n4269);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1675, CK => n5256, Q => 
                           n_1735, QN => n4270);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1674, CK => n5259, Q => 
                           n_1736, QN => n4271);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1673, CK => n5262, Q => 
                           n_1737, QN => n4272);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1672, CK => n5266, Q => 
                           n_1738, QN => n4273);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1671, CK => n5269, Q => 
                           n_1739, QN => n4274);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1670, CK => n5272, Q => 
                           n_1740, QN => n4275);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1669, CK => n5275, Q => 
                           n_1741, QN => n4276);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1668, CK => n5278, Q => 
                           n_1742, QN => n4277);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1667, CK => n5281, Q => 
                           n_1743, QN => n4278);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1666, CK => n5284, Q => 
                           n_1744, QN => n4279);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1665, CK => n5204, Q => 
                           n_1745, QN => n4280);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1664, CK => n5207, Q => 
                           n_1746, QN => n4281);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1663, CK => n5210, Q => 
                           n_1747, QN => n4282);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1662, CK => n5213, Q => 
                           n_1748, QN => n4283);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1661, CK => n5216, Q => 
                           n_1749, QN => n4284);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1660, CK => n5219, Q => 
                           n_1750, QN => n4285);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1659, CK => n5222, Q => 
                           n_1751, QN => n4286);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1658, CK => n5198, Q => 
                           n_1752, QN => n4287);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1657, CK => n5201, Q => 
                           n_1753, QN => n4288);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1656, CK => n5290, Q => 
                           n_1754, QN => n4289);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1655, CK => n5293, Q => 
                           n_1755, QN => n4290);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1654, CK => n5287, Q => 
                           n_1756, QN => n4291);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1653, CK => n5225, Q => 
                           n_1757, QN => n4292);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1652, CK => n5229, Q => 
                           n_1758, QN => n4293);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1651, CK => n5232, Q => 
                           n_1759, QN => n4294);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1650, CK => n5235, Q => 
                           n_1760, QN => n4295);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1649, CK => n5238, Q => 
                           n_1761, QN => n4296);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1648, CK => n5241, Q => 
                           n_1762, QN => n4297);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1647, CK => n5244, Q => 
                           n_1763, QN => n4298);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1646, CK => n5247, Q => 
                           n_1764, QN => n4299);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1645, CK => n5250, Q => 
                           n_1765, QN => n4300);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1644, CK => n5253, Q => 
                           n_1766, QN => n4301);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1643, CK => n5256, Q => 
                           n_1767, QN => n4302);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1642, CK => n5259, Q => 
                           n_1768, QN => n4303);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1641, CK => n5263, Q => 
                           n_1769, QN => n4304);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1640, CK => n5266, Q => 
                           n_1770, QN => n4305);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1639, CK => n5269, Q => 
                           n_1771, QN => n4306);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1638, CK => n5272, Q => 
                           n_1772, QN => n4307);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1637, CK => n5275, Q => 
                           n_1773, QN => n4308);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1636, CK => n5278, Q => 
                           n_1774, QN => n4309);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1635, CK => n5281, Q => 
                           n_1775, QN => n4310);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1634, CK => n5284, Q => 
                           n_1776, QN => n4311);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1633, CK => n5204, Q => 
                           n_1777, QN => n4312);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1632, CK => n5207, Q => 
                           n_1778, QN => n4313);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1631, CK => n5210, Q => 
                           n_1779, QN => n4314);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1630, CK => n5213, Q => 
                           n_1780, QN => n4315);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1629, CK => n5216, Q => 
                           n_1781, QN => n4316);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1628, CK => n5219, Q => 
                           n_1782, QN => n4317);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1627, CK => n5222, Q => 
                           n_1783, QN => n4318);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1626, CK => n5198, Q => 
                           n_1784, QN => n4319);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1625, CK => n5201, Q => 
                           n_1785, QN => n4320);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1624, CK => n5290, Q => 
                           n_1786, QN => n4321);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1623, CK => n5293, Q => 
                           n_1787, QN => n4322);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1622, CK => n5287, Q => 
                           n7023, QN => n4901);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1621, CK => n5226, Q => 
                           n7022, QN => n4902);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1620, CK => n5229, Q => 
                           n7021, QN => n4903);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1619, CK => n5232, Q => 
                           n7020, QN => n4904);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1618, CK => n5235, Q => 
                           n7019, QN => n4905);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1617, CK => n5238, Q => 
                           n7018, QN => n4906);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1616, CK => n5241, Q => 
                           n7017, QN => n4907);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1615, CK => n5244, Q => 
                           n7016, QN => n4908);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1614, CK => n5247, Q => 
                           n7015, QN => n4909);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1613, CK => n5250, Q => 
                           n7014, QN => n4910);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1612, CK => n5253, Q => 
                           n7013, QN => n4911);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1611, CK => n5256, Q => 
                           n7012, QN => n4912);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1610, CK => n5260, Q => 
                           n7011, QN => n4913);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1609, CK => n5263, Q => 
                           n7010, QN => n4914);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1608, CK => n5266, Q => 
                           n7009, QN => n4915);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1607, CK => n5269, Q => 
                           n7008, QN => n4916);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1606, CK => n5272, Q => 
                           n7007, QN => n4917);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1605, CK => n5275, Q => 
                           n7006, QN => n4918);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1604, CK => n5278, Q => 
                           n7005, QN => n4919);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1603, CK => n5281, Q => 
                           n7004, QN => n4920);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1602, CK => n5284, Q => 
                           n7003, QN => n4921);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1601, CK => n5204, Q => 
                           n7002, QN => n4922);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1600, CK => n5207, Q => 
                           n7001, QN => n4923);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1599, CK => n5210, Q => 
                           n7000, QN => n4924);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1598, CK => n5213, Q => 
                           n6999, QN => n4925);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1597, CK => n5216, Q => 
                           n6998, QN => n4926);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1596, CK => n5219, Q => 
                           n6997, QN => n4927);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1595, CK => n5222, Q => 
                           n6996, QN => n4928);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1594, CK => n5198, Q => 
                           n6995, QN => n4929);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1593, CK => n5201, Q => 
                           n6994, QN => n4930);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1592, CK => n5290, Q => 
                           n6993, QN => n4931);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1591, CK => n5294, Q => 
                           n6992, QN => n4932);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1590, CK => n5287, Q => 
                           n_1788, QN => n4549);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1589, CK => n5226, Q => 
                           n_1789, QN => n4550);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1588, CK => n5229, Q => 
                           n_1790, QN => n4551);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1587, CK => n5232, Q => 
                           n_1791, QN => n4552);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1586, CK => n5235, Q => 
                           n_1792, QN => n4553);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1585, CK => n5238, Q => 
                           n_1793, QN => n4554);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1584, CK => n5241, Q => 
                           n_1794, QN => n4555);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1583, CK => n5244, Q => 
                           n_1795, QN => n4556);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1582, CK => n5247, Q => 
                           n_1796, QN => n4557);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1581, CK => n5250, Q => 
                           n_1797, QN => n4558);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1580, CK => n5253, Q => 
                           n_1798, QN => n4559);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1579, CK => n5257, Q => 
                           n_1799, QN => n4560);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1578, CK => n5260, Q => 
                           n_1800, QN => n4561);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1577, CK => n5263, Q => 
                           n_1801, QN => n4562);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1576, CK => n5266, Q => 
                           n_1802, QN => n4563);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1575, CK => n5269, Q => 
                           n_1803, QN => n4564);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1574, CK => n5272, Q => 
                           n_1804, QN => n4565);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1573, CK => n5275, Q => 
                           n_1805, QN => n4566);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1572, CK => n5278, Q => 
                           n_1806, QN => n4567);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1571, CK => n5281, Q => 
                           n_1807, QN => n4568);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1570, CK => n5284, Q => 
                           n_1808, QN => n4569);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1569, CK => n5204, Q => 
                           n_1809, QN => n4570);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1568, CK => n5207, Q => 
                           n_1810, QN => n4571);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1567, CK => n5210, Q => 
                           n_1811, QN => n4572);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1566, CK => n5213, Q => 
                           n_1812, QN => n4573);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1565, CK => n5216, Q => 
                           n_1813, QN => n4574);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1564, CK => n5219, Q => 
                           n_1814, QN => n4575);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1563, CK => n5223, Q => 
                           n_1815, QN => n4576);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1562, CK => n5198, Q => 
                           n_1816, QN => n4577);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1561, CK => n5201, Q => 
                           n_1817, QN => n4578);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1560, CK => n5291, Q => 
                           n_1818, QN => n4579);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1559, CK => n5294, Q => 
                           n_1819, QN => n4580);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1558, CK => n5288, Q => 
                           n_1820, QN => n4581);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1557, CK => n5226, Q => 
                           n_1821, QN => n4582);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1556, CK => n5229, Q => 
                           n_1822, QN => n4583);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1555, CK => n5232, Q => 
                           n_1823, QN => n4584);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1554, CK => n5235, Q => 
                           n_1824, QN => n4585);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1553, CK => n5238, Q => 
                           n_1825, QN => n4586);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1552, CK => n5241, Q => 
                           n_1826, QN => n4587);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1551, CK => n5244, Q => 
                           n_1827, QN => n4588);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1550, CK => n5247, Q => 
                           n_1828, QN => n4589);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1549, CK => n5250, Q => 
                           n_1829, QN => n4590);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1548, CK => n5254, Q => 
                           n_1830, QN => n4591);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1547, CK => n5257, Q => 
                           n_1831, QN => n4592);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1546, CK => n5260, Q => 
                           n_1832, QN => n4593);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1545, CK => n5263, Q => 
                           n_1833, QN => n4594);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1544, CK => n5266, Q => 
                           n_1834, QN => n4595);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1543, CK => n5269, Q => 
                           n_1835, QN => n4596);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1542, CK => n5272, Q => 
                           n_1836, QN => n4597);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1541, CK => n5275, Q => 
                           n_1837, QN => n4598);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1540, CK => n5278, Q => 
                           n_1838, QN => n4599);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1539, CK => n5281, Q => 
                           n_1839, QN => n4600);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1538, CK => n5284, Q => 
                           n_1840, QN => n4601);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1537, CK => n5204, Q => 
                           n_1841, QN => n4602);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1536, CK => n5207, Q => 
                           n_1842, QN => n4603);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1535, CK => n5210, Q => 
                           n_1843, QN => n4604);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1534, CK => n5213, Q => 
                           n_1844, QN => n4605);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1533, CK => n5216, Q => 
                           n_1845, QN => n4606);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1532, CK => n5220, Q => 
                           n_1846, QN => n4607);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1531, CK => n5223, Q => 
                           n_1847, QN => n4608);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1530, CK => n5198, Q => 
                           n_1848, QN => n4609);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1529, CK => n5201, Q => 
                           n_1849, QN => n4610);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1528, CK => n5291, Q => 
                           n_1850, QN => n4611);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1527, CK => n5294, Q => 
                           n_1851, QN => n4612);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1526, CK => n5288, Q => 
                           n_1852, QN => n4323);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1525, CK => n5226, Q => 
                           n_1853, QN => n4324);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1524, CK => n5229, Q => 
                           n_1854, QN => n4325);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1523, CK => n5232, Q => 
                           n_1855, QN => n4326);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1522, CK => n5235, Q => 
                           n_1856, QN => n4327);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1521, CK => n5238, Q => 
                           n_1857, QN => n4328);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1520, CK => n5241, Q => 
                           n_1858, QN => n4329);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1519, CK => n5244, Q => 
                           n_1859, QN => n4330);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1518, CK => n5247, Q => 
                           n_1860, QN => n4331);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1517, CK => n5251, Q => 
                           n_1861, QN => n4332);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1516, CK => n5254, Q => 
                           n_1862, QN => n4333);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1515, CK => n5257, Q => 
                           n_1863, QN => n4334);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1514, CK => n5260, Q => 
                           n_1864, QN => n4335);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1513, CK => n5263, Q => 
                           n_1865, QN => n4336);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1512, CK => n5266, Q => 
                           n_1866, QN => n4337);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1511, CK => n5269, Q => 
                           n_1867, QN => n4338);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1510, CK => n5272, Q => 
                           n_1868, QN => n4339);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1509, CK => n5275, Q => 
                           n_1869, QN => n4340);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1508, CK => n5278, Q => 
                           n_1870, QN => n4341);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1507, CK => n5281, Q => 
                           n_1871, QN => n4342);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1506, CK => n5285, Q => 
                           n_1872, QN => n4343);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1505, CK => n5204, Q => 
                           n_1873, QN => n4344);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1504, CK => n5207, Q => 
                           n_1874, QN => n4345);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1503, CK => n5210, Q => 
                           n_1875, QN => n4346);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1502, CK => n5213, Q => 
                           n_1876, QN => n4347);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1501, CK => n5217, Q => 
                           n_1877, QN => n4348);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1500, CK => n5220, Q => 
                           n_1878, QN => n4349);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1499, CK => n5223, Q => 
                           n_1879, QN => n4350);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1498, CK => n5198, Q => 
                           n_1880, QN => n4351);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1497, CK => n5201, Q => 
                           n_1881, QN => n4352);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1496, CK => n5291, Q => 
                           n_1882, QN => n4353);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1495, CK => n5294, Q => 
                           n_1883, QN => n4354);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1494, CK => n5288, Q => 
                           n6991, QN => n4933);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1493, CK => n5226, Q => 
                           n6990, QN => n4934);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1492, CK => n5229, Q => 
                           n6989, QN => n4935);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1491, CK => n5232, Q => 
                           n6988, QN => n4936);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1490, CK => n5235, Q => 
                           n6987, QN => n4937);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1489, CK => n5238, Q => 
                           n6986, QN => n4938);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1488, CK => n5241, Q => 
                           n6985, QN => n4939);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1487, CK => n5244, Q => 
                           n6984, QN => n4940);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1486, CK => n5248, Q => 
                           n6983, QN => n4941);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1485, CK => n5251, Q => 
                           n6982, QN => n4942);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1484, CK => n5254, Q => 
                           n6981, QN => n4943);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1483, CK => n5257, Q => 
                           n6980, QN => n4944);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1482, CK => n5260, Q => 
                           n6979, QN => n4945);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1481, CK => n5263, Q => 
                           n6978, QN => n4946);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1480, CK => n5266, Q => 
                           n6977, QN => n4947);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1479, CK => n5269, Q => 
                           n6976, QN => n4948);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1478, CK => n5272, Q => 
                           n6975, QN => n4949);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1477, CK => n5275, Q => 
                           n6974, QN => n4950);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1476, CK => n5278, Q => 
                           n6973, QN => n4951);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1475, CK => n5282, Q => 
                           n6972, QN => n4952);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1474, CK => n5285, Q => 
                           n6971, QN => n4953);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1473, CK => n5204, Q => 
                           n6970, QN => n4954);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1472, CK => n5207, Q => 
                           n6969, QN => n4955);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1471, CK => n5210, Q => 
                           n6968, QN => n4956);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1470, CK => n5214, Q => 
                           n6967, QN => n4957);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1469, CK => n5217, Q => 
                           n6966, QN => n4958);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1468, CK => n5220, Q => 
                           n6965, QN => n4959);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1467, CK => n5223, Q => 
                           n6964, QN => n4960);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1466, CK => n5198, Q => 
                           n6963, QN => n4961);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1465, CK => n5201, Q => 
                           n6962, QN => n4962);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1464, CK => n5291, Q => 
                           n6961, QN => n4963);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1463, CK => n5294, Q => 
                           n6960, QN => n4964);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1462, CK => n5288, Q => 
                           n_1884, QN => n4355);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1461, CK => n5226, Q => 
                           n_1885, QN => n4356);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1460, CK => n5229, Q => 
                           n_1886, QN => n4357);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1459, CK => n5232, Q => 
                           n_1887, QN => n4358);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1458, CK => n5235, Q => 
                           n_1888, QN => n4359);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1457, CK => n5238, Q => 
                           n_1889, QN => n4360);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1456, CK => n5241, Q => 
                           n_1890, QN => n4361);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1455, CK => n5245, Q => 
                           n_1891, QN => n4362);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1454, CK => n5248, Q => 
                           n_1892, QN => n4363);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1453, CK => n5251, Q => 
                           n_1893, QN => n4364);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1452, CK => n5254, Q => 
                           n_1894, QN => n4365);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1451, CK => n5257, Q => 
                           n_1895, QN => n4366);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1450, CK => n5260, Q => 
                           n_1896, QN => n4367);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1449, CK => n5263, Q => 
                           n_1897, QN => n4368);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1448, CK => n5266, Q => 
                           n_1898, QN => n4369);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1447, CK => n5269, Q => 
                           n_1899, QN => n4370);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1446, CK => n5272, Q => 
                           n_1900, QN => n4371);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1445, CK => n5275, Q => 
                           n_1901, QN => n4372);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1444, CK => n5279, Q => 
                           n_1902, QN => n4373);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1443, CK => n5282, Q => 
                           n_1903, QN => n4374);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1442, CK => n5285, Q => 
                           n_1904, QN => n4375);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1441, CK => n5204, Q => 
                           n_1905, QN => n4376);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1440, CK => n5207, Q => 
                           n_1906, QN => n4377);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1439, CK => n5211, Q => 
                           n_1907, QN => n4378);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1438, CK => n5214, Q => 
                           n_1908, QN => n4379);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1437, CK => n5217, Q => 
                           n_1909, QN => n4380);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1436, CK => n5220, Q => 
                           n_1910, QN => n4381);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1435, CK => n5223, Q => 
                           n_1911, QN => n4382);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1434, CK => n5198, Q => 
                           n_1912, QN => n4383);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1433, CK => n5201, Q => 
                           n_1913, QN => n4384);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1432, CK => n5291, Q => 
                           n_1914, QN => n4385);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1431, CK => n5294, Q => 
                           n_1915, QN => n4386);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1430, CK => n5288, Q => 
                           n_1916, QN => n4613);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1429, CK => n5226, Q => 
                           n_1917, QN => n4614);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1428, CK => n5229, Q => 
                           n_1918, QN => n4615);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1427, CK => n5232, Q => 
                           n_1919, QN => n4616);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1426, CK => n5235, Q => 
                           n_1920, QN => n4617);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1425, CK => n5238, Q => 
                           n_1921, QN => n4618);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1424, CK => n5242, Q => 
                           n_1922, QN => n4619);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1423, CK => n5245, Q => 
                           n_1923, QN => n4620);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1422, CK => n5248, Q => 
                           n_1924, QN => n4621);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1421, CK => n5251, Q => 
                           n_1925, QN => n4622);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1420, CK => n5254, Q => 
                           n_1926, QN => n4623);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1419, CK => n5257, Q => 
                           n_1927, QN => n4624);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1418, CK => n5260, Q => 
                           n_1928, QN => n4625);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1417, CK => n5263, Q => 
                           n_1929, QN => n4626);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1416, CK => n5266, Q => 
                           n_1930, QN => n4627);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1415, CK => n5269, Q => 
                           n_1931, QN => n4628);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1414, CK => n5272, Q => 
                           n_1932, QN => n4629);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1413, CK => n5276, Q => 
                           n_1933, QN => n4630);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1412, CK => n5279, Q => 
                           n_1934, QN => n4631);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1411, CK => n5282, Q => 
                           n_1935, QN => n4632);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1410, CK => n5285, Q => 
                           n_1936, QN => n4633);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1409, CK => n5204, Q => 
                           n_1937, QN => n4634);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1408, CK => n5208, Q => 
                           n_1938, QN => n4635);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1407, CK => n5211, Q => 
                           n_1939, QN => n4636);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1406, CK => n5214, Q => 
                           n_1940, QN => n4637);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1405, CK => n5217, Q => 
                           n_1941, QN => n4638);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1404, CK => n5220, Q => 
                           n_1942, QN => n4639);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1403, CK => n5223, Q => 
                           n_1943, QN => n4640);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1402, CK => n5198, Q => 
                           n_1944, QN => n4641);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1401, CK => n5201, Q => 
                           n_1945, QN => n4642);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1400, CK => n5291, Q => 
                           n_1946, QN => n4643);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1399, CK => n5294, Q => 
                           n_1947, QN => n4644);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1398, CK => n5288, Q => 
                           n_1948, QN => n4387);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1397, CK => n5226, Q => 
                           n_1949, QN => n4388);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1396, CK => n5229, Q => 
                           n_1950, QN => n4389);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1395, CK => n5232, Q => 
                           n_1951, QN => n4390);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1394, CK => n5235, Q => 
                           n_1952, QN => n4391);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1393, CK => n5239, Q => 
                           n_1953, QN => n4392);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1392, CK => n5242, Q => 
                           n_1954, QN => n4393);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1391, CK => n5245, Q => 
                           n_1955, QN => n4394);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1390, CK => n5248, Q => 
                           n_1956, QN => n4395);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1389, CK => n5251, Q => 
                           n_1957, QN => n4396);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1388, CK => n5254, Q => 
                           n_1958, QN => n4397);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1387, CK => n5257, Q => 
                           n_1959, QN => n4398);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1386, CK => n5260, Q => 
                           n_1960, QN => n4399);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1385, CK => n5263, Q => 
                           n_1961, QN => n4400);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1384, CK => n5266, Q => 
                           n_1962, QN => n4401);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1383, CK => n5269, Q => 
                           n_1963, QN => n4402);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1382, CK => n5273, Q => 
                           n_1964, QN => n4403);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1381, CK => n5276, Q => 
                           n_1965, QN => n4404);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1380, CK => n5279, Q => 
                           n_1966, QN => n4405);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1379, CK => n5282, Q => 
                           n_1967, QN => n4406);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1378, CK => n5285, Q => 
                           n_1968, QN => n4407);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1377, CK => n5205, Q => 
                           n_1969, QN => n4408);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1376, CK => n5208, Q => 
                           n_1970, QN => n4409);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1375, CK => n5211, Q => 
                           n_1971, QN => n4410);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1374, CK => n5214, Q => 
                           n_1972, QN => n4411);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1373, CK => n5217, Q => 
                           n_1973, QN => n4412);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1372, CK => n5220, Q => 
                           n_1974, QN => n4413);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1371, CK => n5223, Q => 
                           n_1975, QN => n4414);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1370, CK => n5198, Q => 
                           n_1976, QN => n4415);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1369, CK => n5202, Q => 
                           n_1977, QN => n4416);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1368, CK => n5291, Q => 
                           n_1978, QN => n4417);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1367, CK => n5294, Q => 
                           n_1979, QN => n4418);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1366, CK => n5288, Q => 
                           n6959, QN => n5157);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1365, CK => n5226, Q => 
                           n6958, QN => n5158);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1364, CK => n5229, Q => 
                           n6957, QN => n5159);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1363, CK => n5232, Q => 
                           n6956, QN => n5160);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1362, CK => n5236, Q => 
                           n6955, QN => n5161);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1361, CK => n5239, Q => 
                           n6954, QN => n5162);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1360, CK => n5242, Q => 
                           n6953, QN => n5163);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1359, CK => n5245, Q => 
                           n6952, QN => n5164);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1358, CK => n5248, Q => 
                           n6951, QN => n5165);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1357, CK => n5251, Q => 
                           n6950, QN => n5166);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1356, CK => n5254, Q => 
                           n6949, QN => n5167);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1355, CK => n5257, Q => 
                           n6948, QN => n5168);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1354, CK => n5260, Q => 
                           n6947, QN => n5169);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1353, CK => n5263, Q => 
                           n6946, QN => n5170);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1352, CK => n5266, Q => 
                           n6945, QN => n5171);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1351, CK => n5270, Q => 
                           n6944, QN => n5172);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1350, CK => n5273, Q => 
                           n6943, QN => n5173);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1349, CK => n5276, Q => 
                           n6942, QN => n5174);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1348, CK => n5279, Q => 
                           n6941, QN => n5175);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1347, CK => n5282, Q => 
                           n6940, QN => n5176);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1346, CK => n5285, Q => 
                           n6939, QN => n5177);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1345, CK => n5205, Q => 
                           n6938, QN => n5178);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1344, CK => n5208, Q => 
                           n6937, QN => n5179);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1343, CK => n5211, Q => 
                           n6936, QN => n5180);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1342, CK => n5214, Q => 
                           n6935, QN => n5181);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1341, CK => n5217, Q => 
                           n6934, QN => n5182);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1340, CK => n5220, Q => 
                           n6933, QN => n5183);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1339, CK => n5223, Q => 
                           n6932, QN => n5184);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1338, CK => n5199, Q => 
                           n6931, QN => n5185);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1337, CK => n5202, Q => 
                           n6930, QN => n5186);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1336, CK => n5291, Q => 
                           n6929, QN => n5187);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1335, CK => n5294, Q => 
                           n6928, QN => n5188);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1334, CK => n5288, Q => 
                           n_1980, QN => n4645);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1333, CK => n5226, Q => 
                           n_1981, QN => n4646);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1332, CK => n5229, Q => 
                           n_1982, QN => n4647);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1331, CK => n5233, Q => 
                           n_1983, QN => n4648);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1330, CK => n5236, Q => 
                           n_1984, QN => n4649);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1329, CK => n5239, Q => 
                           n_1985, QN => n4650);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1328, CK => n5242, Q => 
                           n_1986, QN => n4651);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1327, CK => n5245, Q => 
                           n_1987, QN => n4652);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1326, CK => n5248, Q => 
                           n_1988, QN => n4653);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1325, CK => n5251, Q => 
                           n_1989, QN => n4654);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1324, CK => n5254, Q => 
                           n_1990, QN => n4655);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1323, CK => n5257, Q => 
                           n_1991, QN => n4656);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1322, CK => n5260, Q => 
                           n_1992, QN => n4657);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1321, CK => n5263, Q => 
                           n_1993, QN => n4658);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1320, CK => n5267, Q => 
                           n_1994, QN => n4659);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1319, CK => n5270, Q => 
                           n_1995, QN => n4660);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1318, CK => n5273, Q => 
                           n_1996, QN => n4661);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1317, CK => n5276, Q => 
                           n_1997, QN => n4662);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1316, CK => n5279, Q => 
                           n_1998, QN => n4663);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1315, CK => n5282, Q => 
                           n_1999, QN => n4664);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1314, CK => n5285, Q => 
                           n_2000, QN => n4665);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1313, CK => n5205, Q => 
                           n_2001, QN => n4666);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1312, CK => n5208, Q => 
                           n_2002, QN => n4667);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1311, CK => n5211, Q => 
                           n_2003, QN => n4668);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1310, CK => n5214, Q => 
                           n_2004, QN => n4669);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1309, CK => n5217, Q => 
                           n_2005, QN => n4670);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1308, CK => n5220, Q => 
                           n_2006, QN => n4671);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1307, CK => n5223, Q => 
                           n_2007, QN => n4672);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1306, CK => n5199, Q => 
                           n_2008, QN => n4673);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1305, CK => n5202, Q => 
                           n_2009, QN => n4674);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1304, CK => n5291, Q => 
                           n_2010, QN => n4675);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1303, CK => n5294, Q => 
                           n_2011, QN => n4676);
   OUT1_reg_31_inst : DFF_X1 port map( D => n4162, CK => n5285, Q => 
                           OUT1_31_port, QN => n_2012);
   OUT1_reg_30_inst : DFF_X1 port map( D => n4161, CK => n5223, Q => 
                           OUT1_30_port, QN => n_2013);
   OUT1_reg_29_inst : DFF_X1 port map( D => n4160, CK => n5226, Q => 
                           OUT1_29_port, QN => n_2014);
   OUT1_reg_28_inst : DFF_X1 port map( D => n4159, CK => n5230, Q => 
                           OUT1_28_port, QN => n_2015);
   OUT1_reg_27_inst : DFF_X1 port map( D => n4158, CK => n5233, Q => 
                           OUT1_27_port, QN => n_2016);
   OUT1_reg_26_inst : DFF_X1 port map( D => n4157, CK => n5236, Q => 
                           OUT1_26_port, QN => n_2017);
   OUT1_reg_25_inst : DFF_X1 port map( D => n4156, CK => n5239, Q => 
                           OUT1_25_port, QN => n_2018);
   OUT1_reg_24_inst : DFF_X1 port map( D => n4155, CK => n5242, Q => 
                           OUT1_24_port, QN => n_2019);
   OUT1_reg_23_inst : DFF_X1 port map( D => n4154, CK => n5245, Q => 
                           OUT1_23_port, QN => n_2020);
   OUT1_reg_22_inst : DFF_X1 port map( D => n4153, CK => n5248, Q => 
                           OUT1_22_port, QN => n_2021);
   OUT1_reg_21_inst : DFF_X1 port map( D => n4152, CK => n5251, Q => 
                           OUT1_21_port, QN => n_2022);
   OUT1_reg_20_inst : DFF_X1 port map( D => n4151, CK => n5254, Q => 
                           OUT1_20_port, QN => n_2023);
   OUT1_reg_19_inst : DFF_X1 port map( D => n4150, CK => n5257, Q => 
                           OUT1_19_port, QN => n_2024);
   OUT1_reg_18_inst : DFF_X1 port map( D => n4149, CK => n5260, Q => 
                           OUT1_18_port, QN => n_2025);
   OUT1_reg_17_inst : DFF_X1 port map( D => n4148, CK => n5264, Q => 
                           OUT1_17_port, QN => n_2026);
   OUT1_reg_16_inst : DFF_X1 port map( D => n4147, CK => n5267, Q => 
                           OUT1_16_port, QN => n_2027);
   OUT1_reg_15_inst : DFF_X1 port map( D => n4146, CK => n5270, Q => 
                           OUT1_15_port, QN => n_2028);
   OUT1_reg_14_inst : DFF_X1 port map( D => n4145, CK => n5273, Q => 
                           OUT1_14_port, QN => n_2029);
   OUT1_reg_13_inst : DFF_X1 port map( D => n4144, CK => n5276, Q => 
                           OUT1_13_port, QN => n_2030);
   OUT1_reg_12_inst : DFF_X1 port map( D => n4143, CK => n5279, Q => 
                           OUT1_12_port, QN => n_2031);
   OUT1_reg_11_inst : DFF_X1 port map( D => n4142, CK => n5282, Q => 
                           OUT1_11_port, QN => n_2032);
   OUT1_reg_10_inst : DFF_X1 port map( D => n4141, CK => n5196, Q => 
                           OUT1_10_port, QN => n_2033);
   OUT1_reg_9_inst : DFF_X1 port map( D => n4140, CK => n5205, Q => OUT1_9_port
                           , QN => n_2034);
   OUT1_reg_8_inst : DFF_X1 port map( D => n4139, CK => n5208, Q => OUT1_8_port
                           , QN => n_2035);
   OUT1_reg_7_inst : DFF_X1 port map( D => n4138, CK => n5211, Q => OUT1_7_port
                           , QN => n_2036);
   OUT1_reg_6_inst : DFF_X1 port map( D => n4137, CK => n5214, Q => OUT1_6_port
                           , QN => n_2037);
   OUT1_reg_5_inst : DFF_X1 port map( D => n4136, CK => n5217, Q => OUT1_5_port
                           , QN => n_2038);
   OUT1_reg_4_inst : DFF_X1 port map( D => n4135, CK => n5220, Q => OUT1_4_port
                           , QN => n_2039);
   OUT1_reg_3_inst : DFF_X1 port map( D => n4134, CK => n5196, Q => OUT1_3_port
                           , QN => n_2040);
   OUT1_reg_2_inst : DFF_X1 port map( D => n4133, CK => n5199, Q => OUT1_2_port
                           , QN => n_2041);
   OUT1_reg_1_inst : DFF_X1 port map( D => n4132, CK => n5288, Q => OUT1_1_port
                           , QN => n_2042);
   OUT1_reg_0_inst : DFF_X1 port map( D => n4131, CK => n5291, Q => OUT1_0_port
                           , QN => n_2043);
   U3 : OR2_X1 port map( A1 => n5195, A2 => n5358, ZN => n4483);
   U4 : OR2_X1 port map( A1 => n5195, A2 => n5952, ZN => n4484);
   U5 : NAND2_X2 port map( A1 => n5192, A2 => n6563, ZN => n6564);
   U6 : NAND2_X2 port map( A1 => n5193, A2 => n6566, ZN => n6567);
   U7 : NAND2_X2 port map( A1 => n5192, A2 => n6572, ZN => n6573);
   U8 : NAND2_X2 port map( A1 => n5193, A2 => n6575, ZN => n6576);
   U9 : NAND2_X2 port map( A1 => n5192, A2 => n6578, ZN => n6579);
   U10 : NAND2_X2 port map( A1 => n5193, A2 => n6581, ZN => n6582);
   U11 : NAND2_X2 port map( A1 => n5193, A2 => n6590, ZN => n6591);
   U12 : NAND2_X2 port map( A1 => n5193, A2 => n6592, ZN => n6593);
   U13 : NAND2_X2 port map( A1 => n5193, A2 => n6598, ZN => n6599);
   U14 : NAND2_X2 port map( A1 => n5192, A2 => n6613, ZN => n6614);
   U15 : NAND2_X2 port map( A1 => n5192, A2 => n6615, ZN => n6616);
   U16 : NAND2_X2 port map( A1 => n5192, A2 => n6619, ZN => n6620);
   U17 : INV_X2 port map( A => n4483, ZN => n5189);
   U18 : INV_X2 port map( A => n4484, ZN => n5190);
   U19 : NAND2_X2 port map( A1 => n5193, A2 => n6600, ZN => n6601);
   U20 : NAND2_X2 port map( A1 => n5192, A2 => n6621, ZN => n6622);
   U21 : NAND2_X2 port map( A1 => n6589, A2 => n6565, ZN => n6590);
   U22 : AND2_X2 port map( A1 => n6519, A2 => n6501, ZN => n5967);
   U23 : AND2_X2 port map( A1 => n6505, A2 => n6507, ZN => n5947);
   U24 : AND2_X2 port map( A1 => n6518, A2 => n6498, ZN => n5978);
   U25 : NAND2_X2 port map( A1 => n5924, A2 => n5908, ZN => n5381);
   U26 : NAND2_X2 port map( A1 => n5925, A2 => n5910, ZN => n5370);
   U27 : AND2_X2 port map( A1 => n5911, A2 => n5913, ZN => n5353);
   U28 : NAND2_X2 port map( A1 => n5193, A2 => n6607, ZN => n6608);
   U29 : NAND2_X2 port map( A1 => n5192, A2 => n6624, ZN => n6625);
   U30 : NAND2_X2 port map( A1 => n6577, A2 => n6562, ZN => n6575);
   U31 : NAND2_X2 port map( A1 => n6606, A2 => n6565, ZN => n6607);
   U32 : NAND2_X2 port map( A1 => n6623, A2 => n6561, ZN => n6621);
   U33 : AND2_X2 port map( A1 => n6519, A2 => n6506, ZN => n5961);
   U34 : AND2_X2 port map( A1 => n6518, A2 => n6508, ZN => n5972);
   U35 : NAND2_X2 port map( A1 => n6505, A2 => n6498, ZN => n5955);
   U36 : AND2_X2 port map( A1 => n5925, A2 => n5912, ZN => n5367);
   U37 : AND2_X2 port map( A1 => n5924, A2 => n5904, ZN => n5384);
   U38 : NAND2_X2 port map( A1 => n5192, A2 => n6630, ZN => n6631);
   U39 : NAND2_X2 port map( A1 => n5193, A2 => n6587, ZN => n6588);
   U40 : NAND2_X2 port map( A1 => n5911, A2 => n5914, ZN => n5362);
   U41 : NAND2_X2 port map( A1 => n6580, A2 => n6562, ZN => n6578);
   U42 : NAND2_X2 port map( A1 => n6589, A2 => n6577, ZN => n6598);
   U43 : NAND2_X2 port map( A1 => n6606, A2 => n6574, ZN => n6613);
   U44 : NAND2_X2 port map( A1 => n6623, A2 => n6565, ZN => n6624);
   U45 : AND2_X2 port map( A1 => n6508, A2 => n6499, ZN => n5942);
   U46 : NAND2_X2 port map( A1 => n6518, A2 => n6506, ZN => n5966);
   U47 : NAND2_X2 port map( A1 => n6519, A2 => n6502, ZN => n5977);
   U48 : NAND2_X2 port map( A1 => n6505, A2 => n6501, ZN => n5950);
   U49 : AND2_X2 port map( A1 => n5908, A2 => n5905, ZN => n5343);
   U50 : AND2_X2 port map( A1 => n5924, A2 => n5914, ZN => n5378);
   U51 : AND2_X2 port map( A1 => n5925, A2 => n5907, ZN => n5373);
   U52 : NAND2_X2 port map( A1 => n5192, A2 => n6632, ZN => n6633);
   U53 : NAND2_X2 port map( A1 => n5193, A2 => n6594, ZN => n6595);
   U54 : NAND2_X2 port map( A1 => n5911, A2 => n5906, ZN => n5357);
   U55 : NAND2_X2 port map( A1 => n6583, A2 => n6562, ZN => n6581);
   U56 : NAND2_X2 port map( A1 => n6589, A2 => n6568, ZN => n6592);
   U57 : NAND2_X2 port map( A1 => n6606, A2 => n6577, ZN => n6615);
   U58 : NAND2_X2 port map( A1 => n6623, A2 => n6571, ZN => n6630);
   U59 : AND2_X2 port map( A1 => n6502, A2 => n6499, ZN => n5937);
   U60 : NAND2_X2 port map( A1 => n6506, A2 => n6505, ZN => n5945);
   U61 : NAND2_X2 port map( A1 => n6518, A2 => n6501, ZN => n5970);
   U62 : AND2_X2 port map( A1 => n5914, A2 => n5905, ZN => n5348);
   U63 : AND2_X2 port map( A1 => n6519, A2 => n6498, ZN => n5979);
   U64 : NAND2_X2 port map( A1 => n5924, A2 => n5912, ZN => n5372);
   U65 : NAND2_X2 port map( A1 => n5192, A2 => n6634, ZN => n6635);
   U66 : NAND2_X2 port map( A1 => n5193, A2 => n6596, ZN => n6597);
   U67 : NAND2_X2 port map( A1 => n5925, A2 => n5913, ZN => n5382);
   U68 : NAND2_X2 port map( A1 => n5910, A2 => n5911, ZN => n5352);
   U69 : NAND2_X2 port map( A1 => n6606, A2 => n6583, ZN => n6619);
   U70 : NAND2_X2 port map( A1 => n6623, A2 => n6574, ZN => n6632);
   U71 : NAND2_X2 port map( A1 => n6565, A2 => n6562, ZN => n6563);
   U72 : NAND2_X2 port map( A1 => n6589, A2 => n6561, ZN => n6587);
   U73 : NAND2_X2 port map( A1 => n6500, A2 => n6499, ZN => n5940);
   U74 : AND2_X2 port map( A1 => n6518, A2 => n6507, ZN => n5968);
   U75 : AND2_X2 port map( A1 => n6505, A2 => n6502, ZN => n5948);
   U76 : NAND2_X2 port map( A1 => n6519, A2 => n6504, ZN => n5964);
   U77 : NAND2_X2 port map( A1 => n5192, A2 => n6638, ZN => n6639);
   U78 : NAND2_X2 port map( A1 => n5193, A2 => n6604, ZN => n6605);
   U79 : NAND2_X2 port map( A1 => n5924, A2 => n5910, ZN => n5371);
   U80 : NAND2_X2 port map( A1 => n5904, A2 => n5905, ZN => n5347);
   U81 : NAND2_X2 port map( A1 => n5925, A2 => n5906, ZN => n5377);
   U82 : AND2_X2 port map( A1 => n5911, A2 => n5908, ZN => n5354);
   U83 : NAND2_X2 port map( A1 => n6589, A2 => n6580, ZN => n6600);
   U84 : NAND2_X2 port map( A1 => n6623, A2 => n6577, ZN => n6634);
   U85 : NAND2_X2 port map( A1 => n6568, A2 => n6562, ZN => n6566);
   U86 : NAND2_X2 port map( A1 => n6606, A2 => n6561, ZN => n6604);
   U87 : AND2_X2 port map( A1 => n6507, A2 => n6499, ZN => n5943);
   U88 : AND2_X2 port map( A1 => n6518, A2 => n6500, ZN => n5962);
   U89 : AND2_X2 port map( A1 => n6519, A2 => n6508, ZN => n5973);
   U90 : NAND2_X2 port map( A1 => n5925, A2 => n5908, ZN => n5383);
   U91 : NAND2_X2 port map( A1 => n6504, A2 => n6505, ZN => n5946);
   U92 : NAND2_X2 port map( A1 => n5193, A2 => n6609, ZN => n6610);
   U93 : NAND2_X2 port map( A1 => n5192, A2 => n6617, ZN => n6618);
   U94 : AND2_X2 port map( A1 => n5924, A2 => n5906, ZN => n5368);
   U95 : AND2_X2 port map( A1 => n5913, A2 => n5905, ZN => n5349);
   U96 : NAND2_X2 port map( A1 => n5911, A2 => n5907, ZN => n5356);
   U97 : NAND2_X2 port map( A1 => n6623, A2 => n6583, ZN => n6638);
   U98 : NAND2_X2 port map( A1 => n6574, A2 => n6562, ZN => n6572);
   U99 : NAND2_X2 port map( A1 => n6589, A2 => n6571, ZN => n6594);
   U100 : NAND2_X2 port map( A1 => n6606, A2 => n6568, ZN => n6609);
   U101 : AND2_X2 port map( A1 => n6501, A2 => n6499, ZN => n5938);
   U102 : NAND2_X2 port map( A1 => n6518, A2 => n6502, ZN => n5975);
   U103 : NAND2_X2 port map( A1 => n6505, A2 => n6508, ZN => n5956);
   U104 : NAND2_X2 port map( A1 => n6504, A2 => n6509, ZN => n5982);
   U105 : NAND2_X2 port map( A1 => n6519, A2 => n6500, ZN => n5971);
   U106 : NAND2_X2 port map( A1 => n5192, A2 => n6569, ZN => n6570);
   U107 : NAND2_X2 port map( A1 => n5193, A2 => n6602, ZN => n6603);
   U108 : NAND2_X2 port map( A1 => n5192, A2 => n6627, ZN => n6628);
   U109 : NAND2_X2 port map( A1 => n5910, A2 => n5915, ZN => n5388);
   U110 : AND2_X2 port map( A1 => n5907, A2 => n5905, ZN => n5344);
   U111 : AND2_X2 port map( A1 => n5925, A2 => n5904, ZN => n5385);
   U112 : AND2_X2 port map( A1 => n5924, A2 => n5913, ZN => n5374);
   U113 : NAND2_X2 port map( A1 => n5912, A2 => n5911, ZN => n5351);
   U114 : NAND2_X2 port map( A1 => n6571, A2 => n6562, ZN => n6569);
   U115 : NAND2_X2 port map( A1 => n6589, A2 => n6574, ZN => n6596);
   U116 : NAND2_X2 port map( A1 => n6606, A2 => n6580, ZN => n6617);
   U117 : NAND2_X2 port map( A1 => n6623, A2 => n6568, ZN => n6627);
   U118 : NAND2_X2 port map( A1 => n6506, A2 => n6509, ZN => n5981);
   U119 : NAND2_X2 port map( A1 => n5193, A2 => n6527, ZN => n6529);
   U120 : NAND2_X2 port map( A1 => n6498, A2 => n6499, ZN => n5941);
   U121 : NAND2_X2 port map( A1 => n6505, A2 => n6500, ZN => n5951);
   U122 : NAND2_X2 port map( A1 => n5193, A2 => n6611, ZN => n6612);
   U123 : NAND2_X2 port map( A1 => n5192, A2 => n6636, ZN => n6637);
   U124 : NAND2_X2 port map( A1 => n6518, A2 => n6504, ZN => n5965);
   U125 : NAND2_X2 port map( A1 => n6519, A2 => n6507, ZN => n5976);
   U126 : INV_X2 port map( A => DATAIN(31), ZN => n6528);
   U127 : INV_X2 port map( A => DATAIN(30), ZN => n6530);
   U128 : INV_X2 port map( A => DATAIN(29), ZN => n6531);
   U129 : INV_X2 port map( A => DATAIN(28), ZN => n6532);
   U130 : INV_X2 port map( A => DATAIN(27), ZN => n6533);
   U131 : INV_X2 port map( A => DATAIN(26), ZN => n6534);
   U132 : INV_X2 port map( A => DATAIN(25), ZN => n6535);
   U133 : INV_X2 port map( A => DATAIN(24), ZN => n6536);
   U134 : INV_X2 port map( A => DATAIN(23), ZN => n6537);
   U135 : INV_X2 port map( A => DATAIN(22), ZN => n6538);
   U136 : INV_X2 port map( A => DATAIN(21), ZN => n6539);
   U137 : INV_X2 port map( A => DATAIN(20), ZN => n6540);
   U138 : INV_X2 port map( A => DATAIN(19), ZN => n6541);
   U139 : INV_X2 port map( A => DATAIN(18), ZN => n6542);
   U140 : INV_X2 port map( A => DATAIN(17), ZN => n6543);
   U141 : INV_X2 port map( A => DATAIN(16), ZN => n6544);
   U142 : INV_X2 port map( A => DATAIN(15), ZN => n6545);
   U143 : INV_X2 port map( A => DATAIN(14), ZN => n6546);
   U144 : INV_X2 port map( A => DATAIN(13), ZN => n6547);
   U145 : INV_X2 port map( A => DATAIN(12), ZN => n6548);
   U146 : INV_X2 port map( A => DATAIN(11), ZN => n6549);
   U147 : INV_X2 port map( A => DATAIN(10), ZN => n6550);
   U148 : INV_X2 port map( A => DATAIN(9), ZN => n6551);
   U149 : INV_X2 port map( A => DATAIN(8), ZN => n6552);
   U150 : INV_X2 port map( A => DATAIN(7), ZN => n6553);
   U151 : INV_X2 port map( A => DATAIN(6), ZN => n6554);
   U152 : INV_X2 port map( A => DATAIN(5), ZN => n6555);
   U153 : INV_X2 port map( A => DATAIN(4), ZN => n6556);
   U154 : INV_X2 port map( A => DATAIN(3), ZN => n6557);
   U155 : INV_X2 port map( A => DATAIN(2), ZN => n6558);
   U156 : INV_X2 port map( A => DATAIN(1), ZN => n6559);
   U157 : INV_X2 port map( A => DATAIN(0), ZN => n6560);
   U158 : AND2_X2 port map( A1 => n5925, A2 => n5914, ZN => n5379);
   U159 : NAND2_X2 port map( A1 => n5911, A2 => n5904, ZN => n5361);
   U160 : NAND2_X2 port map( A1 => n5906, A2 => n5905, ZN => n5346);
   U161 : NAND2_X2 port map( A1 => n5912, A2 => n5915, ZN => n5387);
   U162 : NAND2_X2 port map( A1 => n5924, A2 => n5907, ZN => n5376);
   U163 : NAND2_X2 port map( A1 => n6589, A2 => n6583, ZN => n6602);
   U164 : NAND2_X2 port map( A1 => n6606, A2 => n6571, ZN => n6611);
   U165 : NAND2_X2 port map( A1 => n6623, A2 => n6580, ZN => n6636);
   U166 : NAND2_X2 port map( A1 => n6561, A2 => n6562, ZN => n6527);
   U167 : AND2_X2 port map( A1 => RD2, A2 => ENABLE, ZN => n5952);
   U168 : AND2_X2 port map( A1 => RD1, A2 => ENABLE, ZN => n5358);
   U169 : BUF_X1 port map( A => n5335, Z => n5332);
   U170 : BUF_X1 port map( A => n5336, Z => n5331);
   U171 : BUF_X1 port map( A => n5336, Z => n5330);
   U172 : BUF_X1 port map( A => n5336, Z => n5329);
   U173 : BUF_X1 port map( A => n5335, Z => n5333);
   U174 : BUF_X1 port map( A => n5337, Z => n5328);
   U175 : BUF_X1 port map( A => n5338, Z => n5336);
   U176 : BUF_X1 port map( A => n5338, Z => n5335);
   U177 : BUF_X1 port map( A => n5191, Z => n5194);
   U178 : BUF_X1 port map( A => CLK, Z => n5338);
   U179 : BUF_X1 port map( A => n5306, Z => n5260);
   U180 : BUF_X1 port map( A => n5317, Z => n5226);
   U181 : BUF_X1 port map( A => n5305, Z => n5263);
   U182 : BUF_X1 port map( A => n5316, Z => n5229);
   U183 : BUF_X1 port map( A => n5304, Z => n5266);
   U184 : BUF_X1 port map( A => n5315, Z => n5232);
   U185 : BUF_X1 port map( A => n5303, Z => n5269);
   U186 : BUF_X1 port map( A => n5314, Z => n5235);
   U187 : BUF_X1 port map( A => n5302, Z => n5272);
   U188 : BUF_X1 port map( A => n5313, Z => n5238);
   U189 : BUF_X1 port map( A => n5301, Z => n5275);
   U190 : BUF_X1 port map( A => n5312, Z => n5241);
   U191 : BUF_X1 port map( A => n5300, Z => n5278);
   U192 : BUF_X1 port map( A => n5311, Z => n5244);
   U193 : BUF_X1 port map( A => n5322, Z => n5213);
   U194 : BUF_X1 port map( A => n5299, Z => n5281);
   U195 : BUF_X1 port map( A => n5310, Z => n5247);
   U196 : BUF_X1 port map( A => n5321, Z => n5216);
   U197 : BUF_X1 port map( A => n5298, Z => n5284);
   U198 : BUF_X1 port map( A => n5309, Z => n5250);
   U199 : BUF_X1 port map( A => n5320, Z => n5219);
   U200 : BUF_X1 port map( A => n5308, Z => n5253);
   U201 : BUF_X1 port map( A => n5297, Z => n5287);
   U202 : BUF_X1 port map( A => n5296, Z => n5290);
   U203 : BUF_X1 port map( A => n5319, Z => n5222);
   U204 : BUF_X1 port map( A => n5307, Z => n5256);
   U205 : BUF_X1 port map( A => n5295, Z => n5293);
   U206 : BUF_X1 port map( A => n5306, Z => n5259);
   U207 : BUF_X1 port map( A => n5318, Z => n5225);
   U208 : BUF_X1 port map( A => n5305, Z => n5262);
   U209 : BUF_X1 port map( A => n5317, Z => n5228);
   U210 : BUF_X1 port map( A => n5304, Z => n5265);
   U211 : BUF_X1 port map( A => n5316, Z => n5231);
   U212 : BUF_X1 port map( A => n5303, Z => n5268);
   U213 : BUF_X1 port map( A => n5315, Z => n5234);
   U214 : BUF_X1 port map( A => n5302, Z => n5271);
   U215 : BUF_X1 port map( A => n5314, Z => n5237);
   U216 : BUF_X1 port map( A => n5301, Z => n5274);
   U217 : BUF_X1 port map( A => n5313, Z => n5240);
   U218 : BUF_X1 port map( A => n5300, Z => n5277);
   U219 : BUF_X1 port map( A => n5312, Z => n5243);
   U220 : BUF_X1 port map( A => n5322, Z => n5212);
   U221 : BUF_X1 port map( A => n5299, Z => n5280);
   U222 : BUF_X1 port map( A => n5311, Z => n5246);
   U223 : BUF_X1 port map( A => n5321, Z => n5215);
   U224 : BUF_X1 port map( A => n5298, Z => n5283);
   U225 : BUF_X1 port map( A => n5310, Z => n5249);
   U226 : BUF_X1 port map( A => n5320, Z => n5218);
   U227 : BUF_X1 port map( A => n5309, Z => n5252);
   U228 : BUF_X1 port map( A => n5297, Z => n5286);
   U229 : BUF_X1 port map( A => n5296, Z => n5289);
   U230 : BUF_X1 port map( A => n5319, Z => n5221);
   U231 : BUF_X1 port map( A => n5308, Z => n5255);
   U232 : BUF_X1 port map( A => n5295, Z => n5292);
   U233 : BUF_X1 port map( A => n5307, Z => n5258);
   U234 : BUF_X1 port map( A => n5318, Z => n5224);
   U235 : BUF_X1 port map( A => n5296, Z => n5291);
   U236 : BUF_X1 port map( A => n5297, Z => n5288);
   U237 : BUF_X1 port map( A => n5319, Z => n5220);
   U238 : BUF_X1 port map( A => n5320, Z => n5217);
   U239 : BUF_X1 port map( A => n5321, Z => n5214);
   U240 : BUF_X1 port map( A => n5322, Z => n5211);
   U241 : BUF_X1 port map( A => n5299, Z => n5282);
   U242 : BUF_X1 port map( A => n5300, Z => n5279);
   U243 : BUF_X1 port map( A => n5301, Z => n5276);
   U244 : BUF_X1 port map( A => n5302, Z => n5273);
   U245 : BUF_X1 port map( A => n5303, Z => n5270);
   U246 : BUF_X1 port map( A => n5304, Z => n5267);
   U247 : BUF_X1 port map( A => n5305, Z => n5264);
   U248 : BUF_X1 port map( A => n5306, Z => n5261);
   U249 : BUF_X1 port map( A => n5307, Z => n5257);
   U250 : BUF_X1 port map( A => n5308, Z => n5254);
   U251 : BUF_X1 port map( A => n5309, Z => n5251);
   U252 : BUF_X1 port map( A => n5310, Z => n5248);
   U253 : BUF_X1 port map( A => n5311, Z => n5245);
   U254 : BUF_X1 port map( A => n5312, Z => n5242);
   U255 : BUF_X1 port map( A => n5313, Z => n5239);
   U256 : BUF_X1 port map( A => n5314, Z => n5236);
   U257 : BUF_X1 port map( A => n5315, Z => n5233);
   U258 : BUF_X1 port map( A => n5316, Z => n5230);
   U259 : BUF_X1 port map( A => n5317, Z => n5227);
   U260 : BUF_X1 port map( A => n5318, Z => n5223);
   U261 : BUF_X1 port map( A => n5298, Z => n5285);
   U262 : BUF_X1 port map( A => n5295, Z => n5294);
   U263 : BUF_X1 port map( A => n5329, Z => n5319);
   U264 : BUF_X1 port map( A => n5329, Z => n5320);
   U265 : BUF_X1 port map( A => n5329, Z => n5321);
   U266 : BUF_X1 port map( A => n5329, Z => n5322);
   U267 : BUF_X1 port map( A => n5333, Z => n5299);
   U268 : BUF_X1 port map( A => n5333, Z => n5300);
   U269 : BUF_X1 port map( A => n5333, Z => n5301);
   U270 : BUF_X1 port map( A => n5333, Z => n5302);
   U271 : BUF_X1 port map( A => n5332, Z => n5303);
   U272 : BUF_X1 port map( A => n5332, Z => n5304);
   U273 : BUF_X1 port map( A => n5332, Z => n5305);
   U274 : BUF_X1 port map( A => n5332, Z => n5306);
   U275 : BUF_X1 port map( A => n5332, Z => n5307);
   U276 : BUF_X1 port map( A => n5331, Z => n5308);
   U277 : BUF_X1 port map( A => n5331, Z => n5309);
   U278 : BUF_X1 port map( A => n5331, Z => n5310);
   U279 : BUF_X1 port map( A => n5331, Z => n5311);
   U280 : BUF_X1 port map( A => n5331, Z => n5312);
   U281 : BUF_X1 port map( A => n5330, Z => n5313);
   U282 : BUF_X1 port map( A => n5330, Z => n5314);
   U283 : BUF_X1 port map( A => n5330, Z => n5315);
   U284 : BUF_X1 port map( A => n5330, Z => n5316);
   U285 : BUF_X1 port map( A => n5330, Z => n5317);
   U286 : BUF_X1 port map( A => n5329, Z => n5318);
   U287 : BUF_X1 port map( A => n5333, Z => n5298);
   U288 : BUF_X1 port map( A => n5334, Z => n5295);
   U289 : BUF_X1 port map( A => n5334, Z => n5296);
   U290 : BUF_X1 port map( A => n5334, Z => n5297);
   U291 : BUF_X1 port map( A => n5327, Z => n5198);
   U292 : BUF_X1 port map( A => n5326, Z => n5201);
   U293 : BUF_X1 port map( A => n5325, Z => n5204);
   U294 : BUF_X1 port map( A => n5324, Z => n5207);
   U295 : BUF_X1 port map( A => n5323, Z => n5210);
   U296 : BUF_X1 port map( A => n5327, Z => n5197);
   U297 : BUF_X1 port map( A => n5326, Z => n5200);
   U298 : BUF_X1 port map( A => n5325, Z => n5203);
   U299 : BUF_X1 port map( A => n5324, Z => n5206);
   U300 : BUF_X1 port map( A => n5323, Z => n5209);
   U301 : BUF_X1 port map( A => n5326, Z => n5199);
   U302 : BUF_X1 port map( A => n5327, Z => n5196);
   U303 : BUF_X1 port map( A => n5323, Z => n5208);
   U304 : BUF_X1 port map( A => n5324, Z => n5205);
   U305 : BUF_X1 port map( A => n5325, Z => n5202);
   U306 : BUF_X1 port map( A => n5328, Z => n5326);
   U307 : BUF_X1 port map( A => n5328, Z => n5327);
   U308 : BUF_X1 port map( A => n5328, Z => n5323);
   U309 : BUF_X1 port map( A => n5328, Z => n5324);
   U310 : BUF_X1 port map( A => n5328, Z => n5325);
   U311 : BUF_X1 port map( A => n5335, Z => n5334);
   U312 : INV_X1 port map( A => n5194, ZN => n5192);
   U313 : INV_X1 port map( A => n5194, ZN => n5193);
   U314 : BUF_X1 port map( A => n5338, Z => n5337);
   U315 : BUF_X1 port map( A => n5191, Z => n5195);
   U316 : BUF_X1 port map( A => RESET, Z => n5191);
   U317 : NAND4_X1 port map( A1 => n5339, A2 => n5340, A3 => n5341, A4 => n5342
                           , ZN => n4162);
   U318 : AOI221_X1 port map( B1 => n7023, B2 => n5343, C1 => n7087, C2 => 
                           n5344, A => n5345, ZN => n5342);
   U319 : OAI22_X1 port map( A1 => n5346, A2 => n4517, B1 => n5347, B2 => n4259
                           , ZN => n5345);
   U320 : AOI221_X1 port map( B1 => n6896, B2 => n5348, C1 => n7055, C2 => 
                           n5349, A => n5350, ZN => n5341);
   U321 : OAI22_X1 port map( A1 => n5351, A2 => n4645, B1 => n5352, B2 => n4387
                           , ZN => n5350);
   U322 : AOI221_X1 port map( B1 => n6991, B2 => n5353, C1 => n6959, C2 => 
                           n5354, A => n5355, ZN => n5340);
   U323 : OAI22_X1 port map( A1 => n5356, A2 => n4581, B1 => n5357, B2 => n4323
                           , ZN => n5355);
   U324 : AOI221_X1 port map( B1 => n5358, B2 => n5359, C1 => n5189, C2 => 
                           OUT1_31_port, A => n5360, ZN => n5339);
   U325 : OAI22_X1 port map( A1 => n5361, A2 => n4613, B1 => n5362, B2 => n4355
                           , ZN => n5360);
   U326 : NAND4_X1 port map( A1 => n5363, A2 => n5364, A3 => n5365, A4 => n5366
                           , ZN => n5359);
   U327 : AOI221_X1 port map( B1 => n6864, B2 => n5367, C1 => n6640, C2 => 
                           n5368, A => n5369, ZN => n5366);
   U328 : OAI222_X1 port map( A1 => n5370, A2 => n4709, B1 => n5371, B2 => 
                           n4163, C1 => n5372, C2 => n4419, ZN => n5369);
   U329 : AOI221_X1 port map( B1 => n6768, B2 => n5373, C1 => n6672, C2 => 
                           n5374, A => n5375, ZN => n5365);
   U330 : OAI22_X1 port map( A1 => n5376, A2 => n4485, B1 => n5377, B2 => n4227
                           , ZN => n5375);
   U331 : AOI221_X1 port map( B1 => n6704, B2 => n5378, C1 => n6800, C2 => 
                           n5379, A => n5380, ZN => n5364);
   U332 : OAI222_X1 port map( A1 => n5381, A2 => n4677, B1 => n5382, B2 => 
                           n4195, C1 => n5383, C2 => n4451, ZN => n5380);
   U333 : AOI221_X1 port map( B1 => n6736, B2 => n5384, C1 => n6832, C2 => 
                           n5385, A => n5386, ZN => n5363);
   U334 : OAI22_X1 port map( A1 => n5387, A2 => n4549, B1 => n5388, B2 => n4291
                           , ZN => n5386);
   U335 : NAND4_X1 port map( A1 => n5389, A2 => n5390, A3 => n5391, A4 => n5392
                           , ZN => n4161);
   U336 : AOI221_X1 port map( B1 => n7022, B2 => n5343, C1 => n7086, C2 => 
                           n5344, A => n5393, ZN => n5392);
   U337 : OAI22_X1 port map( A1 => n5346, A2 => n4518, B1 => n5347, B2 => n4260
                           , ZN => n5393);
   U338 : AOI221_X1 port map( B1 => n6897, B2 => n5348, C1 => n7054, C2 => 
                           n5349, A => n5394, ZN => n5391);
   U339 : OAI22_X1 port map( A1 => n5351, A2 => n4646, B1 => n5352, B2 => n4388
                           , ZN => n5394);
   U340 : AOI221_X1 port map( B1 => n6990, B2 => n5353, C1 => n6958, C2 => 
                           n5354, A => n5395, ZN => n5390);
   U341 : OAI22_X1 port map( A1 => n5356, A2 => n4582, B1 => n5357, B2 => n4324
                           , ZN => n5395);
   U342 : AOI221_X1 port map( B1 => n5358, B2 => n5396, C1 => n5189, C2 => 
                           OUT1_30_port, A => n5397, ZN => n5389);
   U343 : OAI22_X1 port map( A1 => n5361, A2 => n4614, B1 => n5362, B2 => n4356
                           , ZN => n5397);
   U344 : NAND4_X1 port map( A1 => n5398, A2 => n5399, A3 => n5400, A4 => n5401
                           , ZN => n5396);
   U345 : AOI221_X1 port map( B1 => n6865, B2 => n5367, C1 => n6641, C2 => 
                           n5368, A => n5402, ZN => n5401);
   U346 : OAI222_X1 port map( A1 => n5370, A2 => n4710, B1 => n5371, B2 => 
                           n4164, C1 => n5372, C2 => n4420, ZN => n5402);
   U347 : AOI221_X1 port map( B1 => n6769, B2 => n5373, C1 => n6673, C2 => 
                           n5374, A => n5403, ZN => n5400);
   U348 : OAI22_X1 port map( A1 => n5376, A2 => n4486, B1 => n5377, B2 => n4228
                           , ZN => n5403);
   U349 : AOI221_X1 port map( B1 => n6705, B2 => n5378, C1 => n6801, C2 => 
                           n5379, A => n5404, ZN => n5399);
   U350 : OAI222_X1 port map( A1 => n5381, A2 => n4678, B1 => n5382, B2 => 
                           n4196, C1 => n5383, C2 => n4452, ZN => n5404);
   U351 : AOI221_X1 port map( B1 => n6737, B2 => n5384, C1 => n6833, C2 => 
                           n5385, A => n5405, ZN => n5398);
   U352 : OAI22_X1 port map( A1 => n5387, A2 => n4550, B1 => n5388, B2 => n4292
                           , ZN => n5405);
   U353 : NAND4_X1 port map( A1 => n5406, A2 => n5407, A3 => n5408, A4 => n5409
                           , ZN => n4160);
   U354 : AOI221_X1 port map( B1 => n7021, B2 => n5343, C1 => n7085, C2 => 
                           n5344, A => n5410, ZN => n5409);
   U355 : OAI22_X1 port map( A1 => n5346, A2 => n4519, B1 => n5347, B2 => n4261
                           , ZN => n5410);
   U356 : AOI221_X1 port map( B1 => n6898, B2 => n5348, C1 => n7053, C2 => 
                           n5349, A => n5411, ZN => n5408);
   U357 : OAI22_X1 port map( A1 => n5351, A2 => n4647, B1 => n5352, B2 => n4389
                           , ZN => n5411);
   U358 : AOI221_X1 port map( B1 => n6989, B2 => n5353, C1 => n6957, C2 => 
                           n5354, A => n5412, ZN => n5407);
   U359 : OAI22_X1 port map( A1 => n5356, A2 => n4583, B1 => n5357, B2 => n4325
                           , ZN => n5412);
   U360 : AOI221_X1 port map( B1 => n5358, B2 => n5413, C1 => n5189, C2 => 
                           OUT1_29_port, A => n5414, ZN => n5406);
   U361 : OAI22_X1 port map( A1 => n5361, A2 => n4615, B1 => n5362, B2 => n4357
                           , ZN => n5414);
   U362 : NAND4_X1 port map( A1 => n5415, A2 => n5416, A3 => n5417, A4 => n5418
                           , ZN => n5413);
   U363 : AOI221_X1 port map( B1 => n6866, B2 => n5367, C1 => n6642, C2 => 
                           n5368, A => n5419, ZN => n5418);
   U364 : OAI222_X1 port map( A1 => n5370, A2 => n4711, B1 => n5371, B2 => 
                           n4165, C1 => n5372, C2 => n4421, ZN => n5419);
   U365 : AOI221_X1 port map( B1 => n6770, B2 => n5373, C1 => n6674, C2 => 
                           n5374, A => n5420, ZN => n5417);
   U366 : OAI22_X1 port map( A1 => n5376, A2 => n4487, B1 => n5377, B2 => n4229
                           , ZN => n5420);
   U367 : AOI221_X1 port map( B1 => n6706, B2 => n5378, C1 => n6802, C2 => 
                           n5379, A => n5421, ZN => n5416);
   U368 : OAI222_X1 port map( A1 => n5381, A2 => n4679, B1 => n5382, B2 => 
                           n4197, C1 => n5383, C2 => n4453, ZN => n5421);
   U369 : AOI221_X1 port map( B1 => n6738, B2 => n5384, C1 => n6834, C2 => 
                           n5385, A => n5422, ZN => n5415);
   U370 : OAI22_X1 port map( A1 => n5387, A2 => n4551, B1 => n5388, B2 => n4293
                           , ZN => n5422);
   U371 : NAND4_X1 port map( A1 => n5423, A2 => n5424, A3 => n5425, A4 => n5426
                           , ZN => n4159);
   U372 : AOI221_X1 port map( B1 => n7020, B2 => n5343, C1 => n7084, C2 => 
                           n5344, A => n5427, ZN => n5426);
   U373 : OAI22_X1 port map( A1 => n5346, A2 => n4520, B1 => n5347, B2 => n4262
                           , ZN => n5427);
   U374 : AOI221_X1 port map( B1 => n6899, B2 => n5348, C1 => n7052, C2 => 
                           n5349, A => n5428, ZN => n5425);
   U375 : OAI22_X1 port map( A1 => n5351, A2 => n4648, B1 => n5352, B2 => n4390
                           , ZN => n5428);
   U376 : AOI221_X1 port map( B1 => n6988, B2 => n5353, C1 => n6956, C2 => 
                           n5354, A => n5429, ZN => n5424);
   U377 : OAI22_X1 port map( A1 => n5356, A2 => n4584, B1 => n5357, B2 => n4326
                           , ZN => n5429);
   U378 : AOI221_X1 port map( B1 => n5358, B2 => n5430, C1 => n5189, C2 => 
                           OUT1_28_port, A => n5431, ZN => n5423);
   U379 : OAI22_X1 port map( A1 => n5361, A2 => n4616, B1 => n5362, B2 => n4358
                           , ZN => n5431);
   U380 : NAND4_X1 port map( A1 => n5432, A2 => n5433, A3 => n5434, A4 => n5435
                           , ZN => n5430);
   U381 : AOI221_X1 port map( B1 => n6867, B2 => n5367, C1 => n6643, C2 => 
                           n5368, A => n5436, ZN => n5435);
   U382 : OAI222_X1 port map( A1 => n5370, A2 => n4712, B1 => n5371, B2 => 
                           n4166, C1 => n5372, C2 => n4422, ZN => n5436);
   U383 : AOI221_X1 port map( B1 => n6771, B2 => n5373, C1 => n6675, C2 => 
                           n5374, A => n5437, ZN => n5434);
   U384 : OAI22_X1 port map( A1 => n5376, A2 => n4488, B1 => n5377, B2 => n4230
                           , ZN => n5437);
   U385 : AOI221_X1 port map( B1 => n6707, B2 => n5378, C1 => n6803, C2 => 
                           n5379, A => n5438, ZN => n5433);
   U386 : OAI222_X1 port map( A1 => n5381, A2 => n4680, B1 => n5382, B2 => 
                           n4198, C1 => n5383, C2 => n4454, ZN => n5438);
   U387 : AOI221_X1 port map( B1 => n6739, B2 => n5384, C1 => n6835, C2 => 
                           n5385, A => n5439, ZN => n5432);
   U388 : OAI22_X1 port map( A1 => n5387, A2 => n4552, B1 => n5388, B2 => n4294
                           , ZN => n5439);
   U389 : NAND4_X1 port map( A1 => n5440, A2 => n5441, A3 => n5442, A4 => n5443
                           , ZN => n4158);
   U390 : AOI221_X1 port map( B1 => n7019, B2 => n5343, C1 => n7083, C2 => 
                           n5344, A => n5444, ZN => n5443);
   U391 : OAI22_X1 port map( A1 => n5346, A2 => n4521, B1 => n5347, B2 => n4263
                           , ZN => n5444);
   U392 : AOI221_X1 port map( B1 => n6900, B2 => n5348, C1 => n7051, C2 => 
                           n5349, A => n5445, ZN => n5442);
   U393 : OAI22_X1 port map( A1 => n5351, A2 => n4649, B1 => n5352, B2 => n4391
                           , ZN => n5445);
   U394 : AOI221_X1 port map( B1 => n6987, B2 => n5353, C1 => n6955, C2 => 
                           n5354, A => n5446, ZN => n5441);
   U395 : OAI22_X1 port map( A1 => n5356, A2 => n4585, B1 => n5357, B2 => n4327
                           , ZN => n5446);
   U396 : AOI221_X1 port map( B1 => n5358, B2 => n5447, C1 => n5189, C2 => 
                           OUT1_27_port, A => n5448, ZN => n5440);
   U397 : OAI22_X1 port map( A1 => n5361, A2 => n4617, B1 => n5362, B2 => n4359
                           , ZN => n5448);
   U398 : NAND4_X1 port map( A1 => n5449, A2 => n5450, A3 => n5451, A4 => n5452
                           , ZN => n5447);
   U399 : AOI221_X1 port map( B1 => n6868, B2 => n5367, C1 => n6644, C2 => 
                           n5368, A => n5453, ZN => n5452);
   U400 : OAI222_X1 port map( A1 => n5370, A2 => n4713, B1 => n5371, B2 => 
                           n4167, C1 => n5372, C2 => n4423, ZN => n5453);
   U401 : AOI221_X1 port map( B1 => n6772, B2 => n5373, C1 => n6676, C2 => 
                           n5374, A => n5454, ZN => n5451);
   U402 : OAI22_X1 port map( A1 => n5376, A2 => n4489, B1 => n5377, B2 => n4231
                           , ZN => n5454);
   U403 : AOI221_X1 port map( B1 => n6708, B2 => n5378, C1 => n6804, C2 => 
                           n5379, A => n5455, ZN => n5450);
   U404 : OAI222_X1 port map( A1 => n5381, A2 => n4681, B1 => n5382, B2 => 
                           n4199, C1 => n5383, C2 => n4455, ZN => n5455);
   U405 : AOI221_X1 port map( B1 => n6740, B2 => n5384, C1 => n6836, C2 => 
                           n5385, A => n5456, ZN => n5449);
   U406 : OAI22_X1 port map( A1 => n5387, A2 => n4553, B1 => n5388, B2 => n4295
                           , ZN => n5456);
   U407 : NAND4_X1 port map( A1 => n5457, A2 => n5458, A3 => n5459, A4 => n5460
                           , ZN => n4157);
   U408 : AOI221_X1 port map( B1 => n7018, B2 => n5343, C1 => n7082, C2 => 
                           n5344, A => n5461, ZN => n5460);
   U409 : OAI22_X1 port map( A1 => n5346, A2 => n4522, B1 => n5347, B2 => n4264
                           , ZN => n5461);
   U410 : AOI221_X1 port map( B1 => n6901, B2 => n5348, C1 => n7050, C2 => 
                           n5349, A => n5462, ZN => n5459);
   U411 : OAI22_X1 port map( A1 => n5351, A2 => n4650, B1 => n5352, B2 => n4392
                           , ZN => n5462);
   U412 : AOI221_X1 port map( B1 => n6986, B2 => n5353, C1 => n6954, C2 => 
                           n5354, A => n5463, ZN => n5458);
   U413 : OAI22_X1 port map( A1 => n5356, A2 => n4586, B1 => n5357, B2 => n4328
                           , ZN => n5463);
   U414 : AOI221_X1 port map( B1 => n5358, B2 => n5464, C1 => n5189, C2 => 
                           OUT1_26_port, A => n5465, ZN => n5457);
   U415 : OAI22_X1 port map( A1 => n5361, A2 => n4618, B1 => n5362, B2 => n4360
                           , ZN => n5465);
   U416 : NAND4_X1 port map( A1 => n5466, A2 => n5467, A3 => n5468, A4 => n5469
                           , ZN => n5464);
   U417 : AOI221_X1 port map( B1 => n6869, B2 => n5367, C1 => n6645, C2 => 
                           n5368, A => n5470, ZN => n5469);
   U418 : OAI222_X1 port map( A1 => n5370, A2 => n4714, B1 => n5371, B2 => 
                           n4168, C1 => n5372, C2 => n4424, ZN => n5470);
   U419 : AOI221_X1 port map( B1 => n6773, B2 => n5373, C1 => n6677, C2 => 
                           n5374, A => n5471, ZN => n5468);
   U420 : OAI22_X1 port map( A1 => n5376, A2 => n4490, B1 => n5377, B2 => n4232
                           , ZN => n5471);
   U421 : AOI221_X1 port map( B1 => n6709, B2 => n5378, C1 => n6805, C2 => 
                           n5379, A => n5472, ZN => n5467);
   U422 : OAI222_X1 port map( A1 => n5381, A2 => n4682, B1 => n5382, B2 => 
                           n4200, C1 => n5383, C2 => n4456, ZN => n5472);
   U423 : AOI221_X1 port map( B1 => n6741, B2 => n5384, C1 => n6837, C2 => 
                           n5385, A => n5473, ZN => n5466);
   U424 : OAI22_X1 port map( A1 => n5387, A2 => n4554, B1 => n5388, B2 => n4296
                           , ZN => n5473);
   U425 : NAND4_X1 port map( A1 => n5474, A2 => n5475, A3 => n5476, A4 => n5477
                           , ZN => n4156);
   U426 : AOI221_X1 port map( B1 => n7017, B2 => n5343, C1 => n7081, C2 => 
                           n5344, A => n5478, ZN => n5477);
   U427 : OAI22_X1 port map( A1 => n5346, A2 => n4523, B1 => n5347, B2 => n4265
                           , ZN => n5478);
   U428 : AOI221_X1 port map( B1 => n6902, B2 => n5348, C1 => n7049, C2 => 
                           n5349, A => n5479, ZN => n5476);
   U429 : OAI22_X1 port map( A1 => n5351, A2 => n4651, B1 => n5352, B2 => n4393
                           , ZN => n5479);
   U430 : AOI221_X1 port map( B1 => n6985, B2 => n5353, C1 => n6953, C2 => 
                           n5354, A => n5480, ZN => n5475);
   U431 : OAI22_X1 port map( A1 => n5356, A2 => n4587, B1 => n5357, B2 => n4329
                           , ZN => n5480);
   U432 : AOI221_X1 port map( B1 => n5358, B2 => n5481, C1 => n5189, C2 => 
                           OUT1_25_port, A => n5482, ZN => n5474);
   U433 : OAI22_X1 port map( A1 => n5361, A2 => n4619, B1 => n5362, B2 => n4361
                           , ZN => n5482);
   U434 : NAND4_X1 port map( A1 => n5483, A2 => n5484, A3 => n5485, A4 => n5486
                           , ZN => n5481);
   U435 : AOI221_X1 port map( B1 => n6870, B2 => n5367, C1 => n6646, C2 => 
                           n5368, A => n5487, ZN => n5486);
   U436 : OAI222_X1 port map( A1 => n5370, A2 => n4715, B1 => n5371, B2 => 
                           n4169, C1 => n5372, C2 => n4425, ZN => n5487);
   U437 : AOI221_X1 port map( B1 => n6774, B2 => n5373, C1 => n6678, C2 => 
                           n5374, A => n5488, ZN => n5485);
   U438 : OAI22_X1 port map( A1 => n5376, A2 => n4491, B1 => n5377, B2 => n4233
                           , ZN => n5488);
   U439 : AOI221_X1 port map( B1 => n6710, B2 => n5378, C1 => n6806, C2 => 
                           n5379, A => n5489, ZN => n5484);
   U440 : OAI222_X1 port map( A1 => n5381, A2 => n4683, B1 => n5382, B2 => 
                           n4201, C1 => n5383, C2 => n4457, ZN => n5489);
   U441 : AOI221_X1 port map( B1 => n6742, B2 => n5384, C1 => n6838, C2 => 
                           n5385, A => n5490, ZN => n5483);
   U442 : OAI22_X1 port map( A1 => n5387, A2 => n4555, B1 => n5388, B2 => n4297
                           , ZN => n5490);
   U443 : NAND4_X1 port map( A1 => n5491, A2 => n5492, A3 => n5493, A4 => n5494
                           , ZN => n4155);
   U444 : AOI221_X1 port map( B1 => n7016, B2 => n5343, C1 => n7080, C2 => 
                           n5344, A => n5495, ZN => n5494);
   U445 : OAI22_X1 port map( A1 => n5346, A2 => n4524, B1 => n5347, B2 => n4266
                           , ZN => n5495);
   U446 : AOI221_X1 port map( B1 => n6903, B2 => n5348, C1 => n7048, C2 => 
                           n5349, A => n5496, ZN => n5493);
   U447 : OAI22_X1 port map( A1 => n5351, A2 => n4652, B1 => n5352, B2 => n4394
                           , ZN => n5496);
   U448 : AOI221_X1 port map( B1 => n6984, B2 => n5353, C1 => n6952, C2 => 
                           n5354, A => n5497, ZN => n5492);
   U449 : OAI22_X1 port map( A1 => n5356, A2 => n4588, B1 => n5357, B2 => n4330
                           , ZN => n5497);
   U450 : AOI221_X1 port map( B1 => n5358, B2 => n5498, C1 => n5189, C2 => 
                           OUT1_24_port, A => n5499, ZN => n5491);
   U451 : OAI22_X1 port map( A1 => n5361, A2 => n4620, B1 => n5362, B2 => n4362
                           , ZN => n5499);
   U452 : NAND4_X1 port map( A1 => n5500, A2 => n5501, A3 => n5502, A4 => n5503
                           , ZN => n5498);
   U453 : AOI221_X1 port map( B1 => n6871, B2 => n5367, C1 => n6647, C2 => 
                           n5368, A => n5504, ZN => n5503);
   U454 : OAI222_X1 port map( A1 => n5370, A2 => n4716, B1 => n5371, B2 => 
                           n4170, C1 => n5372, C2 => n4426, ZN => n5504);
   U455 : AOI221_X1 port map( B1 => n6775, B2 => n5373, C1 => n6679, C2 => 
                           n5374, A => n5505, ZN => n5502);
   U456 : OAI22_X1 port map( A1 => n5376, A2 => n4492, B1 => n5377, B2 => n4234
                           , ZN => n5505);
   U457 : AOI221_X1 port map( B1 => n6711, B2 => n5378, C1 => n6807, C2 => 
                           n5379, A => n5506, ZN => n5501);
   U458 : OAI222_X1 port map( A1 => n5381, A2 => n4684, B1 => n5382, B2 => 
                           n4202, C1 => n5383, C2 => n4458, ZN => n5506);
   U459 : AOI221_X1 port map( B1 => n6743, B2 => n5384, C1 => n6839, C2 => 
                           n5385, A => n5507, ZN => n5500);
   U460 : OAI22_X1 port map( A1 => n5387, A2 => n4556, B1 => n5388, B2 => n4298
                           , ZN => n5507);
   U461 : NAND4_X1 port map( A1 => n5508, A2 => n5509, A3 => n5510, A4 => n5511
                           , ZN => n4154);
   U462 : AOI221_X1 port map( B1 => n7015, B2 => n5343, C1 => n7079, C2 => 
                           n5344, A => n5512, ZN => n5511);
   U463 : OAI22_X1 port map( A1 => n5346, A2 => n4525, B1 => n5347, B2 => n4267
                           , ZN => n5512);
   U464 : AOI221_X1 port map( B1 => n6904, B2 => n5348, C1 => n7047, C2 => 
                           n5349, A => n5513, ZN => n5510);
   U465 : OAI22_X1 port map( A1 => n5351, A2 => n4653, B1 => n5352, B2 => n4395
                           , ZN => n5513);
   U466 : AOI221_X1 port map( B1 => n6983, B2 => n5353, C1 => n6951, C2 => 
                           n5354, A => n5514, ZN => n5509);
   U467 : OAI22_X1 port map( A1 => n5356, A2 => n4589, B1 => n5357, B2 => n4331
                           , ZN => n5514);
   U468 : AOI221_X1 port map( B1 => n5358, B2 => n5515, C1 => n5189, C2 => 
                           OUT1_23_port, A => n5516, ZN => n5508);
   U469 : OAI22_X1 port map( A1 => n5361, A2 => n4621, B1 => n5362, B2 => n4363
                           , ZN => n5516);
   U470 : NAND4_X1 port map( A1 => n5517, A2 => n5518, A3 => n5519, A4 => n5520
                           , ZN => n5515);
   U471 : AOI221_X1 port map( B1 => n6872, B2 => n5367, C1 => n6648, C2 => 
                           n5368, A => n5521, ZN => n5520);
   U472 : OAI222_X1 port map( A1 => n5370, A2 => n4717, B1 => n5371, B2 => 
                           n4171, C1 => n5372, C2 => n4427, ZN => n5521);
   U473 : AOI221_X1 port map( B1 => n6776, B2 => n5373, C1 => n6680, C2 => 
                           n5374, A => n5522, ZN => n5519);
   U474 : OAI22_X1 port map( A1 => n5376, A2 => n4493, B1 => n5377, B2 => n4235
                           , ZN => n5522);
   U475 : AOI221_X1 port map( B1 => n6712, B2 => n5378, C1 => n6808, C2 => 
                           n5379, A => n5523, ZN => n5518);
   U476 : OAI222_X1 port map( A1 => n5381, A2 => n4685, B1 => n5382, B2 => 
                           n4203, C1 => n5383, C2 => n4459, ZN => n5523);
   U477 : AOI221_X1 port map( B1 => n6744, B2 => n5384, C1 => n6840, C2 => 
                           n5385, A => n5524, ZN => n5517);
   U478 : OAI22_X1 port map( A1 => n5387, A2 => n4557, B1 => n5388, B2 => n4299
                           , ZN => n5524);
   U479 : NAND4_X1 port map( A1 => n5525, A2 => n5526, A3 => n5527, A4 => n5528
                           , ZN => n4153);
   U480 : AOI221_X1 port map( B1 => n7014, B2 => n5343, C1 => n7078, C2 => 
                           n5344, A => n5529, ZN => n5528);
   U481 : OAI22_X1 port map( A1 => n5346, A2 => n4526, B1 => n5347, B2 => n4268
                           , ZN => n5529);
   U482 : AOI221_X1 port map( B1 => n6905, B2 => n5348, C1 => n7046, C2 => 
                           n5349, A => n5530, ZN => n5527);
   U483 : OAI22_X1 port map( A1 => n5351, A2 => n4654, B1 => n5352, B2 => n4396
                           , ZN => n5530);
   U484 : AOI221_X1 port map( B1 => n6982, B2 => n5353, C1 => n6950, C2 => 
                           n5354, A => n5531, ZN => n5526);
   U485 : OAI22_X1 port map( A1 => n5356, A2 => n4590, B1 => n5357, B2 => n4332
                           , ZN => n5531);
   U486 : AOI221_X1 port map( B1 => n5358, B2 => n5532, C1 => n5189, C2 => 
                           OUT1_22_port, A => n5533, ZN => n5525);
   U487 : OAI22_X1 port map( A1 => n5361, A2 => n4622, B1 => n5362, B2 => n4364
                           , ZN => n5533);
   U488 : NAND4_X1 port map( A1 => n5534, A2 => n5535, A3 => n5536, A4 => n5537
                           , ZN => n5532);
   U489 : AOI221_X1 port map( B1 => n6873, B2 => n5367, C1 => n6649, C2 => 
                           n5368, A => n5538, ZN => n5537);
   U490 : OAI222_X1 port map( A1 => n5370, A2 => n4718, B1 => n5371, B2 => 
                           n4172, C1 => n5372, C2 => n4428, ZN => n5538);
   U491 : AOI221_X1 port map( B1 => n6777, B2 => n5373, C1 => n6681, C2 => 
                           n5374, A => n5539, ZN => n5536);
   U492 : OAI22_X1 port map( A1 => n5376, A2 => n4494, B1 => n5377, B2 => n4236
                           , ZN => n5539);
   U493 : AOI221_X1 port map( B1 => n6713, B2 => n5378, C1 => n6809, C2 => 
                           n5379, A => n5540, ZN => n5535);
   U494 : OAI222_X1 port map( A1 => n5381, A2 => n4686, B1 => n5382, B2 => 
                           n4204, C1 => n5383, C2 => n4460, ZN => n5540);
   U495 : AOI221_X1 port map( B1 => n6745, B2 => n5384, C1 => n6841, C2 => 
                           n5385, A => n5541, ZN => n5534);
   U496 : OAI22_X1 port map( A1 => n5387, A2 => n4558, B1 => n5388, B2 => n4300
                           , ZN => n5541);
   U497 : NAND4_X1 port map( A1 => n5542, A2 => n5543, A3 => n5544, A4 => n5545
                           , ZN => n4152);
   U498 : AOI221_X1 port map( B1 => n7013, B2 => n5343, C1 => n7077, C2 => 
                           n5344, A => n5546, ZN => n5545);
   U499 : OAI22_X1 port map( A1 => n5346, A2 => n4527, B1 => n5347, B2 => n4269
                           , ZN => n5546);
   U500 : AOI221_X1 port map( B1 => n6906, B2 => n5348, C1 => n7045, C2 => 
                           n5349, A => n5547, ZN => n5544);
   U501 : OAI22_X1 port map( A1 => n5351, A2 => n4655, B1 => n5352, B2 => n4397
                           , ZN => n5547);
   U502 : AOI221_X1 port map( B1 => n6981, B2 => n5353, C1 => n6949, C2 => 
                           n5354, A => n5548, ZN => n5543);
   U503 : OAI22_X1 port map( A1 => n5356, A2 => n4591, B1 => n5357, B2 => n4333
                           , ZN => n5548);
   U504 : AOI221_X1 port map( B1 => n5358, B2 => n5549, C1 => n5189, C2 => 
                           OUT1_21_port, A => n5550, ZN => n5542);
   U505 : OAI22_X1 port map( A1 => n5361, A2 => n4623, B1 => n5362, B2 => n4365
                           , ZN => n5550);
   U506 : NAND4_X1 port map( A1 => n5551, A2 => n5552, A3 => n5553, A4 => n5554
                           , ZN => n5549);
   U507 : AOI221_X1 port map( B1 => n6874, B2 => n5367, C1 => n6650, C2 => 
                           n5368, A => n5555, ZN => n5554);
   U508 : OAI222_X1 port map( A1 => n5370, A2 => n4719, B1 => n5371, B2 => 
                           n4173, C1 => n5372, C2 => n4429, ZN => n5555);
   U509 : AOI221_X1 port map( B1 => n6778, B2 => n5373, C1 => n6682, C2 => 
                           n5374, A => n5556, ZN => n5553);
   U510 : OAI22_X1 port map( A1 => n5376, A2 => n4495, B1 => n5377, B2 => n4237
                           , ZN => n5556);
   U511 : AOI221_X1 port map( B1 => n6714, B2 => n5378, C1 => n6810, C2 => 
                           n5379, A => n5557, ZN => n5552);
   U512 : OAI222_X1 port map( A1 => n5381, A2 => n4687, B1 => n5382, B2 => 
                           n4205, C1 => n5383, C2 => n4461, ZN => n5557);
   U513 : AOI221_X1 port map( B1 => n6746, B2 => n5384, C1 => n6842, C2 => 
                           n5385, A => n5558, ZN => n5551);
   U514 : OAI22_X1 port map( A1 => n5387, A2 => n4559, B1 => n5388, B2 => n4301
                           , ZN => n5558);
   U515 : NAND4_X1 port map( A1 => n5559, A2 => n5560, A3 => n5561, A4 => n5562
                           , ZN => n4151);
   U516 : AOI221_X1 port map( B1 => n7012, B2 => n5343, C1 => n7076, C2 => 
                           n5344, A => n5563, ZN => n5562);
   U517 : OAI22_X1 port map( A1 => n5346, A2 => n4528, B1 => n5347, B2 => n4270
                           , ZN => n5563);
   U518 : AOI221_X1 port map( B1 => n6907, B2 => n5348, C1 => n7044, C2 => 
                           n5349, A => n5564, ZN => n5561);
   U519 : OAI22_X1 port map( A1 => n5351, A2 => n4656, B1 => n5352, B2 => n4398
                           , ZN => n5564);
   U520 : AOI221_X1 port map( B1 => n6980, B2 => n5353, C1 => n6948, C2 => 
                           n5354, A => n5565, ZN => n5560);
   U521 : OAI22_X1 port map( A1 => n5356, A2 => n4592, B1 => n5357, B2 => n4334
                           , ZN => n5565);
   U522 : AOI221_X1 port map( B1 => n5358, B2 => n5566, C1 => n5189, C2 => 
                           OUT1_20_port, A => n5567, ZN => n5559);
   U523 : OAI22_X1 port map( A1 => n5361, A2 => n4624, B1 => n5362, B2 => n4366
                           , ZN => n5567);
   U524 : NAND4_X1 port map( A1 => n5568, A2 => n5569, A3 => n5570, A4 => n5571
                           , ZN => n5566);
   U525 : AOI221_X1 port map( B1 => n6875, B2 => n5367, C1 => n6651, C2 => 
                           n5368, A => n5572, ZN => n5571);
   U526 : OAI222_X1 port map( A1 => n5370, A2 => n4720, B1 => n5371, B2 => 
                           n4174, C1 => n5372, C2 => n4430, ZN => n5572);
   U527 : AOI221_X1 port map( B1 => n6779, B2 => n5373, C1 => n6683, C2 => 
                           n5374, A => n5573, ZN => n5570);
   U528 : OAI22_X1 port map( A1 => n5376, A2 => n4496, B1 => n5377, B2 => n4238
                           , ZN => n5573);
   U529 : AOI221_X1 port map( B1 => n6715, B2 => n5378, C1 => n6811, C2 => 
                           n5379, A => n5574, ZN => n5569);
   U530 : OAI222_X1 port map( A1 => n5381, A2 => n4688, B1 => n5382, B2 => 
                           n4206, C1 => n5383, C2 => n4462, ZN => n5574);
   U531 : AOI221_X1 port map( B1 => n6747, B2 => n5384, C1 => n6843, C2 => 
                           n5385, A => n5575, ZN => n5568);
   U532 : OAI22_X1 port map( A1 => n5387, A2 => n4560, B1 => n5388, B2 => n4302
                           , ZN => n5575);
   U533 : NAND4_X1 port map( A1 => n5576, A2 => n5577, A3 => n5578, A4 => n5579
                           , ZN => n4150);
   U534 : AOI221_X1 port map( B1 => n7011, B2 => n5343, C1 => n7075, C2 => 
                           n5344, A => n5580, ZN => n5579);
   U535 : OAI22_X1 port map( A1 => n5346, A2 => n4529, B1 => n5347, B2 => n4271
                           , ZN => n5580);
   U536 : AOI221_X1 port map( B1 => n6908, B2 => n5348, C1 => n7043, C2 => 
                           n5349, A => n5581, ZN => n5578);
   U537 : OAI22_X1 port map( A1 => n5351, A2 => n4657, B1 => n5352, B2 => n4399
                           , ZN => n5581);
   U538 : AOI221_X1 port map( B1 => n6979, B2 => n5353, C1 => n6947, C2 => 
                           n5354, A => n5582, ZN => n5577);
   U539 : OAI22_X1 port map( A1 => n5356, A2 => n4593, B1 => n5357, B2 => n4335
                           , ZN => n5582);
   U540 : AOI221_X1 port map( B1 => n5358, B2 => n5583, C1 => n5189, C2 => 
                           OUT1_19_port, A => n5584, ZN => n5576);
   U541 : OAI22_X1 port map( A1 => n5361, A2 => n4625, B1 => n5362, B2 => n4367
                           , ZN => n5584);
   U542 : NAND4_X1 port map( A1 => n5585, A2 => n5586, A3 => n5587, A4 => n5588
                           , ZN => n5583);
   U543 : AOI221_X1 port map( B1 => n6876, B2 => n5367, C1 => n6652, C2 => 
                           n5368, A => n5589, ZN => n5588);
   U544 : OAI222_X1 port map( A1 => n5370, A2 => n4721, B1 => n5371, B2 => 
                           n4175, C1 => n5372, C2 => n4431, ZN => n5589);
   U545 : AOI221_X1 port map( B1 => n6780, B2 => n5373, C1 => n6684, C2 => 
                           n5374, A => n5590, ZN => n5587);
   U546 : OAI22_X1 port map( A1 => n5376, A2 => n4497, B1 => n5377, B2 => n4239
                           , ZN => n5590);
   U547 : AOI221_X1 port map( B1 => n6716, B2 => n5378, C1 => n6812, C2 => 
                           n5379, A => n5591, ZN => n5586);
   U548 : OAI222_X1 port map( A1 => n5381, A2 => n4689, B1 => n5382, B2 => 
                           n4207, C1 => n5383, C2 => n4463, ZN => n5591);
   U549 : AOI221_X1 port map( B1 => n6748, B2 => n5384, C1 => n6844, C2 => 
                           n5385, A => n5592, ZN => n5585);
   U550 : OAI22_X1 port map( A1 => n5387, A2 => n4561, B1 => n5388, B2 => n4303
                           , ZN => n5592);
   U551 : NAND4_X1 port map( A1 => n5593, A2 => n5594, A3 => n5595, A4 => n5596
                           , ZN => n4149);
   U552 : AOI221_X1 port map( B1 => n7010, B2 => n5343, C1 => n7074, C2 => 
                           n5344, A => n5597, ZN => n5596);
   U553 : OAI22_X1 port map( A1 => n5346, A2 => n4530, B1 => n5347, B2 => n4272
                           , ZN => n5597);
   U554 : AOI221_X1 port map( B1 => n6909, B2 => n5348, C1 => n7042, C2 => 
                           n5349, A => n5598, ZN => n5595);
   U555 : OAI22_X1 port map( A1 => n5351, A2 => n4658, B1 => n5352, B2 => n4400
                           , ZN => n5598);
   U556 : AOI221_X1 port map( B1 => n6978, B2 => n5353, C1 => n6946, C2 => 
                           n5354, A => n5599, ZN => n5594);
   U557 : OAI22_X1 port map( A1 => n5356, A2 => n4594, B1 => n5357, B2 => n4336
                           , ZN => n5599);
   U558 : AOI221_X1 port map( B1 => n5358, B2 => n5600, C1 => n5189, C2 => 
                           OUT1_18_port, A => n5601, ZN => n5593);
   U559 : OAI22_X1 port map( A1 => n5361, A2 => n4626, B1 => n5362, B2 => n4368
                           , ZN => n5601);
   U560 : NAND4_X1 port map( A1 => n5602, A2 => n5603, A3 => n5604, A4 => n5605
                           , ZN => n5600);
   U561 : AOI221_X1 port map( B1 => n6877, B2 => n5367, C1 => n6653, C2 => 
                           n5368, A => n5606, ZN => n5605);
   U562 : OAI222_X1 port map( A1 => n5370, A2 => n4722, B1 => n5371, B2 => 
                           n4176, C1 => n5372, C2 => n4432, ZN => n5606);
   U563 : AOI221_X1 port map( B1 => n6781, B2 => n5373, C1 => n6685, C2 => 
                           n5374, A => n5607, ZN => n5604);
   U564 : OAI22_X1 port map( A1 => n5376, A2 => n4498, B1 => n5377, B2 => n4240
                           , ZN => n5607);
   U565 : AOI221_X1 port map( B1 => n6717, B2 => n5378, C1 => n6813, C2 => 
                           n5379, A => n5608, ZN => n5603);
   U566 : OAI222_X1 port map( A1 => n5381, A2 => n4690, B1 => n5382, B2 => 
                           n4208, C1 => n5383, C2 => n4464, ZN => n5608);
   U567 : AOI221_X1 port map( B1 => n6749, B2 => n5384, C1 => n6845, C2 => 
                           n5385, A => n5609, ZN => n5602);
   U568 : OAI22_X1 port map( A1 => n5387, A2 => n4562, B1 => n5388, B2 => n4304
                           , ZN => n5609);
   U569 : NAND4_X1 port map( A1 => n5610, A2 => n5611, A3 => n5612, A4 => n5613
                           , ZN => n4148);
   U570 : AOI221_X1 port map( B1 => n7009, B2 => n5343, C1 => n7073, C2 => 
                           n5344, A => n5614, ZN => n5613);
   U571 : OAI22_X1 port map( A1 => n5346, A2 => n4531, B1 => n5347, B2 => n4273
                           , ZN => n5614);
   U572 : AOI221_X1 port map( B1 => n6910, B2 => n5348, C1 => n7041, C2 => 
                           n5349, A => n5615, ZN => n5612);
   U573 : OAI22_X1 port map( A1 => n5351, A2 => n4659, B1 => n5352, B2 => n4401
                           , ZN => n5615);
   U574 : AOI221_X1 port map( B1 => n6977, B2 => n5353, C1 => n6945, C2 => 
                           n5354, A => n5616, ZN => n5611);
   U575 : OAI22_X1 port map( A1 => n5356, A2 => n4595, B1 => n5357, B2 => n4337
                           , ZN => n5616);
   U576 : AOI221_X1 port map( B1 => n5358, B2 => n5617, C1 => n5189, C2 => 
                           OUT1_17_port, A => n5618, ZN => n5610);
   U577 : OAI22_X1 port map( A1 => n5361, A2 => n4627, B1 => n5362, B2 => n4369
                           , ZN => n5618);
   U578 : NAND4_X1 port map( A1 => n5619, A2 => n5620, A3 => n5621, A4 => n5622
                           , ZN => n5617);
   U579 : AOI221_X1 port map( B1 => n6878, B2 => n5367, C1 => n6654, C2 => 
                           n5368, A => n5623, ZN => n5622);
   U580 : OAI222_X1 port map( A1 => n5370, A2 => n4723, B1 => n5371, B2 => 
                           n4177, C1 => n5372, C2 => n4433, ZN => n5623);
   U581 : AOI221_X1 port map( B1 => n6782, B2 => n5373, C1 => n6686, C2 => 
                           n5374, A => n5624, ZN => n5621);
   U582 : OAI22_X1 port map( A1 => n5376, A2 => n4499, B1 => n5377, B2 => n4241
                           , ZN => n5624);
   U583 : AOI221_X1 port map( B1 => n6718, B2 => n5378, C1 => n6814, C2 => 
                           n5379, A => n5625, ZN => n5620);
   U584 : OAI222_X1 port map( A1 => n5381, A2 => n4691, B1 => n5382, B2 => 
                           n4209, C1 => n5383, C2 => n4465, ZN => n5625);
   U585 : AOI221_X1 port map( B1 => n6750, B2 => n5384, C1 => n6846, C2 => 
                           n5385, A => n5626, ZN => n5619);
   U586 : OAI22_X1 port map( A1 => n5387, A2 => n4563, B1 => n5388, B2 => n4305
                           , ZN => n5626);
   U587 : NAND4_X1 port map( A1 => n5627, A2 => n5628, A3 => n5629, A4 => n5630
                           , ZN => n4147);
   U588 : AOI221_X1 port map( B1 => n7008, B2 => n5343, C1 => n7072, C2 => 
                           n5344, A => n5631, ZN => n5630);
   U589 : OAI22_X1 port map( A1 => n5346, A2 => n4532, B1 => n5347, B2 => n4274
                           , ZN => n5631);
   U590 : AOI221_X1 port map( B1 => n6911, B2 => n5348, C1 => n7040, C2 => 
                           n5349, A => n5632, ZN => n5629);
   U591 : OAI22_X1 port map( A1 => n5351, A2 => n4660, B1 => n5352, B2 => n4402
                           , ZN => n5632);
   U592 : AOI221_X1 port map( B1 => n6976, B2 => n5353, C1 => n6944, C2 => 
                           n5354, A => n5633, ZN => n5628);
   U593 : OAI22_X1 port map( A1 => n5356, A2 => n4596, B1 => n5357, B2 => n4338
                           , ZN => n5633);
   U594 : AOI221_X1 port map( B1 => n5358, B2 => n5634, C1 => n5189, C2 => 
                           OUT1_16_port, A => n5635, ZN => n5627);
   U595 : OAI22_X1 port map( A1 => n5361, A2 => n4628, B1 => n5362, B2 => n4370
                           , ZN => n5635);
   U596 : NAND4_X1 port map( A1 => n5636, A2 => n5637, A3 => n5638, A4 => n5639
                           , ZN => n5634);
   U597 : AOI221_X1 port map( B1 => n6879, B2 => n5367, C1 => n6655, C2 => 
                           n5368, A => n5640, ZN => n5639);
   U598 : OAI222_X1 port map( A1 => n5370, A2 => n4724, B1 => n5371, B2 => 
                           n4178, C1 => n5372, C2 => n4434, ZN => n5640);
   U599 : AOI221_X1 port map( B1 => n6783, B2 => n5373, C1 => n6687, C2 => 
                           n5374, A => n5641, ZN => n5638);
   U600 : OAI22_X1 port map( A1 => n5376, A2 => n4500, B1 => n5377, B2 => n4242
                           , ZN => n5641);
   U601 : AOI221_X1 port map( B1 => n6719, B2 => n5378, C1 => n6815, C2 => 
                           n5379, A => n5642, ZN => n5637);
   U602 : OAI222_X1 port map( A1 => n5381, A2 => n4692, B1 => n5382, B2 => 
                           n4210, C1 => n5383, C2 => n4466, ZN => n5642);
   U603 : AOI221_X1 port map( B1 => n6751, B2 => n5384, C1 => n6847, C2 => 
                           n5385, A => n5643, ZN => n5636);
   U604 : OAI22_X1 port map( A1 => n5387, A2 => n4564, B1 => n5388, B2 => n4306
                           , ZN => n5643);
   U605 : NAND4_X1 port map( A1 => n5644, A2 => n5645, A3 => n5646, A4 => n5647
                           , ZN => n4146);
   U606 : AOI221_X1 port map( B1 => n7007, B2 => n5343, C1 => n7071, C2 => 
                           n5344, A => n5648, ZN => n5647);
   U607 : OAI22_X1 port map( A1 => n5346, A2 => n4533, B1 => n5347, B2 => n4275
                           , ZN => n5648);
   U608 : AOI221_X1 port map( B1 => n6912, B2 => n5348, C1 => n7039, C2 => 
                           n5349, A => n5649, ZN => n5646);
   U609 : OAI22_X1 port map( A1 => n5351, A2 => n4661, B1 => n5352, B2 => n4403
                           , ZN => n5649);
   U610 : AOI221_X1 port map( B1 => n6975, B2 => n5353, C1 => n6943, C2 => 
                           n5354, A => n5650, ZN => n5645);
   U611 : OAI22_X1 port map( A1 => n5356, A2 => n4597, B1 => n5357, B2 => n4339
                           , ZN => n5650);
   U612 : AOI221_X1 port map( B1 => n5358, B2 => n5651, C1 => n5189, C2 => 
                           OUT1_15_port, A => n5652, ZN => n5644);
   U613 : OAI22_X1 port map( A1 => n5361, A2 => n4629, B1 => n5362, B2 => n4371
                           , ZN => n5652);
   U614 : NAND4_X1 port map( A1 => n5653, A2 => n5654, A3 => n5655, A4 => n5656
                           , ZN => n5651);
   U615 : AOI221_X1 port map( B1 => n6880, B2 => n5367, C1 => n6656, C2 => 
                           n5368, A => n5657, ZN => n5656);
   U616 : OAI222_X1 port map( A1 => n5370, A2 => n4725, B1 => n5371, B2 => 
                           n4179, C1 => n5372, C2 => n4435, ZN => n5657);
   U617 : AOI221_X1 port map( B1 => n6784, B2 => n5373, C1 => n6688, C2 => 
                           n5374, A => n5658, ZN => n5655);
   U618 : OAI22_X1 port map( A1 => n5376, A2 => n4501, B1 => n5377, B2 => n4243
                           , ZN => n5658);
   U619 : AOI221_X1 port map( B1 => n6720, B2 => n5378, C1 => n6816, C2 => 
                           n5379, A => n5659, ZN => n5654);
   U620 : OAI222_X1 port map( A1 => n5381, A2 => n4693, B1 => n5382, B2 => 
                           n4211, C1 => n5383, C2 => n4467, ZN => n5659);
   U621 : AOI221_X1 port map( B1 => n6752, B2 => n5384, C1 => n6848, C2 => 
                           n5385, A => n5660, ZN => n5653);
   U622 : OAI22_X1 port map( A1 => n5387, A2 => n4565, B1 => n5388, B2 => n4307
                           , ZN => n5660);
   U623 : NAND4_X1 port map( A1 => n5661, A2 => n5662, A3 => n5663, A4 => n5664
                           , ZN => n4145);
   U624 : AOI221_X1 port map( B1 => n7006, B2 => n5343, C1 => n7070, C2 => 
                           n5344, A => n5665, ZN => n5664);
   U625 : OAI22_X1 port map( A1 => n5346, A2 => n4534, B1 => n5347, B2 => n4276
                           , ZN => n5665);
   U626 : AOI221_X1 port map( B1 => n6913, B2 => n5348, C1 => n7038, C2 => 
                           n5349, A => n5666, ZN => n5663);
   U627 : OAI22_X1 port map( A1 => n5351, A2 => n4662, B1 => n5352, B2 => n4404
                           , ZN => n5666);
   U628 : AOI221_X1 port map( B1 => n6974, B2 => n5353, C1 => n6942, C2 => 
                           n5354, A => n5667, ZN => n5662);
   U629 : OAI22_X1 port map( A1 => n5356, A2 => n4598, B1 => n5357, B2 => n4340
                           , ZN => n5667);
   U630 : AOI221_X1 port map( B1 => n5358, B2 => n5668, C1 => n5189, C2 => 
                           OUT1_14_port, A => n5669, ZN => n5661);
   U631 : OAI22_X1 port map( A1 => n5361, A2 => n4630, B1 => n5362, B2 => n4372
                           , ZN => n5669);
   U632 : NAND4_X1 port map( A1 => n5670, A2 => n5671, A3 => n5672, A4 => n5673
                           , ZN => n5668);
   U633 : AOI221_X1 port map( B1 => n6881, B2 => n5367, C1 => n6657, C2 => 
                           n5368, A => n5674, ZN => n5673);
   U634 : OAI222_X1 port map( A1 => n5370, A2 => n4726, B1 => n5371, B2 => 
                           n4180, C1 => n5372, C2 => n4436, ZN => n5674);
   U635 : AOI221_X1 port map( B1 => n6785, B2 => n5373, C1 => n6689, C2 => 
                           n5374, A => n5675, ZN => n5672);
   U636 : OAI22_X1 port map( A1 => n5376, A2 => n4502, B1 => n5377, B2 => n4244
                           , ZN => n5675);
   U637 : AOI221_X1 port map( B1 => n6721, B2 => n5378, C1 => n6817, C2 => 
                           n5379, A => n5676, ZN => n5671);
   U638 : OAI222_X1 port map( A1 => n5381, A2 => n4694, B1 => n5382, B2 => 
                           n4212, C1 => n5383, C2 => n4468, ZN => n5676);
   U639 : AOI221_X1 port map( B1 => n6753, B2 => n5384, C1 => n6849, C2 => 
                           n5385, A => n5677, ZN => n5670);
   U640 : OAI22_X1 port map( A1 => n5387, A2 => n4566, B1 => n5388, B2 => n4308
                           , ZN => n5677);
   U641 : NAND4_X1 port map( A1 => n5678, A2 => n5679, A3 => n5680, A4 => n5681
                           , ZN => n4144);
   U642 : AOI221_X1 port map( B1 => n7005, B2 => n5343, C1 => n7069, C2 => 
                           n5344, A => n5682, ZN => n5681);
   U643 : OAI22_X1 port map( A1 => n5346, A2 => n4535, B1 => n5347, B2 => n4277
                           , ZN => n5682);
   U644 : AOI221_X1 port map( B1 => n6914, B2 => n5348, C1 => n7037, C2 => 
                           n5349, A => n5683, ZN => n5680);
   U645 : OAI22_X1 port map( A1 => n5351, A2 => n4663, B1 => n5352, B2 => n4405
                           , ZN => n5683);
   U646 : AOI221_X1 port map( B1 => n6973, B2 => n5353, C1 => n6941, C2 => 
                           n5354, A => n5684, ZN => n5679);
   U647 : OAI22_X1 port map( A1 => n5356, A2 => n4599, B1 => n5357, B2 => n4341
                           , ZN => n5684);
   U648 : AOI221_X1 port map( B1 => n5358, B2 => n5685, C1 => n5189, C2 => 
                           OUT1_13_port, A => n5686, ZN => n5678);
   U649 : OAI22_X1 port map( A1 => n5361, A2 => n4631, B1 => n5362, B2 => n4373
                           , ZN => n5686);
   U650 : NAND4_X1 port map( A1 => n5687, A2 => n5688, A3 => n5689, A4 => n5690
                           , ZN => n5685);
   U651 : AOI221_X1 port map( B1 => n6882, B2 => n5367, C1 => n6658, C2 => 
                           n5368, A => n5691, ZN => n5690);
   U652 : OAI222_X1 port map( A1 => n5370, A2 => n4727, B1 => n5371, B2 => 
                           n4181, C1 => n5372, C2 => n4437, ZN => n5691);
   U653 : AOI221_X1 port map( B1 => n6786, B2 => n5373, C1 => n6690, C2 => 
                           n5374, A => n5692, ZN => n5689);
   U654 : OAI22_X1 port map( A1 => n5376, A2 => n4503, B1 => n5377, B2 => n4245
                           , ZN => n5692);
   U655 : AOI221_X1 port map( B1 => n6722, B2 => n5378, C1 => n6818, C2 => 
                           n5379, A => n5693, ZN => n5688);
   U656 : OAI222_X1 port map( A1 => n5381, A2 => n4695, B1 => n5382, B2 => 
                           n4213, C1 => n5383, C2 => n4469, ZN => n5693);
   U657 : AOI221_X1 port map( B1 => n6754, B2 => n5384, C1 => n6850, C2 => 
                           n5385, A => n5694, ZN => n5687);
   U658 : OAI22_X1 port map( A1 => n5387, A2 => n4567, B1 => n5388, B2 => n4309
                           , ZN => n5694);
   U659 : NAND4_X1 port map( A1 => n5695, A2 => n5696, A3 => n5697, A4 => n5698
                           , ZN => n4143);
   U660 : AOI221_X1 port map( B1 => n7004, B2 => n5343, C1 => n7068, C2 => 
                           n5344, A => n5699, ZN => n5698);
   U661 : OAI22_X1 port map( A1 => n5346, A2 => n4536, B1 => n5347, B2 => n4278
                           , ZN => n5699);
   U662 : AOI221_X1 port map( B1 => n6915, B2 => n5348, C1 => n7036, C2 => 
                           n5349, A => n5700, ZN => n5697);
   U663 : OAI22_X1 port map( A1 => n5351, A2 => n4664, B1 => n5352, B2 => n4406
                           , ZN => n5700);
   U664 : AOI221_X1 port map( B1 => n6972, B2 => n5353, C1 => n6940, C2 => 
                           n5354, A => n5701, ZN => n5696);
   U665 : OAI22_X1 port map( A1 => n5356, A2 => n4600, B1 => n5357, B2 => n4342
                           , ZN => n5701);
   U666 : AOI221_X1 port map( B1 => n5358, B2 => n5702, C1 => n5189, C2 => 
                           OUT1_12_port, A => n5703, ZN => n5695);
   U667 : OAI22_X1 port map( A1 => n5361, A2 => n4632, B1 => n5362, B2 => n4374
                           , ZN => n5703);
   U668 : NAND4_X1 port map( A1 => n5704, A2 => n5705, A3 => n5706, A4 => n5707
                           , ZN => n5702);
   U669 : AOI221_X1 port map( B1 => n6883, B2 => n5367, C1 => n6659, C2 => 
                           n5368, A => n5708, ZN => n5707);
   U670 : OAI222_X1 port map( A1 => n5370, A2 => n4728, B1 => n5371, B2 => 
                           n4182, C1 => n5372, C2 => n4438, ZN => n5708);
   U671 : AOI221_X1 port map( B1 => n6787, B2 => n5373, C1 => n6691, C2 => 
                           n5374, A => n5709, ZN => n5706);
   U672 : OAI22_X1 port map( A1 => n5376, A2 => n4504, B1 => n5377, B2 => n4246
                           , ZN => n5709);
   U673 : AOI221_X1 port map( B1 => n6723, B2 => n5378, C1 => n6819, C2 => 
                           n5379, A => n5710, ZN => n5705);
   U674 : OAI222_X1 port map( A1 => n5381, A2 => n4696, B1 => n5382, B2 => 
                           n4214, C1 => n5383, C2 => n4470, ZN => n5710);
   U675 : AOI221_X1 port map( B1 => n6755, B2 => n5384, C1 => n6851, C2 => 
                           n5385, A => n5711, ZN => n5704);
   U676 : OAI22_X1 port map( A1 => n5387, A2 => n4568, B1 => n5388, B2 => n4310
                           , ZN => n5711);
   U677 : NAND4_X1 port map( A1 => n5712, A2 => n5713, A3 => n5714, A4 => n5715
                           , ZN => n4142);
   U678 : AOI221_X1 port map( B1 => n7003, B2 => n5343, C1 => n7067, C2 => 
                           n5344, A => n5716, ZN => n5715);
   U679 : OAI22_X1 port map( A1 => n5346, A2 => n4537, B1 => n5347, B2 => n4279
                           , ZN => n5716);
   U680 : AOI221_X1 port map( B1 => n6916, B2 => n5348, C1 => n7035, C2 => 
                           n5349, A => n5717, ZN => n5714);
   U681 : OAI22_X1 port map( A1 => n5351, A2 => n4665, B1 => n5352, B2 => n4407
                           , ZN => n5717);
   U682 : AOI221_X1 port map( B1 => n6971, B2 => n5353, C1 => n6939, C2 => 
                           n5354, A => n5718, ZN => n5713);
   U683 : OAI22_X1 port map( A1 => n5356, A2 => n4601, B1 => n5357, B2 => n4343
                           , ZN => n5718);
   U684 : AOI221_X1 port map( B1 => n5358, B2 => n5719, C1 => n5189, C2 => 
                           OUT1_11_port, A => n5720, ZN => n5712);
   U685 : OAI22_X1 port map( A1 => n5361, A2 => n4633, B1 => n5362, B2 => n4375
                           , ZN => n5720);
   U686 : NAND4_X1 port map( A1 => n5721, A2 => n5722, A3 => n5723, A4 => n5724
                           , ZN => n5719);
   U687 : AOI221_X1 port map( B1 => n6884, B2 => n5367, C1 => n6660, C2 => 
                           n5368, A => n5725, ZN => n5724);
   U688 : OAI222_X1 port map( A1 => n5370, A2 => n4729, B1 => n5371, B2 => 
                           n4183, C1 => n5372, C2 => n4439, ZN => n5725);
   U689 : AOI221_X1 port map( B1 => n6788, B2 => n5373, C1 => n6692, C2 => 
                           n5374, A => n5726, ZN => n5723);
   U690 : OAI22_X1 port map( A1 => n5376, A2 => n4505, B1 => n5377, B2 => n4247
                           , ZN => n5726);
   U691 : AOI221_X1 port map( B1 => n6724, B2 => n5378, C1 => n6820, C2 => 
                           n5379, A => n5727, ZN => n5722);
   U692 : OAI222_X1 port map( A1 => n5381, A2 => n4697, B1 => n5382, B2 => 
                           n4215, C1 => n5383, C2 => n4471, ZN => n5727);
   U693 : AOI221_X1 port map( B1 => n6756, B2 => n5384, C1 => n6852, C2 => 
                           n5385, A => n5728, ZN => n5721);
   U694 : OAI22_X1 port map( A1 => n5387, A2 => n4569, B1 => n5388, B2 => n4311
                           , ZN => n5728);
   U695 : NAND4_X1 port map( A1 => n5729, A2 => n5730, A3 => n5731, A4 => n5732
                           , ZN => n4141);
   U696 : AOI221_X1 port map( B1 => n7002, B2 => n5343, C1 => n7066, C2 => 
                           n5344, A => n5733, ZN => n5732);
   U697 : OAI22_X1 port map( A1 => n5346, A2 => n4538, B1 => n5347, B2 => n4280
                           , ZN => n5733);
   U698 : AOI221_X1 port map( B1 => n6917, B2 => n5348, C1 => n7034, C2 => 
                           n5349, A => n5734, ZN => n5731);
   U699 : OAI22_X1 port map( A1 => n5351, A2 => n4666, B1 => n5352, B2 => n4408
                           , ZN => n5734);
   U700 : AOI221_X1 port map( B1 => n6970, B2 => n5353, C1 => n6938, C2 => 
                           n5354, A => n5735, ZN => n5730);
   U701 : OAI22_X1 port map( A1 => n5356, A2 => n4602, B1 => n5357, B2 => n4344
                           , ZN => n5735);
   U702 : AOI221_X1 port map( B1 => n5358, B2 => n5736, C1 => n5189, C2 => 
                           OUT1_10_port, A => n5737, ZN => n5729);
   U703 : OAI22_X1 port map( A1 => n5361, A2 => n4634, B1 => n5362, B2 => n4376
                           , ZN => n5737);
   U704 : NAND4_X1 port map( A1 => n5738, A2 => n5739, A3 => n5740, A4 => n5741
                           , ZN => n5736);
   U705 : AOI221_X1 port map( B1 => n6885, B2 => n5367, C1 => n6661, C2 => 
                           n5368, A => n5742, ZN => n5741);
   U706 : OAI222_X1 port map( A1 => n5370, A2 => n4730, B1 => n5371, B2 => 
                           n4184, C1 => n5372, C2 => n4440, ZN => n5742);
   U707 : AOI221_X1 port map( B1 => n6789, B2 => n5373, C1 => n6693, C2 => 
                           n5374, A => n5743, ZN => n5740);
   U708 : OAI22_X1 port map( A1 => n5376, A2 => n4506, B1 => n5377, B2 => n4248
                           , ZN => n5743);
   U709 : AOI221_X1 port map( B1 => n6725, B2 => n5378, C1 => n6821, C2 => 
                           n5379, A => n5744, ZN => n5739);
   U710 : OAI222_X1 port map( A1 => n5381, A2 => n4698, B1 => n5382, B2 => 
                           n4216, C1 => n5383, C2 => n4472, ZN => n5744);
   U711 : AOI221_X1 port map( B1 => n6757, B2 => n5384, C1 => n6853, C2 => 
                           n5385, A => n5745, ZN => n5738);
   U712 : OAI22_X1 port map( A1 => n5387, A2 => n4570, B1 => n5388, B2 => n4312
                           , ZN => n5745);
   U713 : NAND4_X1 port map( A1 => n5746, A2 => n5747, A3 => n5748, A4 => n5749
                           , ZN => n4140);
   U714 : AOI221_X1 port map( B1 => n7001, B2 => n5343, C1 => n7065, C2 => 
                           n5344, A => n5750, ZN => n5749);
   U715 : OAI22_X1 port map( A1 => n5346, A2 => n4539, B1 => n5347, B2 => n4281
                           , ZN => n5750);
   U716 : AOI221_X1 port map( B1 => n6918, B2 => n5348, C1 => n7033, C2 => 
                           n5349, A => n5751, ZN => n5748);
   U717 : OAI22_X1 port map( A1 => n5351, A2 => n4667, B1 => n5352, B2 => n4409
                           , ZN => n5751);
   U718 : AOI221_X1 port map( B1 => n6969, B2 => n5353, C1 => n6937, C2 => 
                           n5354, A => n5752, ZN => n5747);
   U719 : OAI22_X1 port map( A1 => n5356, A2 => n4603, B1 => n5357, B2 => n4345
                           , ZN => n5752);
   U720 : AOI221_X1 port map( B1 => n5358, B2 => n5753, C1 => n5189, C2 => 
                           OUT1_9_port, A => n5754, ZN => n5746);
   U721 : OAI22_X1 port map( A1 => n5361, A2 => n4635, B1 => n5362, B2 => n4377
                           , ZN => n5754);
   U722 : NAND4_X1 port map( A1 => n5755, A2 => n5756, A3 => n5757, A4 => n5758
                           , ZN => n5753);
   U723 : AOI221_X1 port map( B1 => n6886, B2 => n5367, C1 => n6662, C2 => 
                           n5368, A => n5759, ZN => n5758);
   U724 : OAI222_X1 port map( A1 => n5370, A2 => n4731, B1 => n5371, B2 => 
                           n4185, C1 => n5372, C2 => n4441, ZN => n5759);
   U725 : AOI221_X1 port map( B1 => n6790, B2 => n5373, C1 => n6694, C2 => 
                           n5374, A => n5760, ZN => n5757);
   U726 : OAI22_X1 port map( A1 => n5376, A2 => n4507, B1 => n5377, B2 => n4249
                           , ZN => n5760);
   U727 : AOI221_X1 port map( B1 => n6726, B2 => n5378, C1 => n6822, C2 => 
                           n5379, A => n5761, ZN => n5756);
   U728 : OAI222_X1 port map( A1 => n5381, A2 => n4699, B1 => n5382, B2 => 
                           n4217, C1 => n5383, C2 => n4473, ZN => n5761);
   U729 : AOI221_X1 port map( B1 => n6758, B2 => n5384, C1 => n6854, C2 => 
                           n5385, A => n5762, ZN => n5755);
   U730 : OAI22_X1 port map( A1 => n5387, A2 => n4571, B1 => n5388, B2 => n4313
                           , ZN => n5762);
   U731 : NAND4_X1 port map( A1 => n5763, A2 => n5764, A3 => n5765, A4 => n5766
                           , ZN => n4139);
   U732 : AOI221_X1 port map( B1 => n7000, B2 => n5343, C1 => n7064, C2 => 
                           n5344, A => n5767, ZN => n5766);
   U733 : OAI22_X1 port map( A1 => n5346, A2 => n4540, B1 => n5347, B2 => n4282
                           , ZN => n5767);
   U734 : AOI221_X1 port map( B1 => n6919, B2 => n5348, C1 => n7032, C2 => 
                           n5349, A => n5768, ZN => n5765);
   U735 : OAI22_X1 port map( A1 => n5351, A2 => n4668, B1 => n5352, B2 => n4410
                           , ZN => n5768);
   U736 : AOI221_X1 port map( B1 => n6968, B2 => n5353, C1 => n6936, C2 => 
                           n5354, A => n5769, ZN => n5764);
   U737 : OAI22_X1 port map( A1 => n5356, A2 => n4604, B1 => n5357, B2 => n4346
                           , ZN => n5769);
   U738 : AOI221_X1 port map( B1 => n5358, B2 => n5770, C1 => n5189, C2 => 
                           OUT1_8_port, A => n5771, ZN => n5763);
   U739 : OAI22_X1 port map( A1 => n5361, A2 => n4636, B1 => n5362, B2 => n4378
                           , ZN => n5771);
   U740 : NAND4_X1 port map( A1 => n5772, A2 => n5773, A3 => n5774, A4 => n5775
                           , ZN => n5770);
   U741 : AOI221_X1 port map( B1 => n6887, B2 => n5367, C1 => n6663, C2 => 
                           n5368, A => n5776, ZN => n5775);
   U742 : OAI222_X1 port map( A1 => n5370, A2 => n4732, B1 => n5371, B2 => 
                           n4186, C1 => n5372, C2 => n4442, ZN => n5776);
   U743 : AOI221_X1 port map( B1 => n6791, B2 => n5373, C1 => n6695, C2 => 
                           n5374, A => n5777, ZN => n5774);
   U744 : OAI22_X1 port map( A1 => n5376, A2 => n4508, B1 => n5377, B2 => n4250
                           , ZN => n5777);
   U745 : AOI221_X1 port map( B1 => n6727, B2 => n5378, C1 => n6823, C2 => 
                           n5379, A => n5778, ZN => n5773);
   U746 : OAI222_X1 port map( A1 => n5381, A2 => n4700, B1 => n5382, B2 => 
                           n4218, C1 => n5383, C2 => n4474, ZN => n5778);
   U747 : AOI221_X1 port map( B1 => n6759, B2 => n5384, C1 => n6855, C2 => 
                           n5385, A => n5779, ZN => n5772);
   U748 : OAI22_X1 port map( A1 => n5387, A2 => n4572, B1 => n5388, B2 => n4314
                           , ZN => n5779);
   U749 : NAND4_X1 port map( A1 => n5780, A2 => n5781, A3 => n5782, A4 => n5783
                           , ZN => n4138);
   U750 : AOI221_X1 port map( B1 => n6999, B2 => n5343, C1 => n7063, C2 => 
                           n5344, A => n5784, ZN => n5783);
   U751 : OAI22_X1 port map( A1 => n5346, A2 => n4541, B1 => n5347, B2 => n4283
                           , ZN => n5784);
   U752 : AOI221_X1 port map( B1 => n6920, B2 => n5348, C1 => n7031, C2 => 
                           n5349, A => n5785, ZN => n5782);
   U753 : OAI22_X1 port map( A1 => n5351, A2 => n4669, B1 => n5352, B2 => n4411
                           , ZN => n5785);
   U754 : AOI221_X1 port map( B1 => n6967, B2 => n5353, C1 => n6935, C2 => 
                           n5354, A => n5786, ZN => n5781);
   U755 : OAI22_X1 port map( A1 => n5356, A2 => n4605, B1 => n5357, B2 => n4347
                           , ZN => n5786);
   U756 : AOI221_X1 port map( B1 => n5358, B2 => n5787, C1 => n5189, C2 => 
                           OUT1_7_port, A => n5788, ZN => n5780);
   U757 : OAI22_X1 port map( A1 => n5361, A2 => n4637, B1 => n5362, B2 => n4379
                           , ZN => n5788);
   U758 : NAND4_X1 port map( A1 => n5789, A2 => n5790, A3 => n5791, A4 => n5792
                           , ZN => n5787);
   U759 : AOI221_X1 port map( B1 => n6888, B2 => n5367, C1 => n6664, C2 => 
                           n5368, A => n5793, ZN => n5792);
   U760 : OAI222_X1 port map( A1 => n5370, A2 => n4733, B1 => n5371, B2 => 
                           n4187, C1 => n5372, C2 => n4443, ZN => n5793);
   U761 : AOI221_X1 port map( B1 => n6792, B2 => n5373, C1 => n6696, C2 => 
                           n5374, A => n5794, ZN => n5791);
   U762 : OAI22_X1 port map( A1 => n5376, A2 => n4509, B1 => n5377, B2 => n4251
                           , ZN => n5794);
   U763 : AOI221_X1 port map( B1 => n6728, B2 => n5378, C1 => n6824, C2 => 
                           n5379, A => n5795, ZN => n5790);
   U764 : OAI222_X1 port map( A1 => n5381, A2 => n4701, B1 => n5382, B2 => 
                           n4219, C1 => n5383, C2 => n4475, ZN => n5795);
   U765 : AOI221_X1 port map( B1 => n6760, B2 => n5384, C1 => n6856, C2 => 
                           n5385, A => n5796, ZN => n5789);
   U766 : OAI22_X1 port map( A1 => n5387, A2 => n4573, B1 => n5388, B2 => n4315
                           , ZN => n5796);
   U767 : NAND4_X1 port map( A1 => n5797, A2 => n5798, A3 => n5799, A4 => n5800
                           , ZN => n4137);
   U768 : AOI221_X1 port map( B1 => n6998, B2 => n5343, C1 => n7062, C2 => 
                           n5344, A => n5801, ZN => n5800);
   U769 : OAI22_X1 port map( A1 => n5346, A2 => n4542, B1 => n5347, B2 => n4284
                           , ZN => n5801);
   U770 : AOI221_X1 port map( B1 => n6921, B2 => n5348, C1 => n7030, C2 => 
                           n5349, A => n5802, ZN => n5799);
   U771 : OAI22_X1 port map( A1 => n5351, A2 => n4670, B1 => n5352, B2 => n4412
                           , ZN => n5802);
   U772 : AOI221_X1 port map( B1 => n6966, B2 => n5353, C1 => n6934, C2 => 
                           n5354, A => n5803, ZN => n5798);
   U773 : OAI22_X1 port map( A1 => n5356, A2 => n4606, B1 => n5357, B2 => n4348
                           , ZN => n5803);
   U774 : AOI221_X1 port map( B1 => n5358, B2 => n5804, C1 => n5189, C2 => 
                           OUT1_6_port, A => n5805, ZN => n5797);
   U775 : OAI22_X1 port map( A1 => n5361, A2 => n4638, B1 => n5362, B2 => n4380
                           , ZN => n5805);
   U776 : NAND4_X1 port map( A1 => n5806, A2 => n5807, A3 => n5808, A4 => n5809
                           , ZN => n5804);
   U777 : AOI221_X1 port map( B1 => n6889, B2 => n5367, C1 => n6665, C2 => 
                           n5368, A => n5810, ZN => n5809);
   U778 : OAI222_X1 port map( A1 => n5370, A2 => n4734, B1 => n5371, B2 => 
                           n4188, C1 => n5372, C2 => n4444, ZN => n5810);
   U779 : AOI221_X1 port map( B1 => n6793, B2 => n5373, C1 => n6697, C2 => 
                           n5374, A => n5811, ZN => n5808);
   U780 : OAI22_X1 port map( A1 => n5376, A2 => n4510, B1 => n5377, B2 => n4252
                           , ZN => n5811);
   U781 : AOI221_X1 port map( B1 => n6729, B2 => n5378, C1 => n6825, C2 => 
                           n5379, A => n5812, ZN => n5807);
   U782 : OAI222_X1 port map( A1 => n5381, A2 => n4702, B1 => n5382, B2 => 
                           n4220, C1 => n5383, C2 => n4476, ZN => n5812);
   U783 : AOI221_X1 port map( B1 => n6761, B2 => n5384, C1 => n6857, C2 => 
                           n5385, A => n5813, ZN => n5806);
   U784 : OAI22_X1 port map( A1 => n5387, A2 => n4574, B1 => n5388, B2 => n4316
                           , ZN => n5813);
   U785 : NAND4_X1 port map( A1 => n5814, A2 => n5815, A3 => n5816, A4 => n5817
                           , ZN => n4136);
   U786 : AOI221_X1 port map( B1 => n6997, B2 => n5343, C1 => n7061, C2 => 
                           n5344, A => n5818, ZN => n5817);
   U787 : OAI22_X1 port map( A1 => n5346, A2 => n4543, B1 => n5347, B2 => n4285
                           , ZN => n5818);
   U788 : AOI221_X1 port map( B1 => n6922, B2 => n5348, C1 => n7029, C2 => 
                           n5349, A => n5819, ZN => n5816);
   U789 : OAI22_X1 port map( A1 => n5351, A2 => n4671, B1 => n5352, B2 => n4413
                           , ZN => n5819);
   U790 : AOI221_X1 port map( B1 => n6965, B2 => n5353, C1 => n6933, C2 => 
                           n5354, A => n5820, ZN => n5815);
   U791 : OAI22_X1 port map( A1 => n5356, A2 => n4607, B1 => n5357, B2 => n4349
                           , ZN => n5820);
   U792 : AOI221_X1 port map( B1 => n5358, B2 => n5821, C1 => n5189, C2 => 
                           OUT1_5_port, A => n5822, ZN => n5814);
   U793 : OAI22_X1 port map( A1 => n5361, A2 => n4639, B1 => n5362, B2 => n4381
                           , ZN => n5822);
   U794 : NAND4_X1 port map( A1 => n5823, A2 => n5824, A3 => n5825, A4 => n5826
                           , ZN => n5821);
   U795 : AOI221_X1 port map( B1 => n6890, B2 => n5367, C1 => n6666, C2 => 
                           n5368, A => n5827, ZN => n5826);
   U796 : OAI222_X1 port map( A1 => n5370, A2 => n4735, B1 => n5371, B2 => 
                           n4189, C1 => n5372, C2 => n4445, ZN => n5827);
   U797 : AOI221_X1 port map( B1 => n6794, B2 => n5373, C1 => n6698, C2 => 
                           n5374, A => n5828, ZN => n5825);
   U798 : OAI22_X1 port map( A1 => n5376, A2 => n4511, B1 => n5377, B2 => n4253
                           , ZN => n5828);
   U799 : AOI221_X1 port map( B1 => n6730, B2 => n5378, C1 => n6826, C2 => 
                           n5379, A => n5829, ZN => n5824);
   U800 : OAI222_X1 port map( A1 => n5381, A2 => n4703, B1 => n5382, B2 => 
                           n4221, C1 => n5383, C2 => n4477, ZN => n5829);
   U801 : AOI221_X1 port map( B1 => n6762, B2 => n5384, C1 => n6858, C2 => 
                           n5385, A => n5830, ZN => n5823);
   U802 : OAI22_X1 port map( A1 => n5387, A2 => n4575, B1 => n5388, B2 => n4317
                           , ZN => n5830);
   U803 : NAND4_X1 port map( A1 => n5831, A2 => n5832, A3 => n5833, A4 => n5834
                           , ZN => n4135);
   U804 : AOI221_X1 port map( B1 => n6996, B2 => n5343, C1 => n7060, C2 => 
                           n5344, A => n5835, ZN => n5834);
   U805 : OAI22_X1 port map( A1 => n5346, A2 => n4544, B1 => n5347, B2 => n4286
                           , ZN => n5835);
   U806 : AOI221_X1 port map( B1 => n6923, B2 => n5348, C1 => n7028, C2 => 
                           n5349, A => n5836, ZN => n5833);
   U807 : OAI22_X1 port map( A1 => n5351, A2 => n4672, B1 => n5352, B2 => n4414
                           , ZN => n5836);
   U808 : AOI221_X1 port map( B1 => n6964, B2 => n5353, C1 => n6932, C2 => 
                           n5354, A => n5837, ZN => n5832);
   U809 : OAI22_X1 port map( A1 => n5356, A2 => n4608, B1 => n5357, B2 => n4350
                           , ZN => n5837);
   U810 : AOI221_X1 port map( B1 => n5358, B2 => n5838, C1 => n5189, C2 => 
                           OUT1_4_port, A => n5839, ZN => n5831);
   U811 : OAI22_X1 port map( A1 => n5361, A2 => n4640, B1 => n5362, B2 => n4382
                           , ZN => n5839);
   U812 : NAND4_X1 port map( A1 => n5840, A2 => n5841, A3 => n5842, A4 => n5843
                           , ZN => n5838);
   U813 : AOI221_X1 port map( B1 => n6891, B2 => n5367, C1 => n6667, C2 => 
                           n5368, A => n5844, ZN => n5843);
   U814 : OAI222_X1 port map( A1 => n5370, A2 => n4736, B1 => n5371, B2 => 
                           n4190, C1 => n5372, C2 => n4446, ZN => n5844);
   U815 : AOI221_X1 port map( B1 => n6795, B2 => n5373, C1 => n6699, C2 => 
                           n5374, A => n5845, ZN => n5842);
   U816 : OAI22_X1 port map( A1 => n5376, A2 => n4512, B1 => n5377, B2 => n4254
                           , ZN => n5845);
   U817 : AOI221_X1 port map( B1 => n6731, B2 => n5378, C1 => n6827, C2 => 
                           n5379, A => n5846, ZN => n5841);
   U818 : OAI222_X1 port map( A1 => n5381, A2 => n4704, B1 => n5382, B2 => 
                           n4222, C1 => n5383, C2 => n4478, ZN => n5846);
   U819 : AOI221_X1 port map( B1 => n6763, B2 => n5384, C1 => n6859, C2 => 
                           n5385, A => n5847, ZN => n5840);
   U820 : OAI22_X1 port map( A1 => n5387, A2 => n4576, B1 => n5388, B2 => n4318
                           , ZN => n5847);
   U821 : NAND4_X1 port map( A1 => n5848, A2 => n5849, A3 => n5850, A4 => n5851
                           , ZN => n4134);
   U822 : AOI221_X1 port map( B1 => n6995, B2 => n5343, C1 => n7059, C2 => 
                           n5344, A => n5852, ZN => n5851);
   U823 : OAI22_X1 port map( A1 => n5346, A2 => n4545, B1 => n5347, B2 => n4287
                           , ZN => n5852);
   U824 : AOI221_X1 port map( B1 => n6924, B2 => n5348, C1 => n7027, C2 => 
                           n5349, A => n5853, ZN => n5850);
   U825 : OAI22_X1 port map( A1 => n5351, A2 => n4673, B1 => n5352, B2 => n4415
                           , ZN => n5853);
   U826 : AOI221_X1 port map( B1 => n6963, B2 => n5353, C1 => n6931, C2 => 
                           n5354, A => n5854, ZN => n5849);
   U827 : OAI22_X1 port map( A1 => n5356, A2 => n4609, B1 => n5357, B2 => n4351
                           , ZN => n5854);
   U828 : AOI221_X1 port map( B1 => n5358, B2 => n5855, C1 => n5189, C2 => 
                           OUT1_3_port, A => n5856, ZN => n5848);
   U829 : OAI22_X1 port map( A1 => n5361, A2 => n4641, B1 => n5362, B2 => n4383
                           , ZN => n5856);
   U830 : NAND4_X1 port map( A1 => n5857, A2 => n5858, A3 => n5859, A4 => n5860
                           , ZN => n5855);
   U831 : AOI221_X1 port map( B1 => n6892, B2 => n5367, C1 => n6668, C2 => 
                           n5368, A => n5861, ZN => n5860);
   U832 : OAI222_X1 port map( A1 => n5370, A2 => n4737, B1 => n5371, B2 => 
                           n4191, C1 => n5372, C2 => n4447, ZN => n5861);
   U833 : AOI221_X1 port map( B1 => n6796, B2 => n5373, C1 => n6700, C2 => 
                           n5374, A => n5862, ZN => n5859);
   U834 : OAI22_X1 port map( A1 => n5376, A2 => n4513, B1 => n5377, B2 => n4255
                           , ZN => n5862);
   U835 : AOI221_X1 port map( B1 => n6732, B2 => n5378, C1 => n6828, C2 => 
                           n5379, A => n5863, ZN => n5858);
   U836 : OAI222_X1 port map( A1 => n5381, A2 => n4705, B1 => n5382, B2 => 
                           n4223, C1 => n5383, C2 => n4479, ZN => n5863);
   U837 : AOI221_X1 port map( B1 => n6764, B2 => n5384, C1 => n6860, C2 => 
                           n5385, A => n5864, ZN => n5857);
   U838 : OAI22_X1 port map( A1 => n5387, A2 => n4577, B1 => n5388, B2 => n4319
                           , ZN => n5864);
   U839 : NAND4_X1 port map( A1 => n5865, A2 => n5866, A3 => n5867, A4 => n5868
                           , ZN => n4133);
   U840 : AOI221_X1 port map( B1 => n6994, B2 => n5343, C1 => n7058, C2 => 
                           n5344, A => n5869, ZN => n5868);
   U841 : OAI22_X1 port map( A1 => n5346, A2 => n4546, B1 => n5347, B2 => n4288
                           , ZN => n5869);
   U842 : AOI221_X1 port map( B1 => n6925, B2 => n5348, C1 => n7026, C2 => 
                           n5349, A => n5870, ZN => n5867);
   U843 : OAI22_X1 port map( A1 => n5351, A2 => n4674, B1 => n5352, B2 => n4416
                           , ZN => n5870);
   U844 : AOI221_X1 port map( B1 => n6962, B2 => n5353, C1 => n6930, C2 => 
                           n5354, A => n5871, ZN => n5866);
   U845 : OAI22_X1 port map( A1 => n5356, A2 => n4610, B1 => n5357, B2 => n4352
                           , ZN => n5871);
   U846 : AOI221_X1 port map( B1 => n5358, B2 => n5872, C1 => n5189, C2 => 
                           OUT1_2_port, A => n5873, ZN => n5865);
   U847 : OAI22_X1 port map( A1 => n5361, A2 => n4642, B1 => n5362, B2 => n4384
                           , ZN => n5873);
   U848 : NAND4_X1 port map( A1 => n5874, A2 => n5875, A3 => n5876, A4 => n5877
                           , ZN => n5872);
   U849 : AOI221_X1 port map( B1 => n6893, B2 => n5367, C1 => n6669, C2 => 
                           n5368, A => n5878, ZN => n5877);
   U850 : OAI222_X1 port map( A1 => n5370, A2 => n4738, B1 => n5371, B2 => 
                           n4192, C1 => n5372, C2 => n4448, ZN => n5878);
   U851 : AOI221_X1 port map( B1 => n6797, B2 => n5373, C1 => n6701, C2 => 
                           n5374, A => n5879, ZN => n5876);
   U852 : OAI22_X1 port map( A1 => n5376, A2 => n4514, B1 => n5377, B2 => n4256
                           , ZN => n5879);
   U853 : AOI221_X1 port map( B1 => n6733, B2 => n5378, C1 => n6829, C2 => 
                           n5379, A => n5880, ZN => n5875);
   U854 : OAI222_X1 port map( A1 => n5381, A2 => n4706, B1 => n5382, B2 => 
                           n4224, C1 => n5383, C2 => n4480, ZN => n5880);
   U855 : AOI221_X1 port map( B1 => n6765, B2 => n5384, C1 => n6861, C2 => 
                           n5385, A => n5881, ZN => n5874);
   U856 : OAI22_X1 port map( A1 => n5387, A2 => n4578, B1 => n5388, B2 => n4320
                           , ZN => n5881);
   U857 : NAND4_X1 port map( A1 => n5882, A2 => n5883, A3 => n5884, A4 => n5885
                           , ZN => n4132);
   U858 : AOI221_X1 port map( B1 => n6993, B2 => n5343, C1 => n7057, C2 => 
                           n5344, A => n5886, ZN => n5885);
   U859 : OAI22_X1 port map( A1 => n5346, A2 => n4547, B1 => n5347, B2 => n4289
                           , ZN => n5886);
   U860 : AOI221_X1 port map( B1 => n6926, B2 => n5348, C1 => n7025, C2 => 
                           n5349, A => n5887, ZN => n5884);
   U861 : OAI22_X1 port map( A1 => n5351, A2 => n4675, B1 => n5352, B2 => n4417
                           , ZN => n5887);
   U862 : AOI221_X1 port map( B1 => n6961, B2 => n5353, C1 => n6929, C2 => 
                           n5354, A => n5888, ZN => n5883);
   U863 : OAI22_X1 port map( A1 => n5356, A2 => n4611, B1 => n5357, B2 => n4353
                           , ZN => n5888);
   U864 : AOI221_X1 port map( B1 => n5358, B2 => n5889, C1 => n5189, C2 => 
                           OUT1_1_port, A => n5890, ZN => n5882);
   U865 : OAI22_X1 port map( A1 => n5361, A2 => n4643, B1 => n5362, B2 => n4385
                           , ZN => n5890);
   U866 : NAND4_X1 port map( A1 => n5891, A2 => n5892, A3 => n5893, A4 => n5894
                           , ZN => n5889);
   U867 : AOI221_X1 port map( B1 => n6894, B2 => n5367, C1 => n6670, C2 => 
                           n5368, A => n5895, ZN => n5894);
   U868 : OAI222_X1 port map( A1 => n5370, A2 => n4739, B1 => n5371, B2 => 
                           n4193, C1 => n5372, C2 => n4449, ZN => n5895);
   U869 : AOI221_X1 port map( B1 => n6798, B2 => n5373, C1 => n6702, C2 => 
                           n5374, A => n5896, ZN => n5893);
   U870 : OAI22_X1 port map( A1 => n5376, A2 => n4515, B1 => n5377, B2 => n4257
                           , ZN => n5896);
   U871 : AOI221_X1 port map( B1 => n6734, B2 => n5378, C1 => n6830, C2 => 
                           n5379, A => n5897, ZN => n5892);
   U872 : OAI222_X1 port map( A1 => n5381, A2 => n4707, B1 => n5382, B2 => 
                           n4225, C1 => n5383, C2 => n4481, ZN => n5897);
   U873 : AOI221_X1 port map( B1 => n6766, B2 => n5384, C1 => n6862, C2 => 
                           n5385, A => n5898, ZN => n5891);
   U874 : OAI22_X1 port map( A1 => n5387, A2 => n4579, B1 => n5388, B2 => n4321
                           , ZN => n5898);
   U875 : NAND4_X1 port map( A1 => n5899, A2 => n5900, A3 => n5901, A4 => n5902
                           , ZN => n4131);
   U876 : AOI221_X1 port map( B1 => n6992, B2 => n5343, C1 => n7056, C2 => 
                           n5344, A => n5903, ZN => n5902);
   U877 : OAI22_X1 port map( A1 => n5346, A2 => n4548, B1 => n5347, B2 => n4290
                           , ZN => n5903);
   U878 : AOI221_X1 port map( B1 => n6927, B2 => n5348, C1 => n7024, C2 => 
                           n5349, A => n5909, ZN => n5901);
   U879 : OAI22_X1 port map( A1 => n5351, A2 => n4676, B1 => n5352, B2 => n4418
                           , ZN => n5909);
   U880 : AND2_X1 port map( A1 => n5915, A2 => n5358, ZN => n5905);
   U881 : AOI221_X1 port map( B1 => n6960, B2 => n5353, C1 => n6928, C2 => 
                           n5354, A => n5916, ZN => n5900);
   U882 : OAI22_X1 port map( A1 => n5356, A2 => n4612, B1 => n5357, B2 => n4354
                           , ZN => n5916);
   U883 : AOI221_X1 port map( B1 => n5358, B2 => n5917, C1 => n5189, C2 => 
                           OUT1_0_port, A => n5918, ZN => n5899);
   U884 : OAI22_X1 port map( A1 => n5361, A2 => n4644, B1 => n5362, B2 => n4386
                           , ZN => n5918);
   U885 : AND3_X1 port map( A1 => n5358, A2 => ADD_RD1(4), A3 => ADD_RD1(3), ZN
                           => n5911);
   U886 : NAND4_X1 port map( A1 => n5919, A2 => n5920, A3 => n5921, A4 => n5922
                           , ZN => n5917);
   U887 : AOI221_X1 port map( B1 => n6895, B2 => n5367, C1 => n6671, C2 => 
                           n5368, A => n5923, ZN => n5922);
   U888 : OAI222_X1 port map( A1 => n5370, A2 => n4740, B1 => n5371, B2 => 
                           n4194, C1 => n5372, C2 => n4450, ZN => n5923);
   U889 : AOI221_X1 port map( B1 => n6799, B2 => n5373, C1 => n6703, C2 => 
                           n5374, A => n5926, ZN => n5921);
   U890 : OAI22_X1 port map( A1 => n5376, A2 => n4516, B1 => n5377, B2 => n4258
                           , ZN => n5926);
   U891 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n5927, ZN
                           => n5906);
   U892 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(0), ZN => n5907);
   U893 : AOI221_X1 port map( B1 => n6735, B2 => n5378, C1 => n6831, C2 => 
                           n5379, A => n5928, ZN => n5920);
   U894 : OAI222_X1 port map( A1 => n5381, A2 => n4708, B1 => n5382, B2 => 
                           n4226, C1 => n5383, C2 => n4482, ZN => n5928);
   U895 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n5929, ZN
                           => n5913);
   U896 : NOR3_X1 port map( A1 => n5929, A2 => ADD_RD1(0), A3 => n5930, ZN => 
                           n5908);
   U897 : NOR3_X1 port map( A1 => n5929, A2 => ADD_RD1(2), A3 => n5927, ZN => 
                           n5914);
   U898 : AOI221_X1 port map( B1 => n6767, B2 => n5384, C1 => n6863, C2 => 
                           n5385, A => n5931, ZN => n5919);
   U899 : OAI22_X1 port map( A1 => n5387, A2 => n4580, B1 => n5388, B2 => n4322
                           , ZN => n5931);
   U900 : NOR3_X1 port map( A1 => n5930, A2 => ADD_RD1(1), A3 => n5927, ZN => 
                           n5910);
   U901 : AND2_X1 port map( A1 => ADD_RD1(4), A2 => n5932, ZN => n5915);
   U902 : NOR3_X1 port map( A1 => n5930, A2 => n5929, A3 => n5927, ZN => n5912)
                           ;
   U903 : INV_X1 port map( A => ADD_RD1(0), ZN => n5927);
   U904 : INV_X1 port map( A => ADD_RD1(1), ZN => n5929);
   U905 : NOR2_X1 port map( A1 => n5932, A2 => ADD_RD1(4), ZN => n5925);
   U906 : INV_X1 port map( A => ADD_RD1(3), ZN => n5932);
   U907 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n5930, ZN
                           => n5904);
   U908 : INV_X1 port map( A => ADD_RD1(2), ZN => n5930);
   U909 : NOR2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n5924);
   U910 : NAND4_X1 port map( A1 => n5933, A2 => n5934, A3 => n5935, A4 => n5936
                           , ZN => n4130);
   U911 : AOI221_X1 port map( B1 => n5937, B2 => n7023, C1 => n5938, C2 => 
                           n7087, A => n5939, ZN => n5936);
   U912 : OAI22_X1 port map( A1 => n4517, A2 => n5940, B1 => n4259, B2 => n5941
                           , ZN => n5939);
   U913 : AOI221_X1 port map( B1 => n5942, B2 => n6896, C1 => n5943, C2 => 
                           n7055, A => n5944, ZN => n5935);
   U914 : OAI22_X1 port map( A1 => n4645, A2 => n5945, B1 => n4387, B2 => n5946
                           , ZN => n5944);
   U915 : AOI221_X1 port map( B1 => n5947, B2 => n6991, C1 => n5948, C2 => 
                           n6959, A => n5949, ZN => n5934);
   U916 : OAI22_X1 port map( A1 => n4581, A2 => n5950, B1 => n4323, B2 => n5951
                           , ZN => n5949);
   U917 : AOI221_X1 port map( B1 => n5952, B2 => n5953, C1 => n5190, C2 => 
                           OUT2_31_port, A => n5954, ZN => n5933);
   U918 : OAI22_X1 port map( A1 => n4613, A2 => n5955, B1 => n4355, B2 => n5956
                           , ZN => n5954);
   U919 : NAND4_X1 port map( A1 => n5957, A2 => n5958, A3 => n5959, A4 => n5960
                           , ZN => n5953);
   U920 : AOI221_X1 port map( B1 => n5961, B2 => n6864, C1 => n5962, C2 => 
                           n6640, A => n5963, ZN => n5960);
   U921 : OAI222_X1 port map( A1 => n4709, A2 => n5964, B1 => n4163, B2 => 
                           n5965, C1 => n4419, C2 => n5966, ZN => n5963);
   U922 : AOI221_X1 port map( B1 => n5967, B2 => n6768, C1 => n5968, C2 => 
                           n6672, A => n5969, ZN => n5959);
   U923 : OAI22_X1 port map( A1 => n4485, A2 => n5970, B1 => n4227, B2 => n5971
                           , ZN => n5969);
   U924 : AOI221_X1 port map( B1 => n5972, B2 => n6704, C1 => n5973, C2 => 
                           n6800, A => n5974, ZN => n5958);
   U925 : OAI222_X1 port map( A1 => n4677, A2 => n5975, B1 => n4195, B2 => 
                           n5976, C1 => n4451, C2 => n5977, ZN => n5974);
   U926 : AOI221_X1 port map( B1 => n5978, B2 => n6736, C1 => n5979, C2 => 
                           n6832, A => n5980, ZN => n5957);
   U927 : OAI22_X1 port map( A1 => n4549, A2 => n5981, B1 => n4291, B2 => n5982
                           , ZN => n5980);
   U928 : NAND4_X1 port map( A1 => n5983, A2 => n5984, A3 => n5985, A4 => n5986
                           , ZN => n4129);
   U929 : AOI221_X1 port map( B1 => n5937, B2 => n7022, C1 => n5938, C2 => 
                           n7086, A => n5987, ZN => n5986);
   U930 : OAI22_X1 port map( A1 => n4518, A2 => n5940, B1 => n4260, B2 => n5941
                           , ZN => n5987);
   U931 : AOI221_X1 port map( B1 => n5942, B2 => n6897, C1 => n5943, C2 => 
                           n7054, A => n5988, ZN => n5985);
   U932 : OAI22_X1 port map( A1 => n4646, A2 => n5945, B1 => n4388, B2 => n5946
                           , ZN => n5988);
   U933 : AOI221_X1 port map( B1 => n5947, B2 => n6990, C1 => n5948, C2 => 
                           n6958, A => n5989, ZN => n5984);
   U934 : OAI22_X1 port map( A1 => n4582, A2 => n5950, B1 => n4324, B2 => n5951
                           , ZN => n5989);
   U935 : AOI221_X1 port map( B1 => n5952, B2 => n5990, C1 => n5190, C2 => 
                           OUT2_30_port, A => n5991, ZN => n5983);
   U936 : OAI22_X1 port map( A1 => n4614, A2 => n5955, B1 => n4356, B2 => n5956
                           , ZN => n5991);
   U937 : NAND4_X1 port map( A1 => n5992, A2 => n5993, A3 => n5994, A4 => n5995
                           , ZN => n5990);
   U938 : AOI221_X1 port map( B1 => n5961, B2 => n6865, C1 => n5962, C2 => 
                           n6641, A => n5996, ZN => n5995);
   U939 : OAI222_X1 port map( A1 => n4710, A2 => n5964, B1 => n4164, B2 => 
                           n5965, C1 => n4420, C2 => n5966, ZN => n5996);
   U940 : AOI221_X1 port map( B1 => n5967, B2 => n6769, C1 => n5968, C2 => 
                           n6673, A => n5997, ZN => n5994);
   U941 : OAI22_X1 port map( A1 => n4486, A2 => n5970, B1 => n4228, B2 => n5971
                           , ZN => n5997);
   U942 : AOI221_X1 port map( B1 => n5972, B2 => n6705, C1 => n5973, C2 => 
                           n6801, A => n5998, ZN => n5993);
   U943 : OAI222_X1 port map( A1 => n4678, A2 => n5975, B1 => n4196, B2 => 
                           n5976, C1 => n4452, C2 => n5977, ZN => n5998);
   U944 : AOI221_X1 port map( B1 => n5978, B2 => n6737, C1 => n5979, C2 => 
                           n6833, A => n5999, ZN => n5992);
   U945 : OAI22_X1 port map( A1 => n4550, A2 => n5981, B1 => n4292, B2 => n5982
                           , ZN => n5999);
   U946 : NAND4_X1 port map( A1 => n6000, A2 => n6001, A3 => n6002, A4 => n6003
                           , ZN => n4128);
   U947 : AOI221_X1 port map( B1 => n5937, B2 => n7021, C1 => n5938, C2 => 
                           n7085, A => n6004, ZN => n6003);
   U948 : OAI22_X1 port map( A1 => n4519, A2 => n5940, B1 => n4261, B2 => n5941
                           , ZN => n6004);
   U949 : AOI221_X1 port map( B1 => n5942, B2 => n6898, C1 => n5943, C2 => 
                           n7053, A => n6005, ZN => n6002);
   U950 : OAI22_X1 port map( A1 => n4647, A2 => n5945, B1 => n4389, B2 => n5946
                           , ZN => n6005);
   U951 : AOI221_X1 port map( B1 => n5947, B2 => n6989, C1 => n5948, C2 => 
                           n6957, A => n6006, ZN => n6001);
   U952 : OAI22_X1 port map( A1 => n4583, A2 => n5950, B1 => n4325, B2 => n5951
                           , ZN => n6006);
   U953 : AOI221_X1 port map( B1 => n5952, B2 => n6007, C1 => n5190, C2 => 
                           OUT2_29_port, A => n6008, ZN => n6000);
   U954 : OAI22_X1 port map( A1 => n4615, A2 => n5955, B1 => n4357, B2 => n5956
                           , ZN => n6008);
   U955 : NAND4_X1 port map( A1 => n6009, A2 => n6010, A3 => n6011, A4 => n6012
                           , ZN => n6007);
   U956 : AOI221_X1 port map( B1 => n5961, B2 => n6866, C1 => n5962, C2 => 
                           n6642, A => n6013, ZN => n6012);
   U957 : OAI222_X1 port map( A1 => n4711, A2 => n5964, B1 => n4165, B2 => 
                           n5965, C1 => n4421, C2 => n5966, ZN => n6013);
   U958 : AOI221_X1 port map( B1 => n5967, B2 => n6770, C1 => n5968, C2 => 
                           n6674, A => n6014, ZN => n6011);
   U959 : OAI22_X1 port map( A1 => n4487, A2 => n5970, B1 => n4229, B2 => n5971
                           , ZN => n6014);
   U960 : AOI221_X1 port map( B1 => n5972, B2 => n6706, C1 => n5973, C2 => 
                           n6802, A => n6015, ZN => n6010);
   U961 : OAI222_X1 port map( A1 => n4679, A2 => n5975, B1 => n4197, B2 => 
                           n5976, C1 => n4453, C2 => n5977, ZN => n6015);
   U962 : AOI221_X1 port map( B1 => n5978, B2 => n6738, C1 => n5979, C2 => 
                           n6834, A => n6016, ZN => n6009);
   U963 : OAI22_X1 port map( A1 => n4551, A2 => n5981, B1 => n4293, B2 => n5982
                           , ZN => n6016);
   U964 : NAND4_X1 port map( A1 => n6017, A2 => n6018, A3 => n6019, A4 => n6020
                           , ZN => n4127);
   U965 : AOI221_X1 port map( B1 => n5937, B2 => n7020, C1 => n5938, C2 => 
                           n7084, A => n6021, ZN => n6020);
   U966 : OAI22_X1 port map( A1 => n4520, A2 => n5940, B1 => n4262, B2 => n5941
                           , ZN => n6021);
   U967 : AOI221_X1 port map( B1 => n5942, B2 => n6899, C1 => n5943, C2 => 
                           n7052, A => n6022, ZN => n6019);
   U968 : OAI22_X1 port map( A1 => n4648, A2 => n5945, B1 => n4390, B2 => n5946
                           , ZN => n6022);
   U969 : AOI221_X1 port map( B1 => n5947, B2 => n6988, C1 => n5948, C2 => 
                           n6956, A => n6023, ZN => n6018);
   U970 : OAI22_X1 port map( A1 => n4584, A2 => n5950, B1 => n4326, B2 => n5951
                           , ZN => n6023);
   U971 : AOI221_X1 port map( B1 => n5952, B2 => n6024, C1 => n5190, C2 => 
                           OUT2_28_port, A => n6025, ZN => n6017);
   U972 : OAI22_X1 port map( A1 => n4616, A2 => n5955, B1 => n4358, B2 => n5956
                           , ZN => n6025);
   U973 : NAND4_X1 port map( A1 => n6026, A2 => n6027, A3 => n6028, A4 => n6029
                           , ZN => n6024);
   U974 : AOI221_X1 port map( B1 => n5961, B2 => n6867, C1 => n5962, C2 => 
                           n6643, A => n6030, ZN => n6029);
   U975 : OAI222_X1 port map( A1 => n4712, A2 => n5964, B1 => n4166, B2 => 
                           n5965, C1 => n4422, C2 => n5966, ZN => n6030);
   U976 : AOI221_X1 port map( B1 => n5967, B2 => n6771, C1 => n5968, C2 => 
                           n6675, A => n6031, ZN => n6028);
   U977 : OAI22_X1 port map( A1 => n4488, A2 => n5970, B1 => n4230, B2 => n5971
                           , ZN => n6031);
   U978 : AOI221_X1 port map( B1 => n5972, B2 => n6707, C1 => n5973, C2 => 
                           n6803, A => n6032, ZN => n6027);
   U979 : OAI222_X1 port map( A1 => n4680, A2 => n5975, B1 => n4198, B2 => 
                           n5976, C1 => n4454, C2 => n5977, ZN => n6032);
   U980 : AOI221_X1 port map( B1 => n5978, B2 => n6739, C1 => n5979, C2 => 
                           n6835, A => n6033, ZN => n6026);
   U981 : OAI22_X1 port map( A1 => n4552, A2 => n5981, B1 => n4294, B2 => n5982
                           , ZN => n6033);
   U982 : NAND4_X1 port map( A1 => n6034, A2 => n6035, A3 => n6036, A4 => n6037
                           , ZN => n4126);
   U983 : AOI221_X1 port map( B1 => n5937, B2 => n7019, C1 => n5938, C2 => 
                           n7083, A => n6038, ZN => n6037);
   U984 : OAI22_X1 port map( A1 => n4521, A2 => n5940, B1 => n4263, B2 => n5941
                           , ZN => n6038);
   U985 : AOI221_X1 port map( B1 => n5942, B2 => n6900, C1 => n5943, C2 => 
                           n7051, A => n6039, ZN => n6036);
   U986 : OAI22_X1 port map( A1 => n4649, A2 => n5945, B1 => n4391, B2 => n5946
                           , ZN => n6039);
   U987 : AOI221_X1 port map( B1 => n5947, B2 => n6987, C1 => n5948, C2 => 
                           n6955, A => n6040, ZN => n6035);
   U988 : OAI22_X1 port map( A1 => n4585, A2 => n5950, B1 => n4327, B2 => n5951
                           , ZN => n6040);
   U989 : AOI221_X1 port map( B1 => n5952, B2 => n6041, C1 => n5190, C2 => 
                           OUT2_27_port, A => n6042, ZN => n6034);
   U990 : OAI22_X1 port map( A1 => n4617, A2 => n5955, B1 => n4359, B2 => n5956
                           , ZN => n6042);
   U991 : NAND4_X1 port map( A1 => n6043, A2 => n6044, A3 => n6045, A4 => n6046
                           , ZN => n6041);
   U992 : AOI221_X1 port map( B1 => n5961, B2 => n6868, C1 => n5962, C2 => 
                           n6644, A => n6047, ZN => n6046);
   U993 : OAI222_X1 port map( A1 => n4713, A2 => n5964, B1 => n4167, B2 => 
                           n5965, C1 => n4423, C2 => n5966, ZN => n6047);
   U994 : AOI221_X1 port map( B1 => n5967, B2 => n6772, C1 => n5968, C2 => 
                           n6676, A => n6048, ZN => n6045);
   U995 : OAI22_X1 port map( A1 => n4489, A2 => n5970, B1 => n4231, B2 => n5971
                           , ZN => n6048);
   U996 : AOI221_X1 port map( B1 => n5972, B2 => n6708, C1 => n5973, C2 => 
                           n6804, A => n6049, ZN => n6044);
   U997 : OAI222_X1 port map( A1 => n4681, A2 => n5975, B1 => n4199, B2 => 
                           n5976, C1 => n4455, C2 => n5977, ZN => n6049);
   U998 : AOI221_X1 port map( B1 => n5978, B2 => n6740, C1 => n5979, C2 => 
                           n6836, A => n6050, ZN => n6043);
   U999 : OAI22_X1 port map( A1 => n4553, A2 => n5981, B1 => n4295, B2 => n5982
                           , ZN => n6050);
   U1000 : NAND4_X1 port map( A1 => n6051, A2 => n6052, A3 => n6053, A4 => 
                           n6054, ZN => n4125);
   U1001 : AOI221_X1 port map( B1 => n5937, B2 => n7018, C1 => n5938, C2 => 
                           n7082, A => n6055, ZN => n6054);
   U1002 : OAI22_X1 port map( A1 => n4522, A2 => n5940, B1 => n4264, B2 => 
                           n5941, ZN => n6055);
   U1003 : AOI221_X1 port map( B1 => n5942, B2 => n6901, C1 => n5943, C2 => 
                           n7050, A => n6056, ZN => n6053);
   U1004 : OAI22_X1 port map( A1 => n4650, A2 => n5945, B1 => n4392, B2 => 
                           n5946, ZN => n6056);
   U1005 : AOI221_X1 port map( B1 => n5947, B2 => n6986, C1 => n5948, C2 => 
                           n6954, A => n6057, ZN => n6052);
   U1006 : OAI22_X1 port map( A1 => n4586, A2 => n5950, B1 => n4328, B2 => 
                           n5951, ZN => n6057);
   U1007 : AOI221_X1 port map( B1 => n5952, B2 => n6058, C1 => n5190, C2 => 
                           OUT2_26_port, A => n6059, ZN => n6051);
   U1008 : OAI22_X1 port map( A1 => n4618, A2 => n5955, B1 => n4360, B2 => 
                           n5956, ZN => n6059);
   U1009 : NAND4_X1 port map( A1 => n6060, A2 => n6061, A3 => n6062, A4 => 
                           n6063, ZN => n6058);
   U1010 : AOI221_X1 port map( B1 => n5961, B2 => n6869, C1 => n5962, C2 => 
                           n6645, A => n6064, ZN => n6063);
   U1011 : OAI222_X1 port map( A1 => n4714, A2 => n5964, B1 => n4168, B2 => 
                           n5965, C1 => n4424, C2 => n5966, ZN => n6064);
   U1012 : AOI221_X1 port map( B1 => n5967, B2 => n6773, C1 => n5968, C2 => 
                           n6677, A => n6065, ZN => n6062);
   U1013 : OAI22_X1 port map( A1 => n4490, A2 => n5970, B1 => n4232, B2 => 
                           n5971, ZN => n6065);
   U1014 : AOI221_X1 port map( B1 => n5972, B2 => n6709, C1 => n5973, C2 => 
                           n6805, A => n6066, ZN => n6061);
   U1015 : OAI222_X1 port map( A1 => n4682, A2 => n5975, B1 => n4200, B2 => 
                           n5976, C1 => n4456, C2 => n5977, ZN => n6066);
   U1016 : AOI221_X1 port map( B1 => n5978, B2 => n6741, C1 => n5979, C2 => 
                           n6837, A => n6067, ZN => n6060);
   U1017 : OAI22_X1 port map( A1 => n4554, A2 => n5981, B1 => n4296, B2 => 
                           n5982, ZN => n6067);
   U1018 : NAND4_X1 port map( A1 => n6068, A2 => n6069, A3 => n6070, A4 => 
                           n6071, ZN => n4124);
   U1019 : AOI221_X1 port map( B1 => n5937, B2 => n7017, C1 => n5938, C2 => 
                           n7081, A => n6072, ZN => n6071);
   U1020 : OAI22_X1 port map( A1 => n4523, A2 => n5940, B1 => n4265, B2 => 
                           n5941, ZN => n6072);
   U1021 : AOI221_X1 port map( B1 => n5942, B2 => n6902, C1 => n5943, C2 => 
                           n7049, A => n6073, ZN => n6070);
   U1022 : OAI22_X1 port map( A1 => n4651, A2 => n5945, B1 => n4393, B2 => 
                           n5946, ZN => n6073);
   U1023 : AOI221_X1 port map( B1 => n5947, B2 => n6985, C1 => n5948, C2 => 
                           n6953, A => n6074, ZN => n6069);
   U1024 : OAI22_X1 port map( A1 => n4587, A2 => n5950, B1 => n4329, B2 => 
                           n5951, ZN => n6074);
   U1025 : AOI221_X1 port map( B1 => n5952, B2 => n6075, C1 => n5190, C2 => 
                           OUT2_25_port, A => n6076, ZN => n6068);
   U1026 : OAI22_X1 port map( A1 => n4619, A2 => n5955, B1 => n4361, B2 => 
                           n5956, ZN => n6076);
   U1027 : NAND4_X1 port map( A1 => n6077, A2 => n6078, A3 => n6079, A4 => 
                           n6080, ZN => n6075);
   U1028 : AOI221_X1 port map( B1 => n5961, B2 => n6870, C1 => n5962, C2 => 
                           n6646, A => n6081, ZN => n6080);
   U1029 : OAI222_X1 port map( A1 => n4715, A2 => n5964, B1 => n4169, B2 => 
                           n5965, C1 => n4425, C2 => n5966, ZN => n6081);
   U1030 : AOI221_X1 port map( B1 => n5967, B2 => n6774, C1 => n5968, C2 => 
                           n6678, A => n6082, ZN => n6079);
   U1031 : OAI22_X1 port map( A1 => n4491, A2 => n5970, B1 => n4233, B2 => 
                           n5971, ZN => n6082);
   U1032 : AOI221_X1 port map( B1 => n5972, B2 => n6710, C1 => n5973, C2 => 
                           n6806, A => n6083, ZN => n6078);
   U1033 : OAI222_X1 port map( A1 => n4683, A2 => n5975, B1 => n4201, B2 => 
                           n5976, C1 => n4457, C2 => n5977, ZN => n6083);
   U1034 : AOI221_X1 port map( B1 => n5978, B2 => n6742, C1 => n5979, C2 => 
                           n6838, A => n6084, ZN => n6077);
   U1035 : OAI22_X1 port map( A1 => n4555, A2 => n5981, B1 => n4297, B2 => 
                           n5982, ZN => n6084);
   U1036 : NAND4_X1 port map( A1 => n6085, A2 => n6086, A3 => n6087, A4 => 
                           n6088, ZN => n4123);
   U1037 : AOI221_X1 port map( B1 => n5937, B2 => n7016, C1 => n5938, C2 => 
                           n7080, A => n6089, ZN => n6088);
   U1038 : OAI22_X1 port map( A1 => n4524, A2 => n5940, B1 => n4266, B2 => 
                           n5941, ZN => n6089);
   U1039 : AOI221_X1 port map( B1 => n5942, B2 => n6903, C1 => n5943, C2 => 
                           n7048, A => n6090, ZN => n6087);
   U1040 : OAI22_X1 port map( A1 => n4652, A2 => n5945, B1 => n4394, B2 => 
                           n5946, ZN => n6090);
   U1041 : AOI221_X1 port map( B1 => n5947, B2 => n6984, C1 => n5948, C2 => 
                           n6952, A => n6091, ZN => n6086);
   U1042 : OAI22_X1 port map( A1 => n4588, A2 => n5950, B1 => n4330, B2 => 
                           n5951, ZN => n6091);
   U1043 : AOI221_X1 port map( B1 => n5952, B2 => n6092, C1 => n5190, C2 => 
                           OUT2_24_port, A => n6093, ZN => n6085);
   U1044 : OAI22_X1 port map( A1 => n4620, A2 => n5955, B1 => n4362, B2 => 
                           n5956, ZN => n6093);
   U1045 : NAND4_X1 port map( A1 => n6094, A2 => n6095, A3 => n6096, A4 => 
                           n6097, ZN => n6092);
   U1046 : AOI221_X1 port map( B1 => n5961, B2 => n6871, C1 => n5962, C2 => 
                           n6647, A => n6098, ZN => n6097);
   U1047 : OAI222_X1 port map( A1 => n4716, A2 => n5964, B1 => n4170, B2 => 
                           n5965, C1 => n4426, C2 => n5966, ZN => n6098);
   U1048 : AOI221_X1 port map( B1 => n5967, B2 => n6775, C1 => n5968, C2 => 
                           n6679, A => n6099, ZN => n6096);
   U1049 : OAI22_X1 port map( A1 => n4492, A2 => n5970, B1 => n4234, B2 => 
                           n5971, ZN => n6099);
   U1050 : AOI221_X1 port map( B1 => n5972, B2 => n6711, C1 => n5973, C2 => 
                           n6807, A => n6100, ZN => n6095);
   U1051 : OAI222_X1 port map( A1 => n4684, A2 => n5975, B1 => n4202, B2 => 
                           n5976, C1 => n4458, C2 => n5977, ZN => n6100);
   U1052 : AOI221_X1 port map( B1 => n5978, B2 => n6743, C1 => n5979, C2 => 
                           n6839, A => n6101, ZN => n6094);
   U1053 : OAI22_X1 port map( A1 => n4556, A2 => n5981, B1 => n4298, B2 => 
                           n5982, ZN => n6101);
   U1054 : NAND4_X1 port map( A1 => n6102, A2 => n6103, A3 => n6104, A4 => 
                           n6105, ZN => n4122);
   U1055 : AOI221_X1 port map( B1 => n5937, B2 => n7015, C1 => n5938, C2 => 
                           n7079, A => n6106, ZN => n6105);
   U1056 : OAI22_X1 port map( A1 => n4525, A2 => n5940, B1 => n4267, B2 => 
                           n5941, ZN => n6106);
   U1057 : AOI221_X1 port map( B1 => n5942, B2 => n6904, C1 => n5943, C2 => 
                           n7047, A => n6107, ZN => n6104);
   U1058 : OAI22_X1 port map( A1 => n4653, A2 => n5945, B1 => n4395, B2 => 
                           n5946, ZN => n6107);
   U1059 : AOI221_X1 port map( B1 => n5947, B2 => n6983, C1 => n5948, C2 => 
                           n6951, A => n6108, ZN => n6103);
   U1060 : OAI22_X1 port map( A1 => n4589, A2 => n5950, B1 => n4331, B2 => 
                           n5951, ZN => n6108);
   U1061 : AOI221_X1 port map( B1 => n5952, B2 => n6109, C1 => n5190, C2 => 
                           OUT2_23_port, A => n6110, ZN => n6102);
   U1062 : OAI22_X1 port map( A1 => n4621, A2 => n5955, B1 => n4363, B2 => 
                           n5956, ZN => n6110);
   U1063 : NAND4_X1 port map( A1 => n6111, A2 => n6112, A3 => n6113, A4 => 
                           n6114, ZN => n6109);
   U1064 : AOI221_X1 port map( B1 => n5961, B2 => n6872, C1 => n5962, C2 => 
                           n6648, A => n6115, ZN => n6114);
   U1065 : OAI222_X1 port map( A1 => n4717, A2 => n5964, B1 => n4171, B2 => 
                           n5965, C1 => n4427, C2 => n5966, ZN => n6115);
   U1066 : AOI221_X1 port map( B1 => n5967, B2 => n6776, C1 => n5968, C2 => 
                           n6680, A => n6116, ZN => n6113);
   U1067 : OAI22_X1 port map( A1 => n4493, A2 => n5970, B1 => n4235, B2 => 
                           n5971, ZN => n6116);
   U1068 : AOI221_X1 port map( B1 => n5972, B2 => n6712, C1 => n5973, C2 => 
                           n6808, A => n6117, ZN => n6112);
   U1069 : OAI222_X1 port map( A1 => n4685, A2 => n5975, B1 => n4203, B2 => 
                           n5976, C1 => n4459, C2 => n5977, ZN => n6117);
   U1070 : AOI221_X1 port map( B1 => n5978, B2 => n6744, C1 => n5979, C2 => 
                           n6840, A => n6118, ZN => n6111);
   U1071 : OAI22_X1 port map( A1 => n4557, A2 => n5981, B1 => n4299, B2 => 
                           n5982, ZN => n6118);
   U1072 : NAND4_X1 port map( A1 => n6119, A2 => n6120, A3 => n6121, A4 => 
                           n6122, ZN => n4121);
   U1073 : AOI221_X1 port map( B1 => n5937, B2 => n7014, C1 => n5938, C2 => 
                           n7078, A => n6123, ZN => n6122);
   U1074 : OAI22_X1 port map( A1 => n4526, A2 => n5940, B1 => n4268, B2 => 
                           n5941, ZN => n6123);
   U1075 : AOI221_X1 port map( B1 => n5942, B2 => n6905, C1 => n5943, C2 => 
                           n7046, A => n6124, ZN => n6121);
   U1076 : OAI22_X1 port map( A1 => n4654, A2 => n5945, B1 => n4396, B2 => 
                           n5946, ZN => n6124);
   U1077 : AOI221_X1 port map( B1 => n5947, B2 => n6982, C1 => n5948, C2 => 
                           n6950, A => n6125, ZN => n6120);
   U1078 : OAI22_X1 port map( A1 => n4590, A2 => n5950, B1 => n4332, B2 => 
                           n5951, ZN => n6125);
   U1079 : AOI221_X1 port map( B1 => n5952, B2 => n6126, C1 => n5190, C2 => 
                           OUT2_22_port, A => n6127, ZN => n6119);
   U1080 : OAI22_X1 port map( A1 => n4622, A2 => n5955, B1 => n4364, B2 => 
                           n5956, ZN => n6127);
   U1081 : NAND4_X1 port map( A1 => n6128, A2 => n6129, A3 => n6130, A4 => 
                           n6131, ZN => n6126);
   U1082 : AOI221_X1 port map( B1 => n5961, B2 => n6873, C1 => n5962, C2 => 
                           n6649, A => n6132, ZN => n6131);
   U1083 : OAI222_X1 port map( A1 => n4718, A2 => n5964, B1 => n4172, B2 => 
                           n5965, C1 => n4428, C2 => n5966, ZN => n6132);
   U1084 : AOI221_X1 port map( B1 => n5967, B2 => n6777, C1 => n5968, C2 => 
                           n6681, A => n6133, ZN => n6130);
   U1085 : OAI22_X1 port map( A1 => n4494, A2 => n5970, B1 => n4236, B2 => 
                           n5971, ZN => n6133);
   U1086 : AOI221_X1 port map( B1 => n5972, B2 => n6713, C1 => n5973, C2 => 
                           n6809, A => n6134, ZN => n6129);
   U1087 : OAI222_X1 port map( A1 => n4686, A2 => n5975, B1 => n4204, B2 => 
                           n5976, C1 => n4460, C2 => n5977, ZN => n6134);
   U1088 : AOI221_X1 port map( B1 => n5978, B2 => n6745, C1 => n5979, C2 => 
                           n6841, A => n6135, ZN => n6128);
   U1089 : OAI22_X1 port map( A1 => n4558, A2 => n5981, B1 => n4300, B2 => 
                           n5982, ZN => n6135);
   U1090 : NAND4_X1 port map( A1 => n6136, A2 => n6137, A3 => n6138, A4 => 
                           n6139, ZN => n4120);
   U1091 : AOI221_X1 port map( B1 => n5937, B2 => n7013, C1 => n5938, C2 => 
                           n7077, A => n6140, ZN => n6139);
   U1092 : OAI22_X1 port map( A1 => n4527, A2 => n5940, B1 => n4269, B2 => 
                           n5941, ZN => n6140);
   U1093 : AOI221_X1 port map( B1 => n5942, B2 => n6906, C1 => n5943, C2 => 
                           n7045, A => n6141, ZN => n6138);
   U1094 : OAI22_X1 port map( A1 => n4655, A2 => n5945, B1 => n4397, B2 => 
                           n5946, ZN => n6141);
   U1095 : AOI221_X1 port map( B1 => n5947, B2 => n6981, C1 => n5948, C2 => 
                           n6949, A => n6142, ZN => n6137);
   U1096 : OAI22_X1 port map( A1 => n4591, A2 => n5950, B1 => n4333, B2 => 
                           n5951, ZN => n6142);
   U1097 : AOI221_X1 port map( B1 => n5952, B2 => n6143, C1 => n5190, C2 => 
                           OUT2_21_port, A => n6144, ZN => n6136);
   U1098 : OAI22_X1 port map( A1 => n4623, A2 => n5955, B1 => n4365, B2 => 
                           n5956, ZN => n6144);
   U1099 : NAND4_X1 port map( A1 => n6145, A2 => n6146, A3 => n6147, A4 => 
                           n6148, ZN => n6143);
   U1100 : AOI221_X1 port map( B1 => n5961, B2 => n6874, C1 => n5962, C2 => 
                           n6650, A => n6149, ZN => n6148);
   U1101 : OAI222_X1 port map( A1 => n4719, A2 => n5964, B1 => n4173, B2 => 
                           n5965, C1 => n4429, C2 => n5966, ZN => n6149);
   U1102 : AOI221_X1 port map( B1 => n5967, B2 => n6778, C1 => n5968, C2 => 
                           n6682, A => n6150, ZN => n6147);
   U1103 : OAI22_X1 port map( A1 => n4495, A2 => n5970, B1 => n4237, B2 => 
                           n5971, ZN => n6150);
   U1104 : AOI221_X1 port map( B1 => n5972, B2 => n6714, C1 => n5973, C2 => 
                           n6810, A => n6151, ZN => n6146);
   U1105 : OAI222_X1 port map( A1 => n4687, A2 => n5975, B1 => n4205, B2 => 
                           n5976, C1 => n4461, C2 => n5977, ZN => n6151);
   U1106 : AOI221_X1 port map( B1 => n5978, B2 => n6746, C1 => n5979, C2 => 
                           n6842, A => n6152, ZN => n6145);
   U1107 : OAI22_X1 port map( A1 => n4559, A2 => n5981, B1 => n4301, B2 => 
                           n5982, ZN => n6152);
   U1108 : NAND4_X1 port map( A1 => n6153, A2 => n6154, A3 => n6155, A4 => 
                           n6156, ZN => n4119);
   U1109 : AOI221_X1 port map( B1 => n5937, B2 => n7012, C1 => n5938, C2 => 
                           n7076, A => n6157, ZN => n6156);
   U1110 : OAI22_X1 port map( A1 => n4528, A2 => n5940, B1 => n4270, B2 => 
                           n5941, ZN => n6157);
   U1111 : AOI221_X1 port map( B1 => n5942, B2 => n6907, C1 => n5943, C2 => 
                           n7044, A => n6158, ZN => n6155);
   U1112 : OAI22_X1 port map( A1 => n4656, A2 => n5945, B1 => n4398, B2 => 
                           n5946, ZN => n6158);
   U1113 : AOI221_X1 port map( B1 => n5947, B2 => n6980, C1 => n5948, C2 => 
                           n6948, A => n6159, ZN => n6154);
   U1114 : OAI22_X1 port map( A1 => n4592, A2 => n5950, B1 => n4334, B2 => 
                           n5951, ZN => n6159);
   U1115 : AOI221_X1 port map( B1 => n5952, B2 => n6160, C1 => n5190, C2 => 
                           OUT2_20_port, A => n6161, ZN => n6153);
   U1116 : OAI22_X1 port map( A1 => n4624, A2 => n5955, B1 => n4366, B2 => 
                           n5956, ZN => n6161);
   U1117 : NAND4_X1 port map( A1 => n6162, A2 => n6163, A3 => n6164, A4 => 
                           n6165, ZN => n6160);
   U1118 : AOI221_X1 port map( B1 => n5961, B2 => n6875, C1 => n5962, C2 => 
                           n6651, A => n6166, ZN => n6165);
   U1119 : OAI222_X1 port map( A1 => n4720, A2 => n5964, B1 => n4174, B2 => 
                           n5965, C1 => n4430, C2 => n5966, ZN => n6166);
   U1120 : AOI221_X1 port map( B1 => n5967, B2 => n6779, C1 => n5968, C2 => 
                           n6683, A => n6167, ZN => n6164);
   U1121 : OAI22_X1 port map( A1 => n4496, A2 => n5970, B1 => n4238, B2 => 
                           n5971, ZN => n6167);
   U1122 : AOI221_X1 port map( B1 => n5972, B2 => n6715, C1 => n5973, C2 => 
                           n6811, A => n6168, ZN => n6163);
   U1123 : OAI222_X1 port map( A1 => n4688, A2 => n5975, B1 => n4206, B2 => 
                           n5976, C1 => n4462, C2 => n5977, ZN => n6168);
   U1124 : AOI221_X1 port map( B1 => n5978, B2 => n6747, C1 => n5979, C2 => 
                           n6843, A => n6169, ZN => n6162);
   U1125 : OAI22_X1 port map( A1 => n4560, A2 => n5981, B1 => n4302, B2 => 
                           n5982, ZN => n6169);
   U1126 : NAND4_X1 port map( A1 => n6170, A2 => n6171, A3 => n6172, A4 => 
                           n6173, ZN => n4118);
   U1127 : AOI221_X1 port map( B1 => n5937, B2 => n7011, C1 => n5938, C2 => 
                           n7075, A => n6174, ZN => n6173);
   U1128 : OAI22_X1 port map( A1 => n4529, A2 => n5940, B1 => n4271, B2 => 
                           n5941, ZN => n6174);
   U1129 : AOI221_X1 port map( B1 => n5942, B2 => n6908, C1 => n5943, C2 => 
                           n7043, A => n6175, ZN => n6172);
   U1130 : OAI22_X1 port map( A1 => n4657, A2 => n5945, B1 => n4399, B2 => 
                           n5946, ZN => n6175);
   U1131 : AOI221_X1 port map( B1 => n5947, B2 => n6979, C1 => n5948, C2 => 
                           n6947, A => n6176, ZN => n6171);
   U1132 : OAI22_X1 port map( A1 => n4593, A2 => n5950, B1 => n4335, B2 => 
                           n5951, ZN => n6176);
   U1133 : AOI221_X1 port map( B1 => n5952, B2 => n6177, C1 => n5190, C2 => 
                           OUT2_19_port, A => n6178, ZN => n6170);
   U1134 : OAI22_X1 port map( A1 => n4625, A2 => n5955, B1 => n4367, B2 => 
                           n5956, ZN => n6178);
   U1135 : NAND4_X1 port map( A1 => n6179, A2 => n6180, A3 => n6181, A4 => 
                           n6182, ZN => n6177);
   U1136 : AOI221_X1 port map( B1 => n5961, B2 => n6876, C1 => n5962, C2 => 
                           n6652, A => n6183, ZN => n6182);
   U1137 : OAI222_X1 port map( A1 => n4721, A2 => n5964, B1 => n4175, B2 => 
                           n5965, C1 => n4431, C2 => n5966, ZN => n6183);
   U1138 : AOI221_X1 port map( B1 => n5967, B2 => n6780, C1 => n5968, C2 => 
                           n6684, A => n6184, ZN => n6181);
   U1139 : OAI22_X1 port map( A1 => n4497, A2 => n5970, B1 => n4239, B2 => 
                           n5971, ZN => n6184);
   U1140 : AOI221_X1 port map( B1 => n5972, B2 => n6716, C1 => n5973, C2 => 
                           n6812, A => n6185, ZN => n6180);
   U1141 : OAI222_X1 port map( A1 => n4689, A2 => n5975, B1 => n4207, B2 => 
                           n5976, C1 => n4463, C2 => n5977, ZN => n6185);
   U1142 : AOI221_X1 port map( B1 => n5978, B2 => n6748, C1 => n5979, C2 => 
                           n6844, A => n6186, ZN => n6179);
   U1143 : OAI22_X1 port map( A1 => n4561, A2 => n5981, B1 => n4303, B2 => 
                           n5982, ZN => n6186);
   U1144 : NAND4_X1 port map( A1 => n6187, A2 => n6188, A3 => n6189, A4 => 
                           n6190, ZN => n4117);
   U1145 : AOI221_X1 port map( B1 => n5937, B2 => n7010, C1 => n5938, C2 => 
                           n7074, A => n6191, ZN => n6190);
   U1146 : OAI22_X1 port map( A1 => n4530, A2 => n5940, B1 => n4272, B2 => 
                           n5941, ZN => n6191);
   U1147 : AOI221_X1 port map( B1 => n5942, B2 => n6909, C1 => n5943, C2 => 
                           n7042, A => n6192, ZN => n6189);
   U1148 : OAI22_X1 port map( A1 => n4658, A2 => n5945, B1 => n4400, B2 => 
                           n5946, ZN => n6192);
   U1149 : AOI221_X1 port map( B1 => n5947, B2 => n6978, C1 => n5948, C2 => 
                           n6946, A => n6193, ZN => n6188);
   U1150 : OAI22_X1 port map( A1 => n4594, A2 => n5950, B1 => n4336, B2 => 
                           n5951, ZN => n6193);
   U1151 : AOI221_X1 port map( B1 => n5952, B2 => n6194, C1 => n5190, C2 => 
                           OUT2_18_port, A => n6195, ZN => n6187);
   U1152 : OAI22_X1 port map( A1 => n4626, A2 => n5955, B1 => n4368, B2 => 
                           n5956, ZN => n6195);
   U1153 : NAND4_X1 port map( A1 => n6196, A2 => n6197, A3 => n6198, A4 => 
                           n6199, ZN => n6194);
   U1154 : AOI221_X1 port map( B1 => n5961, B2 => n6877, C1 => n5962, C2 => 
                           n6653, A => n6200, ZN => n6199);
   U1155 : OAI222_X1 port map( A1 => n4722, A2 => n5964, B1 => n4176, B2 => 
                           n5965, C1 => n4432, C2 => n5966, ZN => n6200);
   U1156 : AOI221_X1 port map( B1 => n5967, B2 => n6781, C1 => n5968, C2 => 
                           n6685, A => n6201, ZN => n6198);
   U1157 : OAI22_X1 port map( A1 => n4498, A2 => n5970, B1 => n4240, B2 => 
                           n5971, ZN => n6201);
   U1158 : AOI221_X1 port map( B1 => n5972, B2 => n6717, C1 => n5973, C2 => 
                           n6813, A => n6202, ZN => n6197);
   U1159 : OAI222_X1 port map( A1 => n4690, A2 => n5975, B1 => n4208, B2 => 
                           n5976, C1 => n4464, C2 => n5977, ZN => n6202);
   U1160 : AOI221_X1 port map( B1 => n5978, B2 => n6749, C1 => n5979, C2 => 
                           n6845, A => n6203, ZN => n6196);
   U1161 : OAI22_X1 port map( A1 => n4562, A2 => n5981, B1 => n4304, B2 => 
                           n5982, ZN => n6203);
   U1162 : NAND4_X1 port map( A1 => n6204, A2 => n6205, A3 => n6206, A4 => 
                           n6207, ZN => n4116);
   U1163 : AOI221_X1 port map( B1 => n5937, B2 => n7009, C1 => n5938, C2 => 
                           n7073, A => n6208, ZN => n6207);
   U1164 : OAI22_X1 port map( A1 => n4531, A2 => n5940, B1 => n4273, B2 => 
                           n5941, ZN => n6208);
   U1165 : AOI221_X1 port map( B1 => n5942, B2 => n6910, C1 => n5943, C2 => 
                           n7041, A => n6209, ZN => n6206);
   U1166 : OAI22_X1 port map( A1 => n4659, A2 => n5945, B1 => n4401, B2 => 
                           n5946, ZN => n6209);
   U1167 : AOI221_X1 port map( B1 => n5947, B2 => n6977, C1 => n5948, C2 => 
                           n6945, A => n6210, ZN => n6205);
   U1168 : OAI22_X1 port map( A1 => n4595, A2 => n5950, B1 => n4337, B2 => 
                           n5951, ZN => n6210);
   U1169 : AOI221_X1 port map( B1 => n5952, B2 => n6211, C1 => n5190, C2 => 
                           OUT2_17_port, A => n6212, ZN => n6204);
   U1170 : OAI22_X1 port map( A1 => n4627, A2 => n5955, B1 => n4369, B2 => 
                           n5956, ZN => n6212);
   U1171 : NAND4_X1 port map( A1 => n6213, A2 => n6214, A3 => n6215, A4 => 
                           n6216, ZN => n6211);
   U1172 : AOI221_X1 port map( B1 => n5961, B2 => n6878, C1 => n5962, C2 => 
                           n6654, A => n6217, ZN => n6216);
   U1173 : OAI222_X1 port map( A1 => n4723, A2 => n5964, B1 => n4177, B2 => 
                           n5965, C1 => n4433, C2 => n5966, ZN => n6217);
   U1174 : AOI221_X1 port map( B1 => n5967, B2 => n6782, C1 => n5968, C2 => 
                           n6686, A => n6218, ZN => n6215);
   U1175 : OAI22_X1 port map( A1 => n4499, A2 => n5970, B1 => n4241, B2 => 
                           n5971, ZN => n6218);
   U1176 : AOI221_X1 port map( B1 => n5972, B2 => n6718, C1 => n5973, C2 => 
                           n6814, A => n6219, ZN => n6214);
   U1177 : OAI222_X1 port map( A1 => n4691, A2 => n5975, B1 => n4209, B2 => 
                           n5976, C1 => n4465, C2 => n5977, ZN => n6219);
   U1178 : AOI221_X1 port map( B1 => n5978, B2 => n6750, C1 => n5979, C2 => 
                           n6846, A => n6220, ZN => n6213);
   U1179 : OAI22_X1 port map( A1 => n4563, A2 => n5981, B1 => n4305, B2 => 
                           n5982, ZN => n6220);
   U1180 : NAND4_X1 port map( A1 => n6221, A2 => n6222, A3 => n6223, A4 => 
                           n6224, ZN => n4115);
   U1181 : AOI221_X1 port map( B1 => n5937, B2 => n7008, C1 => n5938, C2 => 
                           n7072, A => n6225, ZN => n6224);
   U1182 : OAI22_X1 port map( A1 => n4532, A2 => n5940, B1 => n4274, B2 => 
                           n5941, ZN => n6225);
   U1183 : AOI221_X1 port map( B1 => n5942, B2 => n6911, C1 => n5943, C2 => 
                           n7040, A => n6226, ZN => n6223);
   U1184 : OAI22_X1 port map( A1 => n4660, A2 => n5945, B1 => n4402, B2 => 
                           n5946, ZN => n6226);
   U1185 : AOI221_X1 port map( B1 => n5947, B2 => n6976, C1 => n5948, C2 => 
                           n6944, A => n6227, ZN => n6222);
   U1186 : OAI22_X1 port map( A1 => n4596, A2 => n5950, B1 => n4338, B2 => 
                           n5951, ZN => n6227);
   U1187 : AOI221_X1 port map( B1 => n5952, B2 => n6228, C1 => n5190, C2 => 
                           OUT2_16_port, A => n6229, ZN => n6221);
   U1188 : OAI22_X1 port map( A1 => n4628, A2 => n5955, B1 => n4370, B2 => 
                           n5956, ZN => n6229);
   U1189 : NAND4_X1 port map( A1 => n6230, A2 => n6231, A3 => n6232, A4 => 
                           n6233, ZN => n6228);
   U1190 : AOI221_X1 port map( B1 => n5961, B2 => n6879, C1 => n5962, C2 => 
                           n6655, A => n6234, ZN => n6233);
   U1191 : OAI222_X1 port map( A1 => n4724, A2 => n5964, B1 => n4178, B2 => 
                           n5965, C1 => n4434, C2 => n5966, ZN => n6234);
   U1192 : AOI221_X1 port map( B1 => n5967, B2 => n6783, C1 => n5968, C2 => 
                           n6687, A => n6235, ZN => n6232);
   U1193 : OAI22_X1 port map( A1 => n4500, A2 => n5970, B1 => n4242, B2 => 
                           n5971, ZN => n6235);
   U1194 : AOI221_X1 port map( B1 => n5972, B2 => n6719, C1 => n5973, C2 => 
                           n6815, A => n6236, ZN => n6231);
   U1195 : OAI222_X1 port map( A1 => n4692, A2 => n5975, B1 => n4210, B2 => 
                           n5976, C1 => n4466, C2 => n5977, ZN => n6236);
   U1196 : AOI221_X1 port map( B1 => n5978, B2 => n6751, C1 => n5979, C2 => 
                           n6847, A => n6237, ZN => n6230);
   U1197 : OAI22_X1 port map( A1 => n4564, A2 => n5981, B1 => n4306, B2 => 
                           n5982, ZN => n6237);
   U1198 : NAND4_X1 port map( A1 => n6238, A2 => n6239, A3 => n6240, A4 => 
                           n6241, ZN => n4114);
   U1199 : AOI221_X1 port map( B1 => n5937, B2 => n7007, C1 => n5938, C2 => 
                           n7071, A => n6242, ZN => n6241);
   U1200 : OAI22_X1 port map( A1 => n4533, A2 => n5940, B1 => n4275, B2 => 
                           n5941, ZN => n6242);
   U1201 : AOI221_X1 port map( B1 => n5942, B2 => n6912, C1 => n5943, C2 => 
                           n7039, A => n6243, ZN => n6240);
   U1202 : OAI22_X1 port map( A1 => n4661, A2 => n5945, B1 => n4403, B2 => 
                           n5946, ZN => n6243);
   U1203 : AOI221_X1 port map( B1 => n5947, B2 => n6975, C1 => n5948, C2 => 
                           n6943, A => n6244, ZN => n6239);
   U1204 : OAI22_X1 port map( A1 => n4597, A2 => n5950, B1 => n4339, B2 => 
                           n5951, ZN => n6244);
   U1205 : AOI221_X1 port map( B1 => n5952, B2 => n6245, C1 => n5190, C2 => 
                           OUT2_15_port, A => n6246, ZN => n6238);
   U1206 : OAI22_X1 port map( A1 => n4629, A2 => n5955, B1 => n4371, B2 => 
                           n5956, ZN => n6246);
   U1207 : NAND4_X1 port map( A1 => n6247, A2 => n6248, A3 => n6249, A4 => 
                           n6250, ZN => n6245);
   U1208 : AOI221_X1 port map( B1 => n5961, B2 => n6880, C1 => n5962, C2 => 
                           n6656, A => n6251, ZN => n6250);
   U1209 : OAI222_X1 port map( A1 => n4725, A2 => n5964, B1 => n4179, B2 => 
                           n5965, C1 => n4435, C2 => n5966, ZN => n6251);
   U1210 : AOI221_X1 port map( B1 => n5967, B2 => n6784, C1 => n5968, C2 => 
                           n6688, A => n6252, ZN => n6249);
   U1211 : OAI22_X1 port map( A1 => n4501, A2 => n5970, B1 => n4243, B2 => 
                           n5971, ZN => n6252);
   U1212 : AOI221_X1 port map( B1 => n5972, B2 => n6720, C1 => n5973, C2 => 
                           n6816, A => n6253, ZN => n6248);
   U1213 : OAI222_X1 port map( A1 => n4693, A2 => n5975, B1 => n4211, B2 => 
                           n5976, C1 => n4467, C2 => n5977, ZN => n6253);
   U1214 : AOI221_X1 port map( B1 => n5978, B2 => n6752, C1 => n5979, C2 => 
                           n6848, A => n6254, ZN => n6247);
   U1215 : OAI22_X1 port map( A1 => n4565, A2 => n5981, B1 => n4307, B2 => 
                           n5982, ZN => n6254);
   U1216 : NAND4_X1 port map( A1 => n6255, A2 => n6256, A3 => n6257, A4 => 
                           n6258, ZN => n4113);
   U1217 : AOI221_X1 port map( B1 => n5937, B2 => n7006, C1 => n5938, C2 => 
                           n7070, A => n6259, ZN => n6258);
   U1218 : OAI22_X1 port map( A1 => n4534, A2 => n5940, B1 => n4276, B2 => 
                           n5941, ZN => n6259);
   U1219 : AOI221_X1 port map( B1 => n5942, B2 => n6913, C1 => n5943, C2 => 
                           n7038, A => n6260, ZN => n6257);
   U1220 : OAI22_X1 port map( A1 => n4662, A2 => n5945, B1 => n4404, B2 => 
                           n5946, ZN => n6260);
   U1221 : AOI221_X1 port map( B1 => n5947, B2 => n6974, C1 => n5948, C2 => 
                           n6942, A => n6261, ZN => n6256);
   U1222 : OAI22_X1 port map( A1 => n4598, A2 => n5950, B1 => n4340, B2 => 
                           n5951, ZN => n6261);
   U1223 : AOI221_X1 port map( B1 => n5952, B2 => n6262, C1 => n5190, C2 => 
                           OUT2_14_port, A => n6263, ZN => n6255);
   U1224 : OAI22_X1 port map( A1 => n4630, A2 => n5955, B1 => n4372, B2 => 
                           n5956, ZN => n6263);
   U1225 : NAND4_X1 port map( A1 => n6264, A2 => n6265, A3 => n6266, A4 => 
                           n6267, ZN => n6262);
   U1226 : AOI221_X1 port map( B1 => n5961, B2 => n6881, C1 => n5962, C2 => 
                           n6657, A => n6268, ZN => n6267);
   U1227 : OAI222_X1 port map( A1 => n4726, A2 => n5964, B1 => n4180, B2 => 
                           n5965, C1 => n4436, C2 => n5966, ZN => n6268);
   U1228 : AOI221_X1 port map( B1 => n5967, B2 => n6785, C1 => n5968, C2 => 
                           n6689, A => n6269, ZN => n6266);
   U1229 : OAI22_X1 port map( A1 => n4502, A2 => n5970, B1 => n4244, B2 => 
                           n5971, ZN => n6269);
   U1230 : AOI221_X1 port map( B1 => n5972, B2 => n6721, C1 => n5973, C2 => 
                           n6817, A => n6270, ZN => n6265);
   U1231 : OAI222_X1 port map( A1 => n4694, A2 => n5975, B1 => n4212, B2 => 
                           n5976, C1 => n4468, C2 => n5977, ZN => n6270);
   U1232 : AOI221_X1 port map( B1 => n5978, B2 => n6753, C1 => n5979, C2 => 
                           n6849, A => n6271, ZN => n6264);
   U1233 : OAI22_X1 port map( A1 => n4566, A2 => n5981, B1 => n4308, B2 => 
                           n5982, ZN => n6271);
   U1234 : NAND4_X1 port map( A1 => n6272, A2 => n6273, A3 => n6274, A4 => 
                           n6275, ZN => n4112);
   U1235 : AOI221_X1 port map( B1 => n5937, B2 => n7005, C1 => n5938, C2 => 
                           n7069, A => n6276, ZN => n6275);
   U1236 : OAI22_X1 port map( A1 => n4535, A2 => n5940, B1 => n4277, B2 => 
                           n5941, ZN => n6276);
   U1237 : AOI221_X1 port map( B1 => n5942, B2 => n6914, C1 => n5943, C2 => 
                           n7037, A => n6277, ZN => n6274);
   U1238 : OAI22_X1 port map( A1 => n4663, A2 => n5945, B1 => n4405, B2 => 
                           n5946, ZN => n6277);
   U1239 : AOI221_X1 port map( B1 => n5947, B2 => n6973, C1 => n5948, C2 => 
                           n6941, A => n6278, ZN => n6273);
   U1240 : OAI22_X1 port map( A1 => n4599, A2 => n5950, B1 => n4341, B2 => 
                           n5951, ZN => n6278);
   U1241 : AOI221_X1 port map( B1 => n5952, B2 => n6279, C1 => n5190, C2 => 
                           OUT2_13_port, A => n6280, ZN => n6272);
   U1242 : OAI22_X1 port map( A1 => n4631, A2 => n5955, B1 => n4373, B2 => 
                           n5956, ZN => n6280);
   U1243 : NAND4_X1 port map( A1 => n6281, A2 => n6282, A3 => n6283, A4 => 
                           n6284, ZN => n6279);
   U1244 : AOI221_X1 port map( B1 => n5961, B2 => n6882, C1 => n5962, C2 => 
                           n6658, A => n6285, ZN => n6284);
   U1245 : OAI222_X1 port map( A1 => n4727, A2 => n5964, B1 => n4181, B2 => 
                           n5965, C1 => n4437, C2 => n5966, ZN => n6285);
   U1246 : AOI221_X1 port map( B1 => n5967, B2 => n6786, C1 => n5968, C2 => 
                           n6690, A => n6286, ZN => n6283);
   U1247 : OAI22_X1 port map( A1 => n4503, A2 => n5970, B1 => n4245, B2 => 
                           n5971, ZN => n6286);
   U1248 : AOI221_X1 port map( B1 => n5972, B2 => n6722, C1 => n5973, C2 => 
                           n6818, A => n6287, ZN => n6282);
   U1249 : OAI222_X1 port map( A1 => n4695, A2 => n5975, B1 => n4213, B2 => 
                           n5976, C1 => n4469, C2 => n5977, ZN => n6287);
   U1250 : AOI221_X1 port map( B1 => n5978, B2 => n6754, C1 => n5979, C2 => 
                           n6850, A => n6288, ZN => n6281);
   U1251 : OAI22_X1 port map( A1 => n4567, A2 => n5981, B1 => n4309, B2 => 
                           n5982, ZN => n6288);
   U1252 : NAND4_X1 port map( A1 => n6289, A2 => n6290, A3 => n6291, A4 => 
                           n6292, ZN => n4111);
   U1253 : AOI221_X1 port map( B1 => n5937, B2 => n7004, C1 => n5938, C2 => 
                           n7068, A => n6293, ZN => n6292);
   U1254 : OAI22_X1 port map( A1 => n4536, A2 => n5940, B1 => n4278, B2 => 
                           n5941, ZN => n6293);
   U1255 : AOI221_X1 port map( B1 => n5942, B2 => n6915, C1 => n5943, C2 => 
                           n7036, A => n6294, ZN => n6291);
   U1256 : OAI22_X1 port map( A1 => n4664, A2 => n5945, B1 => n4406, B2 => 
                           n5946, ZN => n6294);
   U1257 : AOI221_X1 port map( B1 => n5947, B2 => n6972, C1 => n5948, C2 => 
                           n6940, A => n6295, ZN => n6290);
   U1258 : OAI22_X1 port map( A1 => n4600, A2 => n5950, B1 => n4342, B2 => 
                           n5951, ZN => n6295);
   U1259 : AOI221_X1 port map( B1 => n5952, B2 => n6296, C1 => n5190, C2 => 
                           OUT2_12_port, A => n6297, ZN => n6289);
   U1260 : OAI22_X1 port map( A1 => n4632, A2 => n5955, B1 => n4374, B2 => 
                           n5956, ZN => n6297);
   U1261 : NAND4_X1 port map( A1 => n6298, A2 => n6299, A3 => n6300, A4 => 
                           n6301, ZN => n6296);
   U1262 : AOI221_X1 port map( B1 => n5961, B2 => n6883, C1 => n5962, C2 => 
                           n6659, A => n6302, ZN => n6301);
   U1263 : OAI222_X1 port map( A1 => n4728, A2 => n5964, B1 => n4182, B2 => 
                           n5965, C1 => n4438, C2 => n5966, ZN => n6302);
   U1264 : AOI221_X1 port map( B1 => n5967, B2 => n6787, C1 => n5968, C2 => 
                           n6691, A => n6303, ZN => n6300);
   U1265 : OAI22_X1 port map( A1 => n4504, A2 => n5970, B1 => n4246, B2 => 
                           n5971, ZN => n6303);
   U1266 : AOI221_X1 port map( B1 => n5972, B2 => n6723, C1 => n5973, C2 => 
                           n6819, A => n6304, ZN => n6299);
   U1267 : OAI222_X1 port map( A1 => n4696, A2 => n5975, B1 => n4214, B2 => 
                           n5976, C1 => n4470, C2 => n5977, ZN => n6304);
   U1268 : AOI221_X1 port map( B1 => n5978, B2 => n6755, C1 => n5979, C2 => 
                           n6851, A => n6305, ZN => n6298);
   U1269 : OAI22_X1 port map( A1 => n4568, A2 => n5981, B1 => n4310, B2 => 
                           n5982, ZN => n6305);
   U1270 : NAND4_X1 port map( A1 => n6306, A2 => n6307, A3 => n6308, A4 => 
                           n6309, ZN => n4110);
   U1271 : AOI221_X1 port map( B1 => n5937, B2 => n7003, C1 => n5938, C2 => 
                           n7067, A => n6310, ZN => n6309);
   U1272 : OAI22_X1 port map( A1 => n4537, A2 => n5940, B1 => n4279, B2 => 
                           n5941, ZN => n6310);
   U1273 : AOI221_X1 port map( B1 => n5942, B2 => n6916, C1 => n5943, C2 => 
                           n7035, A => n6311, ZN => n6308);
   U1274 : OAI22_X1 port map( A1 => n4665, A2 => n5945, B1 => n4407, B2 => 
                           n5946, ZN => n6311);
   U1275 : AOI221_X1 port map( B1 => n5947, B2 => n6971, C1 => n5948, C2 => 
                           n6939, A => n6312, ZN => n6307);
   U1276 : OAI22_X1 port map( A1 => n4601, A2 => n5950, B1 => n4343, B2 => 
                           n5951, ZN => n6312);
   U1277 : AOI221_X1 port map( B1 => n5952, B2 => n6313, C1 => n5190, C2 => 
                           OUT2_11_port, A => n6314, ZN => n6306);
   U1278 : OAI22_X1 port map( A1 => n4633, A2 => n5955, B1 => n4375, B2 => 
                           n5956, ZN => n6314);
   U1279 : NAND4_X1 port map( A1 => n6315, A2 => n6316, A3 => n6317, A4 => 
                           n6318, ZN => n6313);
   U1280 : AOI221_X1 port map( B1 => n5961, B2 => n6884, C1 => n5962, C2 => 
                           n6660, A => n6319, ZN => n6318);
   U1281 : OAI222_X1 port map( A1 => n4729, A2 => n5964, B1 => n4183, B2 => 
                           n5965, C1 => n4439, C2 => n5966, ZN => n6319);
   U1282 : AOI221_X1 port map( B1 => n5967, B2 => n6788, C1 => n5968, C2 => 
                           n6692, A => n6320, ZN => n6317);
   U1283 : OAI22_X1 port map( A1 => n4505, A2 => n5970, B1 => n4247, B2 => 
                           n5971, ZN => n6320);
   U1284 : AOI221_X1 port map( B1 => n5972, B2 => n6724, C1 => n5973, C2 => 
                           n6820, A => n6321, ZN => n6316);
   U1285 : OAI222_X1 port map( A1 => n4697, A2 => n5975, B1 => n4215, B2 => 
                           n5976, C1 => n4471, C2 => n5977, ZN => n6321);
   U1286 : AOI221_X1 port map( B1 => n5978, B2 => n6756, C1 => n5979, C2 => 
                           n6852, A => n6322, ZN => n6315);
   U1287 : OAI22_X1 port map( A1 => n4569, A2 => n5981, B1 => n4311, B2 => 
                           n5982, ZN => n6322);
   U1288 : NAND4_X1 port map( A1 => n6323, A2 => n6324, A3 => n6325, A4 => 
                           n6326, ZN => n4109);
   U1289 : AOI221_X1 port map( B1 => n5937, B2 => n7002, C1 => n5938, C2 => 
                           n7066, A => n6327, ZN => n6326);
   U1290 : OAI22_X1 port map( A1 => n4538, A2 => n5940, B1 => n4280, B2 => 
                           n5941, ZN => n6327);
   U1291 : AOI221_X1 port map( B1 => n5942, B2 => n6917, C1 => n5943, C2 => 
                           n7034, A => n6328, ZN => n6325);
   U1292 : OAI22_X1 port map( A1 => n4666, A2 => n5945, B1 => n4408, B2 => 
                           n5946, ZN => n6328);
   U1293 : AOI221_X1 port map( B1 => n5947, B2 => n6970, C1 => n5948, C2 => 
                           n6938, A => n6329, ZN => n6324);
   U1294 : OAI22_X1 port map( A1 => n4602, A2 => n5950, B1 => n4344, B2 => 
                           n5951, ZN => n6329);
   U1295 : AOI221_X1 port map( B1 => n5952, B2 => n6330, C1 => n5190, C2 => 
                           OUT2_10_port, A => n6331, ZN => n6323);
   U1296 : OAI22_X1 port map( A1 => n4634, A2 => n5955, B1 => n4376, B2 => 
                           n5956, ZN => n6331);
   U1297 : NAND4_X1 port map( A1 => n6332, A2 => n6333, A3 => n6334, A4 => 
                           n6335, ZN => n6330);
   U1298 : AOI221_X1 port map( B1 => n5961, B2 => n6885, C1 => n5962, C2 => 
                           n6661, A => n6336, ZN => n6335);
   U1299 : OAI222_X1 port map( A1 => n4730, A2 => n5964, B1 => n4184, B2 => 
                           n5965, C1 => n4440, C2 => n5966, ZN => n6336);
   U1300 : AOI221_X1 port map( B1 => n5967, B2 => n6789, C1 => n5968, C2 => 
                           n6693, A => n6337, ZN => n6334);
   U1301 : OAI22_X1 port map( A1 => n4506, A2 => n5970, B1 => n4248, B2 => 
                           n5971, ZN => n6337);
   U1302 : AOI221_X1 port map( B1 => n5972, B2 => n6725, C1 => n5973, C2 => 
                           n6821, A => n6338, ZN => n6333);
   U1303 : OAI222_X1 port map( A1 => n4698, A2 => n5975, B1 => n4216, B2 => 
                           n5976, C1 => n4472, C2 => n5977, ZN => n6338);
   U1304 : AOI221_X1 port map( B1 => n5978, B2 => n6757, C1 => n5979, C2 => 
                           n6853, A => n6339, ZN => n6332);
   U1305 : OAI22_X1 port map( A1 => n4570, A2 => n5981, B1 => n4312, B2 => 
                           n5982, ZN => n6339);
   U1306 : NAND4_X1 port map( A1 => n6340, A2 => n6341, A3 => n6342, A4 => 
                           n6343, ZN => n4108);
   U1307 : AOI221_X1 port map( B1 => n5937, B2 => n7001, C1 => n5938, C2 => 
                           n7065, A => n6344, ZN => n6343);
   U1308 : OAI22_X1 port map( A1 => n4539, A2 => n5940, B1 => n4281, B2 => 
                           n5941, ZN => n6344);
   U1309 : AOI221_X1 port map( B1 => n5942, B2 => n6918, C1 => n5943, C2 => 
                           n7033, A => n6345, ZN => n6342);
   U1310 : OAI22_X1 port map( A1 => n4667, A2 => n5945, B1 => n4409, B2 => 
                           n5946, ZN => n6345);
   U1311 : AOI221_X1 port map( B1 => n5947, B2 => n6969, C1 => n5948, C2 => 
                           n6937, A => n6346, ZN => n6341);
   U1312 : OAI22_X1 port map( A1 => n4603, A2 => n5950, B1 => n4345, B2 => 
                           n5951, ZN => n6346);
   U1313 : AOI221_X1 port map( B1 => n5952, B2 => n6347, C1 => n5190, C2 => 
                           OUT2_9_port, A => n6348, ZN => n6340);
   U1314 : OAI22_X1 port map( A1 => n4635, A2 => n5955, B1 => n4377, B2 => 
                           n5956, ZN => n6348);
   U1315 : NAND4_X1 port map( A1 => n6349, A2 => n6350, A3 => n6351, A4 => 
                           n6352, ZN => n6347);
   U1316 : AOI221_X1 port map( B1 => n5961, B2 => n6886, C1 => n5962, C2 => 
                           n6662, A => n6353, ZN => n6352);
   U1317 : OAI222_X1 port map( A1 => n4731, A2 => n5964, B1 => n4185, B2 => 
                           n5965, C1 => n4441, C2 => n5966, ZN => n6353);
   U1318 : AOI221_X1 port map( B1 => n5967, B2 => n6790, C1 => n5968, C2 => 
                           n6694, A => n6354, ZN => n6351);
   U1319 : OAI22_X1 port map( A1 => n4507, A2 => n5970, B1 => n4249, B2 => 
                           n5971, ZN => n6354);
   U1320 : AOI221_X1 port map( B1 => n5972, B2 => n6726, C1 => n5973, C2 => 
                           n6822, A => n6355, ZN => n6350);
   U1321 : OAI222_X1 port map( A1 => n4699, A2 => n5975, B1 => n4217, B2 => 
                           n5976, C1 => n4473, C2 => n5977, ZN => n6355);
   U1322 : AOI221_X1 port map( B1 => n5978, B2 => n6758, C1 => n5979, C2 => 
                           n6854, A => n6356, ZN => n6349);
   U1323 : OAI22_X1 port map( A1 => n4571, A2 => n5981, B1 => n4313, B2 => 
                           n5982, ZN => n6356);
   U1324 : NAND4_X1 port map( A1 => n6357, A2 => n6358, A3 => n6359, A4 => 
                           n6360, ZN => n4107);
   U1325 : AOI221_X1 port map( B1 => n5937, B2 => n7000, C1 => n5938, C2 => 
                           n7064, A => n6361, ZN => n6360);
   U1326 : OAI22_X1 port map( A1 => n4540, A2 => n5940, B1 => n4282, B2 => 
                           n5941, ZN => n6361);
   U1327 : AOI221_X1 port map( B1 => n5942, B2 => n6919, C1 => n5943, C2 => 
                           n7032, A => n6362, ZN => n6359);
   U1328 : OAI22_X1 port map( A1 => n4668, A2 => n5945, B1 => n4410, B2 => 
                           n5946, ZN => n6362);
   U1329 : AOI221_X1 port map( B1 => n5947, B2 => n6968, C1 => n5948, C2 => 
                           n6936, A => n6363, ZN => n6358);
   U1330 : OAI22_X1 port map( A1 => n4604, A2 => n5950, B1 => n4346, B2 => 
                           n5951, ZN => n6363);
   U1331 : AOI221_X1 port map( B1 => n5952, B2 => n6364, C1 => n5190, C2 => 
                           OUT2_8_port, A => n6365, ZN => n6357);
   U1332 : OAI22_X1 port map( A1 => n4636, A2 => n5955, B1 => n4378, B2 => 
                           n5956, ZN => n6365);
   U1333 : NAND4_X1 port map( A1 => n6366, A2 => n6367, A3 => n6368, A4 => 
                           n6369, ZN => n6364);
   U1334 : AOI221_X1 port map( B1 => n5961, B2 => n6887, C1 => n5962, C2 => 
                           n6663, A => n6370, ZN => n6369);
   U1335 : OAI222_X1 port map( A1 => n4732, A2 => n5964, B1 => n4186, B2 => 
                           n5965, C1 => n4442, C2 => n5966, ZN => n6370);
   U1336 : AOI221_X1 port map( B1 => n5967, B2 => n6791, C1 => n5968, C2 => 
                           n6695, A => n6371, ZN => n6368);
   U1337 : OAI22_X1 port map( A1 => n4508, A2 => n5970, B1 => n4250, B2 => 
                           n5971, ZN => n6371);
   U1338 : AOI221_X1 port map( B1 => n5972, B2 => n6727, C1 => n5973, C2 => 
                           n6823, A => n6372, ZN => n6367);
   U1339 : OAI222_X1 port map( A1 => n4700, A2 => n5975, B1 => n4218, B2 => 
                           n5976, C1 => n4474, C2 => n5977, ZN => n6372);
   U1340 : AOI221_X1 port map( B1 => n5978, B2 => n6759, C1 => n5979, C2 => 
                           n6855, A => n6373, ZN => n6366);
   U1341 : OAI22_X1 port map( A1 => n4572, A2 => n5981, B1 => n4314, B2 => 
                           n5982, ZN => n6373);
   U1342 : NAND4_X1 port map( A1 => n6374, A2 => n6375, A3 => n6376, A4 => 
                           n6377, ZN => n4106);
   U1343 : AOI221_X1 port map( B1 => n5937, B2 => n6999, C1 => n5938, C2 => 
                           n7063, A => n6378, ZN => n6377);
   U1344 : OAI22_X1 port map( A1 => n4541, A2 => n5940, B1 => n4283, B2 => 
                           n5941, ZN => n6378);
   U1345 : AOI221_X1 port map( B1 => n5942, B2 => n6920, C1 => n5943, C2 => 
                           n7031, A => n6379, ZN => n6376);
   U1346 : OAI22_X1 port map( A1 => n4669, A2 => n5945, B1 => n4411, B2 => 
                           n5946, ZN => n6379);
   U1347 : AOI221_X1 port map( B1 => n5947, B2 => n6967, C1 => n5948, C2 => 
                           n6935, A => n6380, ZN => n6375);
   U1348 : OAI22_X1 port map( A1 => n4605, A2 => n5950, B1 => n4347, B2 => 
                           n5951, ZN => n6380);
   U1349 : AOI221_X1 port map( B1 => n5952, B2 => n6381, C1 => n5190, C2 => 
                           OUT2_7_port, A => n6382, ZN => n6374);
   U1350 : OAI22_X1 port map( A1 => n4637, A2 => n5955, B1 => n4379, B2 => 
                           n5956, ZN => n6382);
   U1351 : NAND4_X1 port map( A1 => n6383, A2 => n6384, A3 => n6385, A4 => 
                           n6386, ZN => n6381);
   U1352 : AOI221_X1 port map( B1 => n5961, B2 => n6888, C1 => n5962, C2 => 
                           n6664, A => n6387, ZN => n6386);
   U1353 : OAI222_X1 port map( A1 => n4733, A2 => n5964, B1 => n4187, B2 => 
                           n5965, C1 => n4443, C2 => n5966, ZN => n6387);
   U1354 : AOI221_X1 port map( B1 => n5967, B2 => n6792, C1 => n5968, C2 => 
                           n6696, A => n6388, ZN => n6385);
   U1355 : OAI22_X1 port map( A1 => n4509, A2 => n5970, B1 => n4251, B2 => 
                           n5971, ZN => n6388);
   U1356 : AOI221_X1 port map( B1 => n5972, B2 => n6728, C1 => n5973, C2 => 
                           n6824, A => n6389, ZN => n6384);
   U1357 : OAI222_X1 port map( A1 => n4701, A2 => n5975, B1 => n4219, B2 => 
                           n5976, C1 => n4475, C2 => n5977, ZN => n6389);
   U1358 : AOI221_X1 port map( B1 => n5978, B2 => n6760, C1 => n5979, C2 => 
                           n6856, A => n6390, ZN => n6383);
   U1359 : OAI22_X1 port map( A1 => n4573, A2 => n5981, B1 => n4315, B2 => 
                           n5982, ZN => n6390);
   U1360 : NAND4_X1 port map( A1 => n6391, A2 => n6392, A3 => n6393, A4 => 
                           n6394, ZN => n4105);
   U1361 : AOI221_X1 port map( B1 => n5937, B2 => n6998, C1 => n5938, C2 => 
                           n7062, A => n6395, ZN => n6394);
   U1362 : OAI22_X1 port map( A1 => n4542, A2 => n5940, B1 => n4284, B2 => 
                           n5941, ZN => n6395);
   U1363 : AOI221_X1 port map( B1 => n5942, B2 => n6921, C1 => n5943, C2 => 
                           n7030, A => n6396, ZN => n6393);
   U1364 : OAI22_X1 port map( A1 => n4670, A2 => n5945, B1 => n4412, B2 => 
                           n5946, ZN => n6396);
   U1365 : AOI221_X1 port map( B1 => n5947, B2 => n6966, C1 => n5948, C2 => 
                           n6934, A => n6397, ZN => n6392);
   U1366 : OAI22_X1 port map( A1 => n4606, A2 => n5950, B1 => n4348, B2 => 
                           n5951, ZN => n6397);
   U1367 : AOI221_X1 port map( B1 => n5952, B2 => n6398, C1 => n5190, C2 => 
                           OUT2_6_port, A => n6399, ZN => n6391);
   U1368 : OAI22_X1 port map( A1 => n4638, A2 => n5955, B1 => n4380, B2 => 
                           n5956, ZN => n6399);
   U1369 : NAND4_X1 port map( A1 => n6400, A2 => n6401, A3 => n6402, A4 => 
                           n6403, ZN => n6398);
   U1370 : AOI221_X1 port map( B1 => n5961, B2 => n6889, C1 => n5962, C2 => 
                           n6665, A => n6404, ZN => n6403);
   U1371 : OAI222_X1 port map( A1 => n4734, A2 => n5964, B1 => n4188, B2 => 
                           n5965, C1 => n4444, C2 => n5966, ZN => n6404);
   U1372 : AOI221_X1 port map( B1 => n5967, B2 => n6793, C1 => n5968, C2 => 
                           n6697, A => n6405, ZN => n6402);
   U1373 : OAI22_X1 port map( A1 => n4510, A2 => n5970, B1 => n4252, B2 => 
                           n5971, ZN => n6405);
   U1374 : AOI221_X1 port map( B1 => n5972, B2 => n6729, C1 => n5973, C2 => 
                           n6825, A => n6406, ZN => n6401);
   U1375 : OAI222_X1 port map( A1 => n4702, A2 => n5975, B1 => n4220, B2 => 
                           n5976, C1 => n4476, C2 => n5977, ZN => n6406);
   U1376 : AOI221_X1 port map( B1 => n5978, B2 => n6761, C1 => n5979, C2 => 
                           n6857, A => n6407, ZN => n6400);
   U1377 : OAI22_X1 port map( A1 => n4574, A2 => n5981, B1 => n4316, B2 => 
                           n5982, ZN => n6407);
   U1378 : NAND4_X1 port map( A1 => n6408, A2 => n6409, A3 => n6410, A4 => 
                           n6411, ZN => n4104);
   U1379 : AOI221_X1 port map( B1 => n5937, B2 => n6997, C1 => n5938, C2 => 
                           n7061, A => n6412, ZN => n6411);
   U1380 : OAI22_X1 port map( A1 => n4543, A2 => n5940, B1 => n4285, B2 => 
                           n5941, ZN => n6412);
   U1381 : AOI221_X1 port map( B1 => n5942, B2 => n6922, C1 => n5943, C2 => 
                           n7029, A => n6413, ZN => n6410);
   U1382 : OAI22_X1 port map( A1 => n4671, A2 => n5945, B1 => n4413, B2 => 
                           n5946, ZN => n6413);
   U1383 : AOI221_X1 port map( B1 => n5947, B2 => n6965, C1 => n5948, C2 => 
                           n6933, A => n6414, ZN => n6409);
   U1384 : OAI22_X1 port map( A1 => n4607, A2 => n5950, B1 => n4349, B2 => 
                           n5951, ZN => n6414);
   U1385 : AOI221_X1 port map( B1 => n5952, B2 => n6415, C1 => n5190, C2 => 
                           OUT2_5_port, A => n6416, ZN => n6408);
   U1386 : OAI22_X1 port map( A1 => n4639, A2 => n5955, B1 => n4381, B2 => 
                           n5956, ZN => n6416);
   U1387 : NAND4_X1 port map( A1 => n6417, A2 => n6418, A3 => n6419, A4 => 
                           n6420, ZN => n6415);
   U1388 : AOI221_X1 port map( B1 => n5961, B2 => n6890, C1 => n5962, C2 => 
                           n6666, A => n6421, ZN => n6420);
   U1389 : OAI222_X1 port map( A1 => n4735, A2 => n5964, B1 => n4189, B2 => 
                           n5965, C1 => n4445, C2 => n5966, ZN => n6421);
   U1390 : AOI221_X1 port map( B1 => n5967, B2 => n6794, C1 => n5968, C2 => 
                           n6698, A => n6422, ZN => n6419);
   U1391 : OAI22_X1 port map( A1 => n4511, A2 => n5970, B1 => n4253, B2 => 
                           n5971, ZN => n6422);
   U1392 : AOI221_X1 port map( B1 => n5972, B2 => n6730, C1 => n5973, C2 => 
                           n6826, A => n6423, ZN => n6418);
   U1393 : OAI222_X1 port map( A1 => n4703, A2 => n5975, B1 => n4221, B2 => 
                           n5976, C1 => n4477, C2 => n5977, ZN => n6423);
   U1394 : AOI221_X1 port map( B1 => n5978, B2 => n6762, C1 => n5979, C2 => 
                           n6858, A => n6424, ZN => n6417);
   U1395 : OAI22_X1 port map( A1 => n4575, A2 => n5981, B1 => n4317, B2 => 
                           n5982, ZN => n6424);
   U1396 : NAND4_X1 port map( A1 => n6425, A2 => n6426, A3 => n6427, A4 => 
                           n6428, ZN => n4103);
   U1397 : AOI221_X1 port map( B1 => n5937, B2 => n6996, C1 => n5938, C2 => 
                           n7060, A => n6429, ZN => n6428);
   U1398 : OAI22_X1 port map( A1 => n4544, A2 => n5940, B1 => n4286, B2 => 
                           n5941, ZN => n6429);
   U1399 : AOI221_X1 port map( B1 => n5942, B2 => n6923, C1 => n5943, C2 => 
                           n7028, A => n6430, ZN => n6427);
   U1400 : OAI22_X1 port map( A1 => n4672, A2 => n5945, B1 => n4414, B2 => 
                           n5946, ZN => n6430);
   U1401 : AOI221_X1 port map( B1 => n5947, B2 => n6964, C1 => n5948, C2 => 
                           n6932, A => n6431, ZN => n6426);
   U1402 : OAI22_X1 port map( A1 => n4608, A2 => n5950, B1 => n4350, B2 => 
                           n5951, ZN => n6431);
   U1403 : AOI221_X1 port map( B1 => n5952, B2 => n6432, C1 => n5190, C2 => 
                           OUT2_4_port, A => n6433, ZN => n6425);
   U1404 : OAI22_X1 port map( A1 => n4640, A2 => n5955, B1 => n4382, B2 => 
                           n5956, ZN => n6433);
   U1405 : NAND4_X1 port map( A1 => n6434, A2 => n6435, A3 => n6436, A4 => 
                           n6437, ZN => n6432);
   U1406 : AOI221_X1 port map( B1 => n5961, B2 => n6891, C1 => n5962, C2 => 
                           n6667, A => n6438, ZN => n6437);
   U1407 : OAI222_X1 port map( A1 => n4736, A2 => n5964, B1 => n4190, B2 => 
                           n5965, C1 => n4446, C2 => n5966, ZN => n6438);
   U1408 : AOI221_X1 port map( B1 => n5967, B2 => n6795, C1 => n5968, C2 => 
                           n6699, A => n6439, ZN => n6436);
   U1409 : OAI22_X1 port map( A1 => n4512, A2 => n5970, B1 => n4254, B2 => 
                           n5971, ZN => n6439);
   U1410 : AOI221_X1 port map( B1 => n5972, B2 => n6731, C1 => n5973, C2 => 
                           n6827, A => n6440, ZN => n6435);
   U1411 : OAI222_X1 port map( A1 => n4704, A2 => n5975, B1 => n4222, B2 => 
                           n5976, C1 => n4478, C2 => n5977, ZN => n6440);
   U1412 : AOI221_X1 port map( B1 => n5978, B2 => n6763, C1 => n5979, C2 => 
                           n6859, A => n6441, ZN => n6434);
   U1413 : OAI22_X1 port map( A1 => n4576, A2 => n5981, B1 => n4318, B2 => 
                           n5982, ZN => n6441);
   U1414 : NAND4_X1 port map( A1 => n6442, A2 => n6443, A3 => n6444, A4 => 
                           n6445, ZN => n4102);
   U1415 : AOI221_X1 port map( B1 => n5937, B2 => n6995, C1 => n5938, C2 => 
                           n7059, A => n6446, ZN => n6445);
   U1416 : OAI22_X1 port map( A1 => n4545, A2 => n5940, B1 => n4287, B2 => 
                           n5941, ZN => n6446);
   U1417 : AOI221_X1 port map( B1 => n5942, B2 => n6924, C1 => n5943, C2 => 
                           n7027, A => n6447, ZN => n6444);
   U1418 : OAI22_X1 port map( A1 => n4673, A2 => n5945, B1 => n4415, B2 => 
                           n5946, ZN => n6447);
   U1419 : AOI221_X1 port map( B1 => n5947, B2 => n6963, C1 => n5948, C2 => 
                           n6931, A => n6448, ZN => n6443);
   U1420 : OAI22_X1 port map( A1 => n4609, A2 => n5950, B1 => n4351, B2 => 
                           n5951, ZN => n6448);
   U1421 : AOI221_X1 port map( B1 => n5952, B2 => n6449, C1 => n5190, C2 => 
                           OUT2_3_port, A => n6450, ZN => n6442);
   U1422 : OAI22_X1 port map( A1 => n4641, A2 => n5955, B1 => n4383, B2 => 
                           n5956, ZN => n6450);
   U1423 : NAND4_X1 port map( A1 => n6451, A2 => n6452, A3 => n6453, A4 => 
                           n6454, ZN => n6449);
   U1424 : AOI221_X1 port map( B1 => n5961, B2 => n6892, C1 => n5962, C2 => 
                           n6668, A => n6455, ZN => n6454);
   U1425 : OAI222_X1 port map( A1 => n4737, A2 => n5964, B1 => n4191, B2 => 
                           n5965, C1 => n4447, C2 => n5966, ZN => n6455);
   U1426 : AOI221_X1 port map( B1 => n5967, B2 => n6796, C1 => n5968, C2 => 
                           n6700, A => n6456, ZN => n6453);
   U1427 : OAI22_X1 port map( A1 => n4513, A2 => n5970, B1 => n4255, B2 => 
                           n5971, ZN => n6456);
   U1428 : AOI221_X1 port map( B1 => n5972, B2 => n6732, C1 => n5973, C2 => 
                           n6828, A => n6457, ZN => n6452);
   U1429 : OAI222_X1 port map( A1 => n4705, A2 => n5975, B1 => n4223, B2 => 
                           n5976, C1 => n4479, C2 => n5977, ZN => n6457);
   U1430 : AOI221_X1 port map( B1 => n5978, B2 => n6764, C1 => n5979, C2 => 
                           n6860, A => n6458, ZN => n6451);
   U1431 : OAI22_X1 port map( A1 => n4577, A2 => n5981, B1 => n4319, B2 => 
                           n5982, ZN => n6458);
   U1432 : NAND4_X1 port map( A1 => n6459, A2 => n6460, A3 => n6461, A4 => 
                           n6462, ZN => n4101);
   U1433 : AOI221_X1 port map( B1 => n5937, B2 => n6994, C1 => n5938, C2 => 
                           n7058, A => n6463, ZN => n6462);
   U1434 : OAI22_X1 port map( A1 => n4546, A2 => n5940, B1 => n4288, B2 => 
                           n5941, ZN => n6463);
   U1435 : AOI221_X1 port map( B1 => n5942, B2 => n6925, C1 => n5943, C2 => 
                           n7026, A => n6464, ZN => n6461);
   U1436 : OAI22_X1 port map( A1 => n4674, A2 => n5945, B1 => n4416, B2 => 
                           n5946, ZN => n6464);
   U1437 : AOI221_X1 port map( B1 => n5947, B2 => n6962, C1 => n5948, C2 => 
                           n6930, A => n6465, ZN => n6460);
   U1438 : OAI22_X1 port map( A1 => n4610, A2 => n5950, B1 => n4352, B2 => 
                           n5951, ZN => n6465);
   U1439 : AOI221_X1 port map( B1 => n5952, B2 => n6466, C1 => n5190, C2 => 
                           OUT2_2_port, A => n6467, ZN => n6459);
   U1440 : OAI22_X1 port map( A1 => n4642, A2 => n5955, B1 => n4384, B2 => 
                           n5956, ZN => n6467);
   U1441 : NAND4_X1 port map( A1 => n6468, A2 => n6469, A3 => n6470, A4 => 
                           n6471, ZN => n6466);
   U1442 : AOI221_X1 port map( B1 => n5961, B2 => n6893, C1 => n5962, C2 => 
                           n6669, A => n6472, ZN => n6471);
   U1443 : OAI222_X1 port map( A1 => n4738, A2 => n5964, B1 => n4192, B2 => 
                           n5965, C1 => n4448, C2 => n5966, ZN => n6472);
   U1444 : AOI221_X1 port map( B1 => n5967, B2 => n6797, C1 => n5968, C2 => 
                           n6701, A => n6473, ZN => n6470);
   U1445 : OAI22_X1 port map( A1 => n4514, A2 => n5970, B1 => n4256, B2 => 
                           n5971, ZN => n6473);
   U1446 : AOI221_X1 port map( B1 => n5972, B2 => n6733, C1 => n5973, C2 => 
                           n6829, A => n6474, ZN => n6469);
   U1447 : OAI222_X1 port map( A1 => n4706, A2 => n5975, B1 => n4224, B2 => 
                           n5976, C1 => n4480, C2 => n5977, ZN => n6474);
   U1448 : AOI221_X1 port map( B1 => n5978, B2 => n6765, C1 => n5979, C2 => 
                           n6861, A => n6475, ZN => n6468);
   U1449 : OAI22_X1 port map( A1 => n4578, A2 => n5981, B1 => n4320, B2 => 
                           n5982, ZN => n6475);
   U1450 : NAND4_X1 port map( A1 => n6476, A2 => n6477, A3 => n6478, A4 => 
                           n6479, ZN => n4100);
   U1451 : AOI221_X1 port map( B1 => n5937, B2 => n6993, C1 => n5938, C2 => 
                           n7057, A => n6480, ZN => n6479);
   U1452 : OAI22_X1 port map( A1 => n4547, A2 => n5940, B1 => n4289, B2 => 
                           n5941, ZN => n6480);
   U1453 : AOI221_X1 port map( B1 => n5942, B2 => n6926, C1 => n5943, C2 => 
                           n7025, A => n6481, ZN => n6478);
   U1454 : OAI22_X1 port map( A1 => n4675, A2 => n5945, B1 => n4417, B2 => 
                           n5946, ZN => n6481);
   U1455 : AOI221_X1 port map( B1 => n5947, B2 => n6961, C1 => n5948, C2 => 
                           n6929, A => n6482, ZN => n6477);
   U1456 : OAI22_X1 port map( A1 => n4611, A2 => n5950, B1 => n4353, B2 => 
                           n5951, ZN => n6482);
   U1457 : AOI221_X1 port map( B1 => n5952, B2 => n6483, C1 => n5190, C2 => 
                           OUT2_1_port, A => n6484, ZN => n6476);
   U1458 : OAI22_X1 port map( A1 => n4643, A2 => n5955, B1 => n4385, B2 => 
                           n5956, ZN => n6484);
   U1459 : NAND4_X1 port map( A1 => n6485, A2 => n6486, A3 => n6487, A4 => 
                           n6488, ZN => n6483);
   U1460 : AOI221_X1 port map( B1 => n5961, B2 => n6894, C1 => n5962, C2 => 
                           n6670, A => n6489, ZN => n6488);
   U1461 : OAI222_X1 port map( A1 => n4739, A2 => n5964, B1 => n4193, B2 => 
                           n5965, C1 => n4449, C2 => n5966, ZN => n6489);
   U1462 : AOI221_X1 port map( B1 => n5967, B2 => n6798, C1 => n5968, C2 => 
                           n6702, A => n6490, ZN => n6487);
   U1463 : OAI22_X1 port map( A1 => n4515, A2 => n5970, B1 => n4257, B2 => 
                           n5971, ZN => n6490);
   U1464 : AOI221_X1 port map( B1 => n5972, B2 => n6734, C1 => n5973, C2 => 
                           n6830, A => n6491, ZN => n6486);
   U1465 : OAI222_X1 port map( A1 => n4707, A2 => n5975, B1 => n4225, B2 => 
                           n5976, C1 => n4481, C2 => n5977, ZN => n6491);
   U1466 : AOI221_X1 port map( B1 => n5978, B2 => n6766, C1 => n5979, C2 => 
                           n6862, A => n6492, ZN => n6485);
   U1467 : OAI22_X1 port map( A1 => n4579, A2 => n5981, B1 => n4321, B2 => 
                           n5982, ZN => n6492);
   U1468 : NAND4_X1 port map( A1 => n6493, A2 => n6494, A3 => n6495, A4 => 
                           n6496, ZN => n4099);
   U1469 : AOI221_X1 port map( B1 => n5937, B2 => n6992, C1 => n5938, C2 => 
                           n7056, A => n6497, ZN => n6496);
   U1470 : OAI22_X1 port map( A1 => n4548, A2 => n5940, B1 => n4290, B2 => 
                           n5941, ZN => n6497);
   U1471 : AOI221_X1 port map( B1 => n5942, B2 => n6927, C1 => n5943, C2 => 
                           n7024, A => n6503, ZN => n6495);
   U1472 : OAI22_X1 port map( A1 => n4676, A2 => n5945, B1 => n4418, B2 => 
                           n5946, ZN => n6503);
   U1473 : AND2_X1 port map( A1 => n6509, A2 => n5952, ZN => n6499);
   U1474 : AOI221_X1 port map( B1 => n5947, B2 => n6960, C1 => n5948, C2 => 
                           n6928, A => n6510, ZN => n6494);
   U1475 : OAI22_X1 port map( A1 => n4612, A2 => n5950, B1 => n4354, B2 => 
                           n5951, ZN => n6510);
   U1476 : AOI221_X1 port map( B1 => n5952, B2 => n6511, C1 => n5190, C2 => 
                           OUT2_0_port, A => n6512, ZN => n6493);
   U1477 : OAI22_X1 port map( A1 => n4644, A2 => n5955, B1 => n4386, B2 => 
                           n5956, ZN => n6512);
   U1478 : AND3_X1 port map( A1 => n5952, A2 => ADD_RD2(4), A3 => ADD_RD2(3), 
                           ZN => n6505);
   U1479 : NAND4_X1 port map( A1 => n6513, A2 => n6514, A3 => n6515, A4 => 
                           n6516, ZN => n6511);
   U1480 : AOI221_X1 port map( B1 => n5961, B2 => n6895, C1 => n5962, C2 => 
                           n6671, A => n6517, ZN => n6516);
   U1481 : OAI222_X1 port map( A1 => n4740, A2 => n5964, B1 => n4194, B2 => 
                           n5965, C1 => n4450, C2 => n5966, ZN => n6517);
   U1482 : AOI221_X1 port map( B1 => n5967, B2 => n6799, C1 => n5968, C2 => 
                           n6703, A => n6520, ZN => n6515);
   U1483 : OAI22_X1 port map( A1 => n4516, A2 => n5970, B1 => n4258, B2 => 
                           n5971, ZN => n6520);
   U1484 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n6521, 
                           ZN => n6500);
   U1485 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n6501);
   U1486 : AOI221_X1 port map( B1 => n5972, B2 => n6735, C1 => n5973, C2 => 
                           n6831, A => n6522, ZN => n6514);
   U1487 : OAI222_X1 port map( A1 => n4708, A2 => n5975, B1 => n4226, B2 => 
                           n5976, C1 => n4482, C2 => n5977, ZN => n6522);
   U1488 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n6523, 
                           ZN => n6507);
   U1489 : NOR3_X1 port map( A1 => n6523, A2 => ADD_RD2(0), A3 => n6524, ZN => 
                           n6502);
   U1490 : NOR3_X1 port map( A1 => n6523, A2 => ADD_RD2(2), A3 => n6521, ZN => 
                           n6508);
   U1491 : AOI221_X1 port map( B1 => n5978, B2 => n6767, C1 => n5979, C2 => 
                           n6863, A => n6525, ZN => n6513);
   U1492 : OAI22_X1 port map( A1 => n4580, A2 => n5981, B1 => n4322, B2 => 
                           n5982, ZN => n6525);
   U1493 : NOR3_X1 port map( A1 => n6524, A2 => ADD_RD2(1), A3 => n6521, ZN => 
                           n6504);
   U1494 : AND2_X1 port map( A1 => ADD_RD2(4), A2 => n6526, ZN => n6509);
   U1495 : NOR3_X1 port map( A1 => n6524, A2 => n6523, A3 => n6521, ZN => n6506
                           );
   U1496 : INV_X1 port map( A => ADD_RD2(0), ZN => n6521);
   U1497 : INV_X1 port map( A => ADD_RD2(1), ZN => n6523);
   U1498 : NOR2_X1 port map( A1 => n6526, A2 => ADD_RD2(4), ZN => n6519);
   U1499 : INV_X1 port map( A => ADD_RD2(3), ZN => n6526);
   U1500 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n6524, 
                           ZN => n6498);
   U1501 : INV_X1 port map( A => ADD_RD2(2), ZN => n6524);
   U1502 : NOR2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n6518);
   U1503 : OAI22_X1 port map( A1 => n6527, A2 => n6528, B1 => n4485, B2 => 
                           n6529, ZN => n2326);
   U1504 : OAI22_X1 port map( A1 => n6527, A2 => n6530, B1 => n4486, B2 => 
                           n6529, ZN => n2325);
   U1505 : OAI22_X1 port map( A1 => n6527, A2 => n6531, B1 => n4487, B2 => 
                           n6529, ZN => n2324);
   U1506 : OAI22_X1 port map( A1 => n6527, A2 => n6532, B1 => n4488, B2 => 
                           n6529, ZN => n2323);
   U1507 : OAI22_X1 port map( A1 => n6527, A2 => n6533, B1 => n4489, B2 => 
                           n6529, ZN => n2322);
   U1508 : OAI22_X1 port map( A1 => n6527, A2 => n6534, B1 => n4490, B2 => 
                           n6529, ZN => n2321);
   U1509 : OAI22_X1 port map( A1 => n6527, A2 => n6535, B1 => n4491, B2 => 
                           n6529, ZN => n2320);
   U1510 : OAI22_X1 port map( A1 => n6527, A2 => n6536, B1 => n4492, B2 => 
                           n6529, ZN => n2319);
   U1511 : OAI22_X1 port map( A1 => n6527, A2 => n6537, B1 => n4493, B2 => 
                           n6529, ZN => n2318);
   U1512 : OAI22_X1 port map( A1 => n6527, A2 => n6538, B1 => n4494, B2 => 
                           n6529, ZN => n2317);
   U1513 : OAI22_X1 port map( A1 => n6527, A2 => n6539, B1 => n4495, B2 => 
                           n6529, ZN => n2316);
   U1514 : OAI22_X1 port map( A1 => n6527, A2 => n6540, B1 => n4496, B2 => 
                           n6529, ZN => n2315);
   U1515 : OAI22_X1 port map( A1 => n6527, A2 => n6541, B1 => n4497, B2 => 
                           n6529, ZN => n2314);
   U1516 : OAI22_X1 port map( A1 => n6527, A2 => n6542, B1 => n4498, B2 => 
                           n6529, ZN => n2313);
   U1517 : OAI22_X1 port map( A1 => n6527, A2 => n6543, B1 => n4499, B2 => 
                           n6529, ZN => n2312);
   U1518 : OAI22_X1 port map( A1 => n6527, A2 => n6544, B1 => n4500, B2 => 
                           n6529, ZN => n2311);
   U1519 : OAI22_X1 port map( A1 => n6527, A2 => n6545, B1 => n4501, B2 => 
                           n6529, ZN => n2310);
   U1520 : OAI22_X1 port map( A1 => n6527, A2 => n6546, B1 => n4502, B2 => 
                           n6529, ZN => n2309);
   U1521 : OAI22_X1 port map( A1 => n6527, A2 => n6547, B1 => n4503, B2 => 
                           n6529, ZN => n2308);
   U1522 : OAI22_X1 port map( A1 => n6527, A2 => n6548, B1 => n4504, B2 => 
                           n6529, ZN => n2307);
   U1523 : OAI22_X1 port map( A1 => n6527, A2 => n6549, B1 => n4505, B2 => 
                           n6529, ZN => n2306);
   U1524 : OAI22_X1 port map( A1 => n6527, A2 => n6550, B1 => n4506, B2 => 
                           n6529, ZN => n2305);
   U1525 : OAI22_X1 port map( A1 => n6527, A2 => n6551, B1 => n4507, B2 => 
                           n6529, ZN => n2304);
   U1526 : OAI22_X1 port map( A1 => n6527, A2 => n6552, B1 => n4508, B2 => 
                           n6529, ZN => n2303);
   U1527 : OAI22_X1 port map( A1 => n6527, A2 => n6553, B1 => n4509, B2 => 
                           n6529, ZN => n2302);
   U1528 : OAI22_X1 port map( A1 => n6527, A2 => n6554, B1 => n4510, B2 => 
                           n6529, ZN => n2301);
   U1529 : OAI22_X1 port map( A1 => n6527, A2 => n6555, B1 => n4511, B2 => 
                           n6529, ZN => n2300);
   U1530 : OAI22_X1 port map( A1 => n6527, A2 => n6556, B1 => n4512, B2 => 
                           n6529, ZN => n2299);
   U1531 : OAI22_X1 port map( A1 => n6527, A2 => n6557, B1 => n4513, B2 => 
                           n6529, ZN => n2298);
   U1532 : OAI22_X1 port map( A1 => n6527, A2 => n6558, B1 => n4514, B2 => 
                           n6529, ZN => n2297);
   U1533 : OAI22_X1 port map( A1 => n6527, A2 => n6559, B1 => n4515, B2 => 
                           n6529, ZN => n2296);
   U1534 : OAI22_X1 port map( A1 => n6527, A2 => n6560, B1 => n4516, B2 => 
                           n6529, ZN => n2295);
   U1535 : OAI22_X1 port map( A1 => n6528, A2 => n6563, B1 => n4965, B2 => 
                           n6564, ZN => n2294);
   U1536 : OAI22_X1 port map( A1 => n6530, A2 => n6563, B1 => n4966, B2 => 
                           n6564, ZN => n2293);
   U1537 : OAI22_X1 port map( A1 => n6531, A2 => n6563, B1 => n4967, B2 => 
                           n6564, ZN => n2292);
   U1538 : OAI22_X1 port map( A1 => n6532, A2 => n6563, B1 => n4968, B2 => 
                           n6564, ZN => n2291);
   U1539 : OAI22_X1 port map( A1 => n6533, A2 => n6563, B1 => n4969, B2 => 
                           n6564, ZN => n2290);
   U1540 : OAI22_X1 port map( A1 => n6534, A2 => n6563, B1 => n4970, B2 => 
                           n6564, ZN => n2289);
   U1541 : OAI22_X1 port map( A1 => n6535, A2 => n6563, B1 => n4971, B2 => 
                           n6564, ZN => n2288);
   U1542 : OAI22_X1 port map( A1 => n6536, A2 => n6563, B1 => n4972, B2 => 
                           n6564, ZN => n2287);
   U1543 : OAI22_X1 port map( A1 => n6537, A2 => n6563, B1 => n4973, B2 => 
                           n6564, ZN => n2286);
   U1544 : OAI22_X1 port map( A1 => n6538, A2 => n6563, B1 => n4974, B2 => 
                           n6564, ZN => n2285);
   U1545 : OAI22_X1 port map( A1 => n6539, A2 => n6563, B1 => n4975, B2 => 
                           n6564, ZN => n2284);
   U1546 : OAI22_X1 port map( A1 => n6540, A2 => n6563, B1 => n4976, B2 => 
                           n6564, ZN => n2283);
   U1547 : OAI22_X1 port map( A1 => n6541, A2 => n6563, B1 => n4977, B2 => 
                           n6564, ZN => n2282);
   U1548 : OAI22_X1 port map( A1 => n6542, A2 => n6563, B1 => n4978, B2 => 
                           n6564, ZN => n2281);
   U1549 : OAI22_X1 port map( A1 => n6543, A2 => n6563, B1 => n4979, B2 => 
                           n6564, ZN => n2280);
   U1550 : OAI22_X1 port map( A1 => n6544, A2 => n6563, B1 => n4980, B2 => 
                           n6564, ZN => n2279);
   U1551 : OAI22_X1 port map( A1 => n6545, A2 => n6563, B1 => n4981, B2 => 
                           n6564, ZN => n2278);
   U1552 : OAI22_X1 port map( A1 => n6546, A2 => n6563, B1 => n4982, B2 => 
                           n6564, ZN => n2277);
   U1553 : OAI22_X1 port map( A1 => n6547, A2 => n6563, B1 => n4983, B2 => 
                           n6564, ZN => n2276);
   U1554 : OAI22_X1 port map( A1 => n6548, A2 => n6563, B1 => n4984, B2 => 
                           n6564, ZN => n2275);
   U1555 : OAI22_X1 port map( A1 => n6549, A2 => n6563, B1 => n4985, B2 => 
                           n6564, ZN => n2274);
   U1556 : OAI22_X1 port map( A1 => n6550, A2 => n6563, B1 => n4986, B2 => 
                           n6564, ZN => n2273);
   U1557 : OAI22_X1 port map( A1 => n6551, A2 => n6563, B1 => n4987, B2 => 
                           n6564, ZN => n2272);
   U1558 : OAI22_X1 port map( A1 => n6552, A2 => n6563, B1 => n4988, B2 => 
                           n6564, ZN => n2271);
   U1559 : OAI22_X1 port map( A1 => n6553, A2 => n6563, B1 => n4989, B2 => 
                           n6564, ZN => n2270);
   U1560 : OAI22_X1 port map( A1 => n6554, A2 => n6563, B1 => n4990, B2 => 
                           n6564, ZN => n2269);
   U1561 : OAI22_X1 port map( A1 => n6555, A2 => n6563, B1 => n4991, B2 => 
                           n6564, ZN => n2268);
   U1562 : OAI22_X1 port map( A1 => n6556, A2 => n6563, B1 => n4992, B2 => 
                           n6564, ZN => n2267);
   U1563 : OAI22_X1 port map( A1 => n6557, A2 => n6563, B1 => n4993, B2 => 
                           n6564, ZN => n2266);
   U1564 : OAI22_X1 port map( A1 => n6558, A2 => n6563, B1 => n4994, B2 => 
                           n6564, ZN => n2265);
   U1565 : OAI22_X1 port map( A1 => n6559, A2 => n6563, B1 => n4995, B2 => 
                           n6564, ZN => n2264);
   U1566 : OAI22_X1 port map( A1 => n6560, A2 => n6563, B1 => n4996, B2 => 
                           n6564, ZN => n2263);
   U1567 : OAI22_X1 port map( A1 => n6528, A2 => n6566, B1 => n4997, B2 => 
                           n6567, ZN => n2262);
   U1568 : OAI22_X1 port map( A1 => n6530, A2 => n6566, B1 => n4998, B2 => 
                           n6567, ZN => n2261);
   U1569 : OAI22_X1 port map( A1 => n6531, A2 => n6566, B1 => n4999, B2 => 
                           n6567, ZN => n2260);
   U1570 : OAI22_X1 port map( A1 => n6532, A2 => n6566, B1 => n5000, B2 => 
                           n6567, ZN => n2259);
   U1571 : OAI22_X1 port map( A1 => n6533, A2 => n6566, B1 => n5001, B2 => 
                           n6567, ZN => n2258);
   U1572 : OAI22_X1 port map( A1 => n6534, A2 => n6566, B1 => n5002, B2 => 
                           n6567, ZN => n2257);
   U1573 : OAI22_X1 port map( A1 => n6535, A2 => n6566, B1 => n5003, B2 => 
                           n6567, ZN => n2256);
   U1574 : OAI22_X1 port map( A1 => n6536, A2 => n6566, B1 => n5004, B2 => 
                           n6567, ZN => n2255);
   U1575 : OAI22_X1 port map( A1 => n6537, A2 => n6566, B1 => n5005, B2 => 
                           n6567, ZN => n2254);
   U1576 : OAI22_X1 port map( A1 => n6538, A2 => n6566, B1 => n5006, B2 => 
                           n6567, ZN => n2253);
   U1577 : OAI22_X1 port map( A1 => n6539, A2 => n6566, B1 => n5007, B2 => 
                           n6567, ZN => n2252);
   U1578 : OAI22_X1 port map( A1 => n6540, A2 => n6566, B1 => n5008, B2 => 
                           n6567, ZN => n2251);
   U1579 : OAI22_X1 port map( A1 => n6541, A2 => n6566, B1 => n5009, B2 => 
                           n6567, ZN => n2250);
   U1580 : OAI22_X1 port map( A1 => n6542, A2 => n6566, B1 => n5010, B2 => 
                           n6567, ZN => n2249);
   U1581 : OAI22_X1 port map( A1 => n6543, A2 => n6566, B1 => n5011, B2 => 
                           n6567, ZN => n2248);
   U1582 : OAI22_X1 port map( A1 => n6544, A2 => n6566, B1 => n5012, B2 => 
                           n6567, ZN => n2247);
   U1583 : OAI22_X1 port map( A1 => n6545, A2 => n6566, B1 => n5013, B2 => 
                           n6567, ZN => n2246);
   U1584 : OAI22_X1 port map( A1 => n6546, A2 => n6566, B1 => n5014, B2 => 
                           n6567, ZN => n2245);
   U1585 : OAI22_X1 port map( A1 => n6547, A2 => n6566, B1 => n5015, B2 => 
                           n6567, ZN => n2244);
   U1586 : OAI22_X1 port map( A1 => n6548, A2 => n6566, B1 => n5016, B2 => 
                           n6567, ZN => n2243);
   U1587 : OAI22_X1 port map( A1 => n6549, A2 => n6566, B1 => n5017, B2 => 
                           n6567, ZN => n2242);
   U1588 : OAI22_X1 port map( A1 => n6550, A2 => n6566, B1 => n5018, B2 => 
                           n6567, ZN => n2241);
   U1589 : OAI22_X1 port map( A1 => n6551, A2 => n6566, B1 => n5019, B2 => 
                           n6567, ZN => n2240);
   U1590 : OAI22_X1 port map( A1 => n6552, A2 => n6566, B1 => n5020, B2 => 
                           n6567, ZN => n2239);
   U1591 : OAI22_X1 port map( A1 => n6553, A2 => n6566, B1 => n5021, B2 => 
                           n6567, ZN => n2238);
   U1592 : OAI22_X1 port map( A1 => n6554, A2 => n6566, B1 => n5022, B2 => 
                           n6567, ZN => n2237);
   U1593 : OAI22_X1 port map( A1 => n6555, A2 => n6566, B1 => n5023, B2 => 
                           n6567, ZN => n2236);
   U1594 : OAI22_X1 port map( A1 => n6556, A2 => n6566, B1 => n5024, B2 => 
                           n6567, ZN => n2235);
   U1595 : OAI22_X1 port map( A1 => n6557, A2 => n6566, B1 => n5025, B2 => 
                           n6567, ZN => n2234);
   U1596 : OAI22_X1 port map( A1 => n6558, A2 => n6566, B1 => n5026, B2 => 
                           n6567, ZN => n2233);
   U1597 : OAI22_X1 port map( A1 => n6559, A2 => n6566, B1 => n5027, B2 => 
                           n6567, ZN => n2232);
   U1598 : OAI22_X1 port map( A1 => n6560, A2 => n6566, B1 => n5028, B2 => 
                           n6567, ZN => n2231);
   U1599 : OAI22_X1 port map( A1 => n6528, A2 => n6569, B1 => n4741, B2 => 
                           n6570, ZN => n2230);
   U1600 : OAI22_X1 port map( A1 => n6530, A2 => n6569, B1 => n4742, B2 => 
                           n6570, ZN => n2229);
   U1601 : OAI22_X1 port map( A1 => n6531, A2 => n6569, B1 => n4743, B2 => 
                           n6570, ZN => n2228);
   U1602 : OAI22_X1 port map( A1 => n6532, A2 => n6569, B1 => n4744, B2 => 
                           n6570, ZN => n2227);
   U1603 : OAI22_X1 port map( A1 => n6533, A2 => n6569, B1 => n4745, B2 => 
                           n6570, ZN => n2226);
   U1604 : OAI22_X1 port map( A1 => n6534, A2 => n6569, B1 => n4746, B2 => 
                           n6570, ZN => n2225);
   U1605 : OAI22_X1 port map( A1 => n6535, A2 => n6569, B1 => n4747, B2 => 
                           n6570, ZN => n2224);
   U1606 : OAI22_X1 port map( A1 => n6536, A2 => n6569, B1 => n4748, B2 => 
                           n6570, ZN => n2223);
   U1607 : OAI22_X1 port map( A1 => n6537, A2 => n6569, B1 => n4749, B2 => 
                           n6570, ZN => n2222);
   U1608 : OAI22_X1 port map( A1 => n6538, A2 => n6569, B1 => n4750, B2 => 
                           n6570, ZN => n2221);
   U1609 : OAI22_X1 port map( A1 => n6539, A2 => n6569, B1 => n4751, B2 => 
                           n6570, ZN => n2220);
   U1610 : OAI22_X1 port map( A1 => n6540, A2 => n6569, B1 => n4752, B2 => 
                           n6570, ZN => n2219);
   U1611 : OAI22_X1 port map( A1 => n6541, A2 => n6569, B1 => n4753, B2 => 
                           n6570, ZN => n2218);
   U1612 : OAI22_X1 port map( A1 => n6542, A2 => n6569, B1 => n4754, B2 => 
                           n6570, ZN => n2217);
   U1613 : OAI22_X1 port map( A1 => n6543, A2 => n6569, B1 => n4755, B2 => 
                           n6570, ZN => n2216);
   U1614 : OAI22_X1 port map( A1 => n6544, A2 => n6569, B1 => n4756, B2 => 
                           n6570, ZN => n2215);
   U1615 : OAI22_X1 port map( A1 => n6545, A2 => n6569, B1 => n4757, B2 => 
                           n6570, ZN => n2214);
   U1616 : OAI22_X1 port map( A1 => n6546, A2 => n6569, B1 => n4758, B2 => 
                           n6570, ZN => n2213);
   U1617 : OAI22_X1 port map( A1 => n6547, A2 => n6569, B1 => n4759, B2 => 
                           n6570, ZN => n2212);
   U1618 : OAI22_X1 port map( A1 => n6548, A2 => n6569, B1 => n4760, B2 => 
                           n6570, ZN => n2211);
   U1619 : OAI22_X1 port map( A1 => n6549, A2 => n6569, B1 => n4761, B2 => 
                           n6570, ZN => n2210);
   U1620 : OAI22_X1 port map( A1 => n6550, A2 => n6569, B1 => n4762, B2 => 
                           n6570, ZN => n2209);
   U1621 : OAI22_X1 port map( A1 => n6551, A2 => n6569, B1 => n4763, B2 => 
                           n6570, ZN => n2208);
   U1622 : OAI22_X1 port map( A1 => n6552, A2 => n6569, B1 => n4764, B2 => 
                           n6570, ZN => n2207);
   U1623 : OAI22_X1 port map( A1 => n6553, A2 => n6569, B1 => n4765, B2 => 
                           n6570, ZN => n2206);
   U1624 : OAI22_X1 port map( A1 => n6554, A2 => n6569, B1 => n4766, B2 => 
                           n6570, ZN => n2205);
   U1625 : OAI22_X1 port map( A1 => n6555, A2 => n6569, B1 => n4767, B2 => 
                           n6570, ZN => n2204);
   U1626 : OAI22_X1 port map( A1 => n6556, A2 => n6569, B1 => n4768, B2 => 
                           n6570, ZN => n2203);
   U1627 : OAI22_X1 port map( A1 => n6557, A2 => n6569, B1 => n4769, B2 => 
                           n6570, ZN => n2202);
   U1628 : OAI22_X1 port map( A1 => n6558, A2 => n6569, B1 => n4770, B2 => 
                           n6570, ZN => n2201);
   U1629 : OAI22_X1 port map( A1 => n6559, A2 => n6569, B1 => n4771, B2 => 
                           n6570, ZN => n2200);
   U1630 : OAI22_X1 port map( A1 => n6560, A2 => n6569, B1 => n4772, B2 => 
                           n6570, ZN => n2199);
   U1631 : OAI22_X1 port map( A1 => n6528, A2 => n6572, B1 => n4773, B2 => 
                           n6573, ZN => n2198);
   U1632 : OAI22_X1 port map( A1 => n6530, A2 => n6572, B1 => n4774, B2 => 
                           n6573, ZN => n2197);
   U1633 : OAI22_X1 port map( A1 => n6531, A2 => n6572, B1 => n4775, B2 => 
                           n6573, ZN => n2196);
   U1634 : OAI22_X1 port map( A1 => n6532, A2 => n6572, B1 => n4776, B2 => 
                           n6573, ZN => n2195);
   U1635 : OAI22_X1 port map( A1 => n6533, A2 => n6572, B1 => n4777, B2 => 
                           n6573, ZN => n2194);
   U1636 : OAI22_X1 port map( A1 => n6534, A2 => n6572, B1 => n4778, B2 => 
                           n6573, ZN => n2193);
   U1637 : OAI22_X1 port map( A1 => n6535, A2 => n6572, B1 => n4779, B2 => 
                           n6573, ZN => n2192);
   U1638 : OAI22_X1 port map( A1 => n6536, A2 => n6572, B1 => n4780, B2 => 
                           n6573, ZN => n2191);
   U1639 : OAI22_X1 port map( A1 => n6537, A2 => n6572, B1 => n4781, B2 => 
                           n6573, ZN => n2190);
   U1640 : OAI22_X1 port map( A1 => n6538, A2 => n6572, B1 => n4782, B2 => 
                           n6573, ZN => n2189);
   U1641 : OAI22_X1 port map( A1 => n6539, A2 => n6572, B1 => n4783, B2 => 
                           n6573, ZN => n2188);
   U1642 : OAI22_X1 port map( A1 => n6540, A2 => n6572, B1 => n4784, B2 => 
                           n6573, ZN => n2187);
   U1643 : OAI22_X1 port map( A1 => n6541, A2 => n6572, B1 => n4785, B2 => 
                           n6573, ZN => n2186);
   U1644 : OAI22_X1 port map( A1 => n6542, A2 => n6572, B1 => n4786, B2 => 
                           n6573, ZN => n2185);
   U1645 : OAI22_X1 port map( A1 => n6543, A2 => n6572, B1 => n4787, B2 => 
                           n6573, ZN => n2184);
   U1646 : OAI22_X1 port map( A1 => n6544, A2 => n6572, B1 => n4788, B2 => 
                           n6573, ZN => n2183);
   U1647 : OAI22_X1 port map( A1 => n6545, A2 => n6572, B1 => n4789, B2 => 
                           n6573, ZN => n2182);
   U1648 : OAI22_X1 port map( A1 => n6546, A2 => n6572, B1 => n4790, B2 => 
                           n6573, ZN => n2181);
   U1649 : OAI22_X1 port map( A1 => n6547, A2 => n6572, B1 => n4791, B2 => 
                           n6573, ZN => n2180);
   U1650 : OAI22_X1 port map( A1 => n6548, A2 => n6572, B1 => n4792, B2 => 
                           n6573, ZN => n2179);
   U1651 : OAI22_X1 port map( A1 => n6549, A2 => n6572, B1 => n4793, B2 => 
                           n6573, ZN => n2178);
   U1652 : OAI22_X1 port map( A1 => n6550, A2 => n6572, B1 => n4794, B2 => 
                           n6573, ZN => n2177);
   U1653 : OAI22_X1 port map( A1 => n6551, A2 => n6572, B1 => n4795, B2 => 
                           n6573, ZN => n2176);
   U1654 : OAI22_X1 port map( A1 => n6552, A2 => n6572, B1 => n4796, B2 => 
                           n6573, ZN => n2175);
   U1655 : OAI22_X1 port map( A1 => n6553, A2 => n6572, B1 => n4797, B2 => 
                           n6573, ZN => n2174);
   U1656 : OAI22_X1 port map( A1 => n6554, A2 => n6572, B1 => n4798, B2 => 
                           n6573, ZN => n2173);
   U1657 : OAI22_X1 port map( A1 => n6555, A2 => n6572, B1 => n4799, B2 => 
                           n6573, ZN => n2172);
   U1658 : OAI22_X1 port map( A1 => n6556, A2 => n6572, B1 => n4800, B2 => 
                           n6573, ZN => n2171);
   U1659 : OAI22_X1 port map( A1 => n6557, A2 => n6572, B1 => n4801, B2 => 
                           n6573, ZN => n2170);
   U1660 : OAI22_X1 port map( A1 => n6558, A2 => n6572, B1 => n4802, B2 => 
                           n6573, ZN => n2169);
   U1661 : OAI22_X1 port map( A1 => n6559, A2 => n6572, B1 => n4803, B2 => 
                           n6573, ZN => n2168);
   U1662 : OAI22_X1 port map( A1 => n6560, A2 => n6572, B1 => n4804, B2 => 
                           n6573, ZN => n2167);
   U1663 : OAI22_X1 port map( A1 => n6528, A2 => n6575, B1 => n4163, B2 => 
                           n6576, ZN => n2166);
   U1664 : OAI22_X1 port map( A1 => n6530, A2 => n6575, B1 => n4164, B2 => 
                           n6576, ZN => n2165);
   U1665 : OAI22_X1 port map( A1 => n6531, A2 => n6575, B1 => n4165, B2 => 
                           n6576, ZN => n2164);
   U1666 : OAI22_X1 port map( A1 => n6532, A2 => n6575, B1 => n4166, B2 => 
                           n6576, ZN => n2163);
   U1667 : OAI22_X1 port map( A1 => n6533, A2 => n6575, B1 => n4167, B2 => 
                           n6576, ZN => n2162);
   U1668 : OAI22_X1 port map( A1 => n6534, A2 => n6575, B1 => n4168, B2 => 
                           n6576, ZN => n2161);
   U1669 : OAI22_X1 port map( A1 => n6535, A2 => n6575, B1 => n4169, B2 => 
                           n6576, ZN => n2160);
   U1670 : OAI22_X1 port map( A1 => n6536, A2 => n6575, B1 => n4170, B2 => 
                           n6576, ZN => n2159);
   U1671 : OAI22_X1 port map( A1 => n6537, A2 => n6575, B1 => n4171, B2 => 
                           n6576, ZN => n2158);
   U1672 : OAI22_X1 port map( A1 => n6538, A2 => n6575, B1 => n4172, B2 => 
                           n6576, ZN => n2157);
   U1673 : OAI22_X1 port map( A1 => n6539, A2 => n6575, B1 => n4173, B2 => 
                           n6576, ZN => n2156);
   U1674 : OAI22_X1 port map( A1 => n6540, A2 => n6575, B1 => n4174, B2 => 
                           n6576, ZN => n2155);
   U1675 : OAI22_X1 port map( A1 => n6541, A2 => n6575, B1 => n4175, B2 => 
                           n6576, ZN => n2154);
   U1676 : OAI22_X1 port map( A1 => n6542, A2 => n6575, B1 => n4176, B2 => 
                           n6576, ZN => n2153);
   U1677 : OAI22_X1 port map( A1 => n6543, A2 => n6575, B1 => n4177, B2 => 
                           n6576, ZN => n2152);
   U1678 : OAI22_X1 port map( A1 => n6544, A2 => n6575, B1 => n4178, B2 => 
                           n6576, ZN => n2151);
   U1679 : OAI22_X1 port map( A1 => n6545, A2 => n6575, B1 => n4179, B2 => 
                           n6576, ZN => n2150);
   U1680 : OAI22_X1 port map( A1 => n6546, A2 => n6575, B1 => n4180, B2 => 
                           n6576, ZN => n2149);
   U1681 : OAI22_X1 port map( A1 => n6547, A2 => n6575, B1 => n4181, B2 => 
                           n6576, ZN => n2148);
   U1682 : OAI22_X1 port map( A1 => n6548, A2 => n6575, B1 => n4182, B2 => 
                           n6576, ZN => n2147);
   U1683 : OAI22_X1 port map( A1 => n6549, A2 => n6575, B1 => n4183, B2 => 
                           n6576, ZN => n2146);
   U1684 : OAI22_X1 port map( A1 => n6550, A2 => n6575, B1 => n4184, B2 => 
                           n6576, ZN => n2145);
   U1685 : OAI22_X1 port map( A1 => n6551, A2 => n6575, B1 => n4185, B2 => 
                           n6576, ZN => n2144);
   U1686 : OAI22_X1 port map( A1 => n6552, A2 => n6575, B1 => n4186, B2 => 
                           n6576, ZN => n2143);
   U1687 : OAI22_X1 port map( A1 => n6553, A2 => n6575, B1 => n4187, B2 => 
                           n6576, ZN => n2142);
   U1688 : OAI22_X1 port map( A1 => n6554, A2 => n6575, B1 => n4188, B2 => 
                           n6576, ZN => n2141);
   U1689 : OAI22_X1 port map( A1 => n6555, A2 => n6575, B1 => n4189, B2 => 
                           n6576, ZN => n2140);
   U1690 : OAI22_X1 port map( A1 => n6556, A2 => n6575, B1 => n4190, B2 => 
                           n6576, ZN => n2139);
   U1691 : OAI22_X1 port map( A1 => n6557, A2 => n6575, B1 => n4191, B2 => 
                           n6576, ZN => n2138);
   U1692 : OAI22_X1 port map( A1 => n6558, A2 => n6575, B1 => n4192, B2 => 
                           n6576, ZN => n2137);
   U1693 : OAI22_X1 port map( A1 => n6559, A2 => n6575, B1 => n4193, B2 => 
                           n6576, ZN => n2136);
   U1694 : OAI22_X1 port map( A1 => n6560, A2 => n6575, B1 => n4194, B2 => 
                           n6576, ZN => n2135);
   U1695 : OAI22_X1 port map( A1 => n6528, A2 => n6578, B1 => n4677, B2 => 
                           n6579, ZN => n2134);
   U1696 : OAI22_X1 port map( A1 => n6530, A2 => n6578, B1 => n4678, B2 => 
                           n6579, ZN => n2133);
   U1697 : OAI22_X1 port map( A1 => n6531, A2 => n6578, B1 => n4679, B2 => 
                           n6579, ZN => n2132);
   U1698 : OAI22_X1 port map( A1 => n6532, A2 => n6578, B1 => n4680, B2 => 
                           n6579, ZN => n2131);
   U1699 : OAI22_X1 port map( A1 => n6533, A2 => n6578, B1 => n4681, B2 => 
                           n6579, ZN => n2130);
   U1700 : OAI22_X1 port map( A1 => n6534, A2 => n6578, B1 => n4682, B2 => 
                           n6579, ZN => n2129);
   U1701 : OAI22_X1 port map( A1 => n6535, A2 => n6578, B1 => n4683, B2 => 
                           n6579, ZN => n2128);
   U1702 : OAI22_X1 port map( A1 => n6536, A2 => n6578, B1 => n4684, B2 => 
                           n6579, ZN => n2127);
   U1703 : OAI22_X1 port map( A1 => n6537, A2 => n6578, B1 => n4685, B2 => 
                           n6579, ZN => n2126);
   U1704 : OAI22_X1 port map( A1 => n6538, A2 => n6578, B1 => n4686, B2 => 
                           n6579, ZN => n2125);
   U1705 : OAI22_X1 port map( A1 => n6539, A2 => n6578, B1 => n4687, B2 => 
                           n6579, ZN => n2124);
   U1706 : OAI22_X1 port map( A1 => n6540, A2 => n6578, B1 => n4688, B2 => 
                           n6579, ZN => n2123);
   U1707 : OAI22_X1 port map( A1 => n6541, A2 => n6578, B1 => n4689, B2 => 
                           n6579, ZN => n2122);
   U1708 : OAI22_X1 port map( A1 => n6542, A2 => n6578, B1 => n4690, B2 => 
                           n6579, ZN => n2121);
   U1709 : OAI22_X1 port map( A1 => n6543, A2 => n6578, B1 => n4691, B2 => 
                           n6579, ZN => n2120);
   U1710 : OAI22_X1 port map( A1 => n6544, A2 => n6578, B1 => n4692, B2 => 
                           n6579, ZN => n2119);
   U1711 : OAI22_X1 port map( A1 => n6545, A2 => n6578, B1 => n4693, B2 => 
                           n6579, ZN => n2118);
   U1712 : OAI22_X1 port map( A1 => n6546, A2 => n6578, B1 => n4694, B2 => 
                           n6579, ZN => n2117);
   U1713 : OAI22_X1 port map( A1 => n6547, A2 => n6578, B1 => n4695, B2 => 
                           n6579, ZN => n2116);
   U1714 : OAI22_X1 port map( A1 => n6548, A2 => n6578, B1 => n4696, B2 => 
                           n6579, ZN => n2115);
   U1715 : OAI22_X1 port map( A1 => n6549, A2 => n6578, B1 => n4697, B2 => 
                           n6579, ZN => n2114);
   U1716 : OAI22_X1 port map( A1 => n6550, A2 => n6578, B1 => n4698, B2 => 
                           n6579, ZN => n2113);
   U1717 : OAI22_X1 port map( A1 => n6551, A2 => n6578, B1 => n4699, B2 => 
                           n6579, ZN => n2112);
   U1718 : OAI22_X1 port map( A1 => n6552, A2 => n6578, B1 => n4700, B2 => 
                           n6579, ZN => n2111);
   U1719 : OAI22_X1 port map( A1 => n6553, A2 => n6578, B1 => n4701, B2 => 
                           n6579, ZN => n2110);
   U1720 : OAI22_X1 port map( A1 => n6554, A2 => n6578, B1 => n4702, B2 => 
                           n6579, ZN => n2109);
   U1721 : OAI22_X1 port map( A1 => n6555, A2 => n6578, B1 => n4703, B2 => 
                           n6579, ZN => n2108);
   U1722 : OAI22_X1 port map( A1 => n6556, A2 => n6578, B1 => n4704, B2 => 
                           n6579, ZN => n2107);
   U1723 : OAI22_X1 port map( A1 => n6557, A2 => n6578, B1 => n4705, B2 => 
                           n6579, ZN => n2106);
   U1724 : OAI22_X1 port map( A1 => n6558, A2 => n6578, B1 => n4706, B2 => 
                           n6579, ZN => n2105);
   U1725 : OAI22_X1 port map( A1 => n6559, A2 => n6578, B1 => n4707, B2 => 
                           n6579, ZN => n2104);
   U1726 : OAI22_X1 port map( A1 => n6560, A2 => n6578, B1 => n4708, B2 => 
                           n6579, ZN => n2103);
   U1727 : OAI22_X1 port map( A1 => n6528, A2 => n6581, B1 => n4419, B2 => 
                           n6582, ZN => n2102);
   U1728 : OAI22_X1 port map( A1 => n6530, A2 => n6581, B1 => n4420, B2 => 
                           n6582, ZN => n2101);
   U1729 : OAI22_X1 port map( A1 => n6531, A2 => n6581, B1 => n4421, B2 => 
                           n6582, ZN => n2100);
   U1730 : OAI22_X1 port map( A1 => n6532, A2 => n6581, B1 => n4422, B2 => 
                           n6582, ZN => n2099);
   U1731 : OAI22_X1 port map( A1 => n6533, A2 => n6581, B1 => n4423, B2 => 
                           n6582, ZN => n2098);
   U1732 : OAI22_X1 port map( A1 => n6534, A2 => n6581, B1 => n4424, B2 => 
                           n6582, ZN => n2097);
   U1733 : OAI22_X1 port map( A1 => n6535, A2 => n6581, B1 => n4425, B2 => 
                           n6582, ZN => n2096);
   U1734 : OAI22_X1 port map( A1 => n6536, A2 => n6581, B1 => n4426, B2 => 
                           n6582, ZN => n2095);
   U1735 : OAI22_X1 port map( A1 => n6537, A2 => n6581, B1 => n4427, B2 => 
                           n6582, ZN => n2094);
   U1736 : OAI22_X1 port map( A1 => n6538, A2 => n6581, B1 => n4428, B2 => 
                           n6582, ZN => n2093);
   U1737 : OAI22_X1 port map( A1 => n6539, A2 => n6581, B1 => n4429, B2 => 
                           n6582, ZN => n2092);
   U1738 : OAI22_X1 port map( A1 => n6540, A2 => n6581, B1 => n4430, B2 => 
                           n6582, ZN => n2091);
   U1739 : OAI22_X1 port map( A1 => n6541, A2 => n6581, B1 => n4431, B2 => 
                           n6582, ZN => n2090);
   U1740 : OAI22_X1 port map( A1 => n6542, A2 => n6581, B1 => n4432, B2 => 
                           n6582, ZN => n2089);
   U1741 : OAI22_X1 port map( A1 => n6543, A2 => n6581, B1 => n4433, B2 => 
                           n6582, ZN => n2088);
   U1742 : OAI22_X1 port map( A1 => n6544, A2 => n6581, B1 => n4434, B2 => 
                           n6582, ZN => n2087);
   U1743 : OAI22_X1 port map( A1 => n6545, A2 => n6581, B1 => n4435, B2 => 
                           n6582, ZN => n2086);
   U1744 : OAI22_X1 port map( A1 => n6546, A2 => n6581, B1 => n4436, B2 => 
                           n6582, ZN => n2085);
   U1745 : OAI22_X1 port map( A1 => n6547, A2 => n6581, B1 => n4437, B2 => 
                           n6582, ZN => n2084);
   U1746 : OAI22_X1 port map( A1 => n6548, A2 => n6581, B1 => n4438, B2 => 
                           n6582, ZN => n2083);
   U1747 : OAI22_X1 port map( A1 => n6549, A2 => n6581, B1 => n4439, B2 => 
                           n6582, ZN => n2082);
   U1748 : OAI22_X1 port map( A1 => n6550, A2 => n6581, B1 => n4440, B2 => 
                           n6582, ZN => n2081);
   U1749 : OAI22_X1 port map( A1 => n6551, A2 => n6581, B1 => n4441, B2 => 
                           n6582, ZN => n2080);
   U1750 : OAI22_X1 port map( A1 => n6552, A2 => n6581, B1 => n4442, B2 => 
                           n6582, ZN => n2079);
   U1751 : OAI22_X1 port map( A1 => n6553, A2 => n6581, B1 => n4443, B2 => 
                           n6582, ZN => n2078);
   U1752 : OAI22_X1 port map( A1 => n6554, A2 => n6581, B1 => n4444, B2 => 
                           n6582, ZN => n2077);
   U1753 : OAI22_X1 port map( A1 => n6555, A2 => n6581, B1 => n4445, B2 => 
                           n6582, ZN => n2076);
   U1754 : OAI22_X1 port map( A1 => n6556, A2 => n6581, B1 => n4446, B2 => 
                           n6582, ZN => n2075);
   U1755 : OAI22_X1 port map( A1 => n6557, A2 => n6581, B1 => n4447, B2 => 
                           n6582, ZN => n2074);
   U1756 : OAI22_X1 port map( A1 => n6558, A2 => n6581, B1 => n4448, B2 => 
                           n6582, ZN => n2073);
   U1757 : OAI22_X1 port map( A1 => n6559, A2 => n6581, B1 => n4449, B2 => 
                           n6582, ZN => n2072);
   U1758 : OAI22_X1 port map( A1 => n6560, A2 => n6581, B1 => n4450, B2 => 
                           n6582, ZN => n2071);
   U1759 : AND3_X1 port map( A1 => n6584, A2 => n6585, A3 => n6586, ZN => n6562
                           );
   U1760 : OAI22_X1 port map( A1 => n6528, A2 => n6587, B1 => n4805, B2 => 
                           n6588, ZN => n2070);
   U1761 : OAI22_X1 port map( A1 => n6530, A2 => n6587, B1 => n4806, B2 => 
                           n6588, ZN => n2069);
   U1762 : OAI22_X1 port map( A1 => n6531, A2 => n6587, B1 => n4807, B2 => 
                           n6588, ZN => n2068);
   U1763 : OAI22_X1 port map( A1 => n6532, A2 => n6587, B1 => n4808, B2 => 
                           n6588, ZN => n2067);
   U1764 : OAI22_X1 port map( A1 => n6533, A2 => n6587, B1 => n4809, B2 => 
                           n6588, ZN => n2066);
   U1765 : OAI22_X1 port map( A1 => n6534, A2 => n6587, B1 => n4810, B2 => 
                           n6588, ZN => n2065);
   U1766 : OAI22_X1 port map( A1 => n6535, A2 => n6587, B1 => n4811, B2 => 
                           n6588, ZN => n2064);
   U1767 : OAI22_X1 port map( A1 => n6536, A2 => n6587, B1 => n4812, B2 => 
                           n6588, ZN => n2063);
   U1768 : OAI22_X1 port map( A1 => n6537, A2 => n6587, B1 => n4813, B2 => 
                           n6588, ZN => n2062);
   U1769 : OAI22_X1 port map( A1 => n6538, A2 => n6587, B1 => n4814, B2 => 
                           n6588, ZN => n2061);
   U1770 : OAI22_X1 port map( A1 => n6539, A2 => n6587, B1 => n4815, B2 => 
                           n6588, ZN => n2060);
   U1771 : OAI22_X1 port map( A1 => n6540, A2 => n6587, B1 => n4816, B2 => 
                           n6588, ZN => n2059);
   U1772 : OAI22_X1 port map( A1 => n6541, A2 => n6587, B1 => n4817, B2 => 
                           n6588, ZN => n2058);
   U1773 : OAI22_X1 port map( A1 => n6542, A2 => n6587, B1 => n4818, B2 => 
                           n6588, ZN => n2057);
   U1774 : OAI22_X1 port map( A1 => n6543, A2 => n6587, B1 => n4819, B2 => 
                           n6588, ZN => n2056);
   U1775 : OAI22_X1 port map( A1 => n6544, A2 => n6587, B1 => n4820, B2 => 
                           n6588, ZN => n2055);
   U1776 : OAI22_X1 port map( A1 => n6545, A2 => n6587, B1 => n4821, B2 => 
                           n6588, ZN => n2054);
   U1777 : OAI22_X1 port map( A1 => n6546, A2 => n6587, B1 => n4822, B2 => 
                           n6588, ZN => n2053);
   U1778 : OAI22_X1 port map( A1 => n6547, A2 => n6587, B1 => n4823, B2 => 
                           n6588, ZN => n2052);
   U1779 : OAI22_X1 port map( A1 => n6548, A2 => n6587, B1 => n4824, B2 => 
                           n6588, ZN => n2051);
   U1780 : OAI22_X1 port map( A1 => n6549, A2 => n6587, B1 => n4825, B2 => 
                           n6588, ZN => n2050);
   U1781 : OAI22_X1 port map( A1 => n6550, A2 => n6587, B1 => n4826, B2 => 
                           n6588, ZN => n2049);
   U1782 : OAI22_X1 port map( A1 => n6551, A2 => n6587, B1 => n4827, B2 => 
                           n6588, ZN => n2048);
   U1783 : OAI22_X1 port map( A1 => n6552, A2 => n6587, B1 => n4828, B2 => 
                           n6588, ZN => n2047);
   U1784 : OAI22_X1 port map( A1 => n6553, A2 => n6587, B1 => n4829, B2 => 
                           n6588, ZN => n2046);
   U1785 : OAI22_X1 port map( A1 => n6554, A2 => n6587, B1 => n4830, B2 => 
                           n6588, ZN => n2045);
   U1786 : OAI22_X1 port map( A1 => n6555, A2 => n6587, B1 => n4831, B2 => 
                           n6588, ZN => n2044);
   U1787 : OAI22_X1 port map( A1 => n6556, A2 => n6587, B1 => n4832, B2 => 
                           n6588, ZN => n2043);
   U1788 : OAI22_X1 port map( A1 => n6557, A2 => n6587, B1 => n4833, B2 => 
                           n6588, ZN => n2042);
   U1789 : OAI22_X1 port map( A1 => n6558, A2 => n6587, B1 => n4834, B2 => 
                           n6588, ZN => n2041);
   U1790 : OAI22_X1 port map( A1 => n6559, A2 => n6587, B1 => n4835, B2 => 
                           n6588, ZN => n2040);
   U1791 : OAI22_X1 port map( A1 => n6560, A2 => n6587, B1 => n4836, B2 => 
                           n6588, ZN => n2039);
   U1792 : OAI22_X1 port map( A1 => n6528, A2 => n6590, B1 => n4227, B2 => 
                           n6591, ZN => n2038);
   U1793 : OAI22_X1 port map( A1 => n6530, A2 => n6590, B1 => n4228, B2 => 
                           n6591, ZN => n2037);
   U1794 : OAI22_X1 port map( A1 => n6531, A2 => n6590, B1 => n4229, B2 => 
                           n6591, ZN => n2036);
   U1795 : OAI22_X1 port map( A1 => n6532, A2 => n6590, B1 => n4230, B2 => 
                           n6591, ZN => n2035);
   U1796 : OAI22_X1 port map( A1 => n6533, A2 => n6590, B1 => n4231, B2 => 
                           n6591, ZN => n2034);
   U1797 : OAI22_X1 port map( A1 => n6534, A2 => n6590, B1 => n4232, B2 => 
                           n6591, ZN => n2033);
   U1798 : OAI22_X1 port map( A1 => n6535, A2 => n6590, B1 => n4233, B2 => 
                           n6591, ZN => n2032);
   U1799 : OAI22_X1 port map( A1 => n6536, A2 => n6590, B1 => n4234, B2 => 
                           n6591, ZN => n2031);
   U1800 : OAI22_X1 port map( A1 => n6537, A2 => n6590, B1 => n4235, B2 => 
                           n6591, ZN => n2030);
   U1801 : OAI22_X1 port map( A1 => n6538, A2 => n6590, B1 => n4236, B2 => 
                           n6591, ZN => n2029);
   U1802 : OAI22_X1 port map( A1 => n6539, A2 => n6590, B1 => n4237, B2 => 
                           n6591, ZN => n2028);
   U1803 : OAI22_X1 port map( A1 => n6540, A2 => n6590, B1 => n4238, B2 => 
                           n6591, ZN => n2027);
   U1804 : OAI22_X1 port map( A1 => n6541, A2 => n6590, B1 => n4239, B2 => 
                           n6591, ZN => n2026);
   U1805 : OAI22_X1 port map( A1 => n6542, A2 => n6590, B1 => n4240, B2 => 
                           n6591, ZN => n2025);
   U1806 : OAI22_X1 port map( A1 => n6543, A2 => n6590, B1 => n4241, B2 => 
                           n6591, ZN => n2024);
   U1807 : OAI22_X1 port map( A1 => n6544, A2 => n6590, B1 => n4242, B2 => 
                           n6591, ZN => n2023);
   U1808 : OAI22_X1 port map( A1 => n6545, A2 => n6590, B1 => n4243, B2 => 
                           n6591, ZN => n2022);
   U1809 : OAI22_X1 port map( A1 => n6546, A2 => n6590, B1 => n4244, B2 => 
                           n6591, ZN => n2021);
   U1810 : OAI22_X1 port map( A1 => n6547, A2 => n6590, B1 => n4245, B2 => 
                           n6591, ZN => n2020);
   U1811 : OAI22_X1 port map( A1 => n6548, A2 => n6590, B1 => n4246, B2 => 
                           n6591, ZN => n2019);
   U1812 : OAI22_X1 port map( A1 => n6549, A2 => n6590, B1 => n4247, B2 => 
                           n6591, ZN => n2018);
   U1813 : OAI22_X1 port map( A1 => n6550, A2 => n6590, B1 => n4248, B2 => 
                           n6591, ZN => n2017);
   U1814 : OAI22_X1 port map( A1 => n6551, A2 => n6590, B1 => n4249, B2 => 
                           n6591, ZN => n2016);
   U1815 : OAI22_X1 port map( A1 => n6552, A2 => n6590, B1 => n4250, B2 => 
                           n6591, ZN => n2015);
   U1816 : OAI22_X1 port map( A1 => n6553, A2 => n6590, B1 => n4251, B2 => 
                           n6591, ZN => n2014);
   U1817 : OAI22_X1 port map( A1 => n6554, A2 => n6590, B1 => n4252, B2 => 
                           n6591, ZN => n2013);
   U1818 : OAI22_X1 port map( A1 => n6555, A2 => n6590, B1 => n4253, B2 => 
                           n6591, ZN => n2012);
   U1819 : OAI22_X1 port map( A1 => n6556, A2 => n6590, B1 => n4254, B2 => 
                           n6591, ZN => n2011);
   U1820 : OAI22_X1 port map( A1 => n6557, A2 => n6590, B1 => n4255, B2 => 
                           n6591, ZN => n2010);
   U1821 : OAI22_X1 port map( A1 => n6558, A2 => n6590, B1 => n4256, B2 => 
                           n6591, ZN => n2009);
   U1822 : OAI22_X1 port map( A1 => n6559, A2 => n6590, B1 => n4257, B2 => 
                           n6591, ZN => n2008);
   U1823 : OAI22_X1 port map( A1 => n6560, A2 => n6590, B1 => n4258, B2 => 
                           n6591, ZN => n2007);
   U1824 : OAI22_X1 port map( A1 => n6528, A2 => n6592, B1 => n4195, B2 => 
                           n6593, ZN => n2006);
   U1825 : OAI22_X1 port map( A1 => n6530, A2 => n6592, B1 => n4196, B2 => 
                           n6593, ZN => n2005);
   U1826 : OAI22_X1 port map( A1 => n6531, A2 => n6592, B1 => n4197, B2 => 
                           n6593, ZN => n2004);
   U1827 : OAI22_X1 port map( A1 => n6532, A2 => n6592, B1 => n4198, B2 => 
                           n6593, ZN => n2003);
   U1828 : OAI22_X1 port map( A1 => n6533, A2 => n6592, B1 => n4199, B2 => 
                           n6593, ZN => n2002);
   U1829 : OAI22_X1 port map( A1 => n6534, A2 => n6592, B1 => n4200, B2 => 
                           n6593, ZN => n2001);
   U1830 : OAI22_X1 port map( A1 => n6535, A2 => n6592, B1 => n4201, B2 => 
                           n6593, ZN => n2000);
   U1831 : OAI22_X1 port map( A1 => n6536, A2 => n6592, B1 => n4202, B2 => 
                           n6593, ZN => n1999);
   U1832 : OAI22_X1 port map( A1 => n6537, A2 => n6592, B1 => n4203, B2 => 
                           n6593, ZN => n1998);
   U1833 : OAI22_X1 port map( A1 => n6538, A2 => n6592, B1 => n4204, B2 => 
                           n6593, ZN => n1997);
   U1834 : OAI22_X1 port map( A1 => n6539, A2 => n6592, B1 => n4205, B2 => 
                           n6593, ZN => n1996);
   U1835 : OAI22_X1 port map( A1 => n6540, A2 => n6592, B1 => n4206, B2 => 
                           n6593, ZN => n1995);
   U1836 : OAI22_X1 port map( A1 => n6541, A2 => n6592, B1 => n4207, B2 => 
                           n6593, ZN => n1994);
   U1837 : OAI22_X1 port map( A1 => n6542, A2 => n6592, B1 => n4208, B2 => 
                           n6593, ZN => n1993);
   U1838 : OAI22_X1 port map( A1 => n6543, A2 => n6592, B1 => n4209, B2 => 
                           n6593, ZN => n1992);
   U1839 : OAI22_X1 port map( A1 => n6544, A2 => n6592, B1 => n4210, B2 => 
                           n6593, ZN => n1991);
   U1840 : OAI22_X1 port map( A1 => n6545, A2 => n6592, B1 => n4211, B2 => 
                           n6593, ZN => n1990);
   U1841 : OAI22_X1 port map( A1 => n6546, A2 => n6592, B1 => n4212, B2 => 
                           n6593, ZN => n1989);
   U1842 : OAI22_X1 port map( A1 => n6547, A2 => n6592, B1 => n4213, B2 => 
                           n6593, ZN => n1988);
   U1843 : OAI22_X1 port map( A1 => n6548, A2 => n6592, B1 => n4214, B2 => 
                           n6593, ZN => n1987);
   U1844 : OAI22_X1 port map( A1 => n6549, A2 => n6592, B1 => n4215, B2 => 
                           n6593, ZN => n1986);
   U1845 : OAI22_X1 port map( A1 => n6550, A2 => n6592, B1 => n4216, B2 => 
                           n6593, ZN => n1985);
   U1846 : OAI22_X1 port map( A1 => n6551, A2 => n6592, B1 => n4217, B2 => 
                           n6593, ZN => n1984);
   U1847 : OAI22_X1 port map( A1 => n6552, A2 => n6592, B1 => n4218, B2 => 
                           n6593, ZN => n1983);
   U1848 : OAI22_X1 port map( A1 => n6553, A2 => n6592, B1 => n4219, B2 => 
                           n6593, ZN => n1982);
   U1849 : OAI22_X1 port map( A1 => n6554, A2 => n6592, B1 => n4220, B2 => 
                           n6593, ZN => n1981);
   U1850 : OAI22_X1 port map( A1 => n6555, A2 => n6592, B1 => n4221, B2 => 
                           n6593, ZN => n1980);
   U1851 : OAI22_X1 port map( A1 => n6556, A2 => n6592, B1 => n4222, B2 => 
                           n6593, ZN => n1979);
   U1852 : OAI22_X1 port map( A1 => n6557, A2 => n6592, B1 => n4223, B2 => 
                           n6593, ZN => n1978);
   U1853 : OAI22_X1 port map( A1 => n6558, A2 => n6592, B1 => n4224, B2 => 
                           n6593, ZN => n1977);
   U1854 : OAI22_X1 port map( A1 => n6559, A2 => n6592, B1 => n4225, B2 => 
                           n6593, ZN => n1976);
   U1855 : OAI22_X1 port map( A1 => n6560, A2 => n6592, B1 => n4226, B2 => 
                           n6593, ZN => n1975);
   U1856 : OAI22_X1 port map( A1 => n6528, A2 => n6594, B1 => n5029, B2 => 
                           n6595, ZN => n1974);
   U1857 : OAI22_X1 port map( A1 => n6530, A2 => n6594, B1 => n5030, B2 => 
                           n6595, ZN => n1973);
   U1858 : OAI22_X1 port map( A1 => n6531, A2 => n6594, B1 => n5031, B2 => 
                           n6595, ZN => n1972);
   U1859 : OAI22_X1 port map( A1 => n6532, A2 => n6594, B1 => n5032, B2 => 
                           n6595, ZN => n1971);
   U1860 : OAI22_X1 port map( A1 => n6533, A2 => n6594, B1 => n5033, B2 => 
                           n6595, ZN => n1970);
   U1861 : OAI22_X1 port map( A1 => n6534, A2 => n6594, B1 => n5034, B2 => 
                           n6595, ZN => n1969);
   U1862 : OAI22_X1 port map( A1 => n6535, A2 => n6594, B1 => n5035, B2 => 
                           n6595, ZN => n1968);
   U1863 : OAI22_X1 port map( A1 => n6536, A2 => n6594, B1 => n5036, B2 => 
                           n6595, ZN => n1967);
   U1864 : OAI22_X1 port map( A1 => n6537, A2 => n6594, B1 => n5037, B2 => 
                           n6595, ZN => n1966);
   U1865 : OAI22_X1 port map( A1 => n6538, A2 => n6594, B1 => n5038, B2 => 
                           n6595, ZN => n1965);
   U1866 : OAI22_X1 port map( A1 => n6539, A2 => n6594, B1 => n5039, B2 => 
                           n6595, ZN => n1964);
   U1867 : OAI22_X1 port map( A1 => n6540, A2 => n6594, B1 => n5040, B2 => 
                           n6595, ZN => n1963);
   U1868 : OAI22_X1 port map( A1 => n6541, A2 => n6594, B1 => n5041, B2 => 
                           n6595, ZN => n1962);
   U1869 : OAI22_X1 port map( A1 => n6542, A2 => n6594, B1 => n5042, B2 => 
                           n6595, ZN => n1961);
   U1870 : OAI22_X1 port map( A1 => n6543, A2 => n6594, B1 => n5043, B2 => 
                           n6595, ZN => n1960);
   U1871 : OAI22_X1 port map( A1 => n6544, A2 => n6594, B1 => n5044, B2 => 
                           n6595, ZN => n1959);
   U1872 : OAI22_X1 port map( A1 => n6545, A2 => n6594, B1 => n5045, B2 => 
                           n6595, ZN => n1958);
   U1873 : OAI22_X1 port map( A1 => n6546, A2 => n6594, B1 => n5046, B2 => 
                           n6595, ZN => n1957);
   U1874 : OAI22_X1 port map( A1 => n6547, A2 => n6594, B1 => n5047, B2 => 
                           n6595, ZN => n1956);
   U1875 : OAI22_X1 port map( A1 => n6548, A2 => n6594, B1 => n5048, B2 => 
                           n6595, ZN => n1955);
   U1876 : OAI22_X1 port map( A1 => n6549, A2 => n6594, B1 => n5049, B2 => 
                           n6595, ZN => n1954);
   U1877 : OAI22_X1 port map( A1 => n6550, A2 => n6594, B1 => n5050, B2 => 
                           n6595, ZN => n1953);
   U1878 : OAI22_X1 port map( A1 => n6551, A2 => n6594, B1 => n5051, B2 => 
                           n6595, ZN => n1952);
   U1879 : OAI22_X1 port map( A1 => n6552, A2 => n6594, B1 => n5052, B2 => 
                           n6595, ZN => n1951);
   U1880 : OAI22_X1 port map( A1 => n6553, A2 => n6594, B1 => n5053, B2 => 
                           n6595, ZN => n1950);
   U1881 : OAI22_X1 port map( A1 => n6554, A2 => n6594, B1 => n5054, B2 => 
                           n6595, ZN => n1949);
   U1882 : OAI22_X1 port map( A1 => n6555, A2 => n6594, B1 => n5055, B2 => 
                           n6595, ZN => n1948);
   U1883 : OAI22_X1 port map( A1 => n6556, A2 => n6594, B1 => n5056, B2 => 
                           n6595, ZN => n1947);
   U1884 : OAI22_X1 port map( A1 => n6557, A2 => n6594, B1 => n5057, B2 => 
                           n6595, ZN => n1946);
   U1885 : OAI22_X1 port map( A1 => n6558, A2 => n6594, B1 => n5058, B2 => 
                           n6595, ZN => n1945);
   U1886 : OAI22_X1 port map( A1 => n6559, A2 => n6594, B1 => n5059, B2 => 
                           n6595, ZN => n1944);
   U1887 : OAI22_X1 port map( A1 => n6560, A2 => n6594, B1 => n5060, B2 => 
                           n6595, ZN => n1943);
   U1888 : OAI22_X1 port map( A1 => n6528, A2 => n6596, B1 => n5061, B2 => 
                           n6597, ZN => n1942);
   U1889 : OAI22_X1 port map( A1 => n6530, A2 => n6596, B1 => n5062, B2 => 
                           n6597, ZN => n1941);
   U1890 : OAI22_X1 port map( A1 => n6531, A2 => n6596, B1 => n5063, B2 => 
                           n6597, ZN => n1940);
   U1891 : OAI22_X1 port map( A1 => n6532, A2 => n6596, B1 => n5064, B2 => 
                           n6597, ZN => n1939);
   U1892 : OAI22_X1 port map( A1 => n6533, A2 => n6596, B1 => n5065, B2 => 
                           n6597, ZN => n1938);
   U1893 : OAI22_X1 port map( A1 => n6534, A2 => n6596, B1 => n5066, B2 => 
                           n6597, ZN => n1937);
   U1894 : OAI22_X1 port map( A1 => n6535, A2 => n6596, B1 => n5067, B2 => 
                           n6597, ZN => n1936);
   U1895 : OAI22_X1 port map( A1 => n6536, A2 => n6596, B1 => n5068, B2 => 
                           n6597, ZN => n1935);
   U1896 : OAI22_X1 port map( A1 => n6537, A2 => n6596, B1 => n5069, B2 => 
                           n6597, ZN => n1934);
   U1897 : OAI22_X1 port map( A1 => n6538, A2 => n6596, B1 => n5070, B2 => 
                           n6597, ZN => n1933);
   U1898 : OAI22_X1 port map( A1 => n6539, A2 => n6596, B1 => n5071, B2 => 
                           n6597, ZN => n1932);
   U1899 : OAI22_X1 port map( A1 => n6540, A2 => n6596, B1 => n5072, B2 => 
                           n6597, ZN => n1931);
   U1900 : OAI22_X1 port map( A1 => n6541, A2 => n6596, B1 => n5073, B2 => 
                           n6597, ZN => n1930);
   U1901 : OAI22_X1 port map( A1 => n6542, A2 => n6596, B1 => n5074, B2 => 
                           n6597, ZN => n1929);
   U1902 : OAI22_X1 port map( A1 => n6543, A2 => n6596, B1 => n5075, B2 => 
                           n6597, ZN => n1928);
   U1903 : OAI22_X1 port map( A1 => n6544, A2 => n6596, B1 => n5076, B2 => 
                           n6597, ZN => n1927);
   U1904 : OAI22_X1 port map( A1 => n6545, A2 => n6596, B1 => n5077, B2 => 
                           n6597, ZN => n1926);
   U1905 : OAI22_X1 port map( A1 => n6546, A2 => n6596, B1 => n5078, B2 => 
                           n6597, ZN => n1925);
   U1906 : OAI22_X1 port map( A1 => n6547, A2 => n6596, B1 => n5079, B2 => 
                           n6597, ZN => n1924);
   U1907 : OAI22_X1 port map( A1 => n6548, A2 => n6596, B1 => n5080, B2 => 
                           n6597, ZN => n1923);
   U1908 : OAI22_X1 port map( A1 => n6549, A2 => n6596, B1 => n5081, B2 => 
                           n6597, ZN => n1922);
   U1909 : OAI22_X1 port map( A1 => n6550, A2 => n6596, B1 => n5082, B2 => 
                           n6597, ZN => n1921);
   U1910 : OAI22_X1 port map( A1 => n6551, A2 => n6596, B1 => n5083, B2 => 
                           n6597, ZN => n1920);
   U1911 : OAI22_X1 port map( A1 => n6552, A2 => n6596, B1 => n5084, B2 => 
                           n6597, ZN => n1919);
   U1912 : OAI22_X1 port map( A1 => n6553, A2 => n6596, B1 => n5085, B2 => 
                           n6597, ZN => n1918);
   U1913 : OAI22_X1 port map( A1 => n6554, A2 => n6596, B1 => n5086, B2 => 
                           n6597, ZN => n1917);
   U1914 : OAI22_X1 port map( A1 => n6555, A2 => n6596, B1 => n5087, B2 => 
                           n6597, ZN => n1916);
   U1915 : OAI22_X1 port map( A1 => n6556, A2 => n6596, B1 => n5088, B2 => 
                           n6597, ZN => n1915);
   U1916 : OAI22_X1 port map( A1 => n6557, A2 => n6596, B1 => n5089, B2 => 
                           n6597, ZN => n1914);
   U1917 : OAI22_X1 port map( A1 => n6558, A2 => n6596, B1 => n5090, B2 => 
                           n6597, ZN => n1913);
   U1918 : OAI22_X1 port map( A1 => n6559, A2 => n6596, B1 => n5091, B2 => 
                           n6597, ZN => n1912);
   U1919 : OAI22_X1 port map( A1 => n6560, A2 => n6596, B1 => n5092, B2 => 
                           n6597, ZN => n1911);
   U1920 : OAI22_X1 port map( A1 => n6528, A2 => n6598, B1 => n4709, B2 => 
                           n6599, ZN => n1910);
   U1921 : OAI22_X1 port map( A1 => n6530, A2 => n6598, B1 => n4710, B2 => 
                           n6599, ZN => n1909);
   U1922 : OAI22_X1 port map( A1 => n6531, A2 => n6598, B1 => n4711, B2 => 
                           n6599, ZN => n1908);
   U1923 : OAI22_X1 port map( A1 => n6532, A2 => n6598, B1 => n4712, B2 => 
                           n6599, ZN => n1907);
   U1924 : OAI22_X1 port map( A1 => n6533, A2 => n6598, B1 => n4713, B2 => 
                           n6599, ZN => n1906);
   U1925 : OAI22_X1 port map( A1 => n6534, A2 => n6598, B1 => n4714, B2 => 
                           n6599, ZN => n1905);
   U1926 : OAI22_X1 port map( A1 => n6535, A2 => n6598, B1 => n4715, B2 => 
                           n6599, ZN => n1904);
   U1927 : OAI22_X1 port map( A1 => n6536, A2 => n6598, B1 => n4716, B2 => 
                           n6599, ZN => n1903);
   U1928 : OAI22_X1 port map( A1 => n6537, A2 => n6598, B1 => n4717, B2 => 
                           n6599, ZN => n1902);
   U1929 : OAI22_X1 port map( A1 => n6538, A2 => n6598, B1 => n4718, B2 => 
                           n6599, ZN => n1901);
   U1930 : OAI22_X1 port map( A1 => n6539, A2 => n6598, B1 => n4719, B2 => 
                           n6599, ZN => n1900);
   U1931 : OAI22_X1 port map( A1 => n6540, A2 => n6598, B1 => n4720, B2 => 
                           n6599, ZN => n1899);
   U1932 : OAI22_X1 port map( A1 => n6541, A2 => n6598, B1 => n4721, B2 => 
                           n6599, ZN => n1898);
   U1933 : OAI22_X1 port map( A1 => n6542, A2 => n6598, B1 => n4722, B2 => 
                           n6599, ZN => n1897);
   U1934 : OAI22_X1 port map( A1 => n6543, A2 => n6598, B1 => n4723, B2 => 
                           n6599, ZN => n1896);
   U1935 : OAI22_X1 port map( A1 => n6544, A2 => n6598, B1 => n4724, B2 => 
                           n6599, ZN => n1895);
   U1936 : OAI22_X1 port map( A1 => n6545, A2 => n6598, B1 => n4725, B2 => 
                           n6599, ZN => n1894);
   U1937 : OAI22_X1 port map( A1 => n6546, A2 => n6598, B1 => n4726, B2 => 
                           n6599, ZN => n1893);
   U1938 : OAI22_X1 port map( A1 => n6547, A2 => n6598, B1 => n4727, B2 => 
                           n6599, ZN => n1892);
   U1939 : OAI22_X1 port map( A1 => n6548, A2 => n6598, B1 => n4728, B2 => 
                           n6599, ZN => n1891);
   U1940 : OAI22_X1 port map( A1 => n6549, A2 => n6598, B1 => n4729, B2 => 
                           n6599, ZN => n1890);
   U1941 : OAI22_X1 port map( A1 => n6550, A2 => n6598, B1 => n4730, B2 => 
                           n6599, ZN => n1889);
   U1942 : OAI22_X1 port map( A1 => n6551, A2 => n6598, B1 => n4731, B2 => 
                           n6599, ZN => n1888);
   U1943 : OAI22_X1 port map( A1 => n6552, A2 => n6598, B1 => n4732, B2 => 
                           n6599, ZN => n1887);
   U1944 : OAI22_X1 port map( A1 => n6553, A2 => n6598, B1 => n4733, B2 => 
                           n6599, ZN => n1886);
   U1945 : OAI22_X1 port map( A1 => n6554, A2 => n6598, B1 => n4734, B2 => 
                           n6599, ZN => n1885);
   U1946 : OAI22_X1 port map( A1 => n6555, A2 => n6598, B1 => n4735, B2 => 
                           n6599, ZN => n1884);
   U1947 : OAI22_X1 port map( A1 => n6556, A2 => n6598, B1 => n4736, B2 => 
                           n6599, ZN => n1883);
   U1948 : OAI22_X1 port map( A1 => n6557, A2 => n6598, B1 => n4737, B2 => 
                           n6599, ZN => n1882);
   U1949 : OAI22_X1 port map( A1 => n6558, A2 => n6598, B1 => n4738, B2 => 
                           n6599, ZN => n1881);
   U1950 : OAI22_X1 port map( A1 => n6559, A2 => n6598, B1 => n4739, B2 => 
                           n6599, ZN => n1880);
   U1951 : OAI22_X1 port map( A1 => n6560, A2 => n6598, B1 => n4740, B2 => 
                           n6599, ZN => n1879);
   U1952 : OAI22_X1 port map( A1 => n6528, A2 => n6600, B1 => n4451, B2 => 
                           n6601, ZN => n1878);
   U1953 : OAI22_X1 port map( A1 => n6530, A2 => n6600, B1 => n4452, B2 => 
                           n6601, ZN => n1877);
   U1954 : OAI22_X1 port map( A1 => n6531, A2 => n6600, B1 => n4453, B2 => 
                           n6601, ZN => n1876);
   U1955 : OAI22_X1 port map( A1 => n6532, A2 => n6600, B1 => n4454, B2 => 
                           n6601, ZN => n1875);
   U1956 : OAI22_X1 port map( A1 => n6533, A2 => n6600, B1 => n4455, B2 => 
                           n6601, ZN => n1874);
   U1957 : OAI22_X1 port map( A1 => n6534, A2 => n6600, B1 => n4456, B2 => 
                           n6601, ZN => n1873);
   U1958 : OAI22_X1 port map( A1 => n6535, A2 => n6600, B1 => n4457, B2 => 
                           n6601, ZN => n1872);
   U1959 : OAI22_X1 port map( A1 => n6536, A2 => n6600, B1 => n4458, B2 => 
                           n6601, ZN => n1871);
   U1960 : OAI22_X1 port map( A1 => n6537, A2 => n6600, B1 => n4459, B2 => 
                           n6601, ZN => n1870);
   U1961 : OAI22_X1 port map( A1 => n6538, A2 => n6600, B1 => n4460, B2 => 
                           n6601, ZN => n1869);
   U1962 : OAI22_X1 port map( A1 => n6539, A2 => n6600, B1 => n4461, B2 => 
                           n6601, ZN => n1868);
   U1963 : OAI22_X1 port map( A1 => n6540, A2 => n6600, B1 => n4462, B2 => 
                           n6601, ZN => n1867);
   U1964 : OAI22_X1 port map( A1 => n6541, A2 => n6600, B1 => n4463, B2 => 
                           n6601, ZN => n1866);
   U1965 : OAI22_X1 port map( A1 => n6542, A2 => n6600, B1 => n4464, B2 => 
                           n6601, ZN => n1865);
   U1966 : OAI22_X1 port map( A1 => n6543, A2 => n6600, B1 => n4465, B2 => 
                           n6601, ZN => n1864);
   U1967 : OAI22_X1 port map( A1 => n6544, A2 => n6600, B1 => n4466, B2 => 
                           n6601, ZN => n1863);
   U1968 : OAI22_X1 port map( A1 => n6545, A2 => n6600, B1 => n4467, B2 => 
                           n6601, ZN => n1862);
   U1969 : OAI22_X1 port map( A1 => n6546, A2 => n6600, B1 => n4468, B2 => 
                           n6601, ZN => n1861);
   U1970 : OAI22_X1 port map( A1 => n6547, A2 => n6600, B1 => n4469, B2 => 
                           n6601, ZN => n1860);
   U1971 : OAI22_X1 port map( A1 => n6548, A2 => n6600, B1 => n4470, B2 => 
                           n6601, ZN => n1859);
   U1972 : OAI22_X1 port map( A1 => n6549, A2 => n6600, B1 => n4471, B2 => 
                           n6601, ZN => n1858);
   U1973 : OAI22_X1 port map( A1 => n6550, A2 => n6600, B1 => n4472, B2 => 
                           n6601, ZN => n1857);
   U1974 : OAI22_X1 port map( A1 => n6551, A2 => n6600, B1 => n4473, B2 => 
                           n6601, ZN => n1856);
   U1975 : OAI22_X1 port map( A1 => n6552, A2 => n6600, B1 => n4474, B2 => 
                           n6601, ZN => n1855);
   U1976 : OAI22_X1 port map( A1 => n6553, A2 => n6600, B1 => n4475, B2 => 
                           n6601, ZN => n1854);
   U1977 : OAI22_X1 port map( A1 => n6554, A2 => n6600, B1 => n4476, B2 => 
                           n6601, ZN => n1853);
   U1978 : OAI22_X1 port map( A1 => n6555, A2 => n6600, B1 => n4477, B2 => 
                           n6601, ZN => n1852);
   U1979 : OAI22_X1 port map( A1 => n6556, A2 => n6600, B1 => n4478, B2 => 
                           n6601, ZN => n1851);
   U1980 : OAI22_X1 port map( A1 => n6557, A2 => n6600, B1 => n4479, B2 => 
                           n6601, ZN => n1850);
   U1981 : OAI22_X1 port map( A1 => n6558, A2 => n6600, B1 => n4480, B2 => 
                           n6601, ZN => n1849);
   U1982 : OAI22_X1 port map( A1 => n6559, A2 => n6600, B1 => n4481, B2 => 
                           n6601, ZN => n1848);
   U1983 : OAI22_X1 port map( A1 => n6560, A2 => n6600, B1 => n4482, B2 => 
                           n6601, ZN => n1847);
   U1984 : OAI22_X1 port map( A1 => n6528, A2 => n6602, B1 => n4837, B2 => 
                           n6603, ZN => n1846);
   U1985 : OAI22_X1 port map( A1 => n6530, A2 => n6602, B1 => n4838, B2 => 
                           n6603, ZN => n1845);
   U1986 : OAI22_X1 port map( A1 => n6531, A2 => n6602, B1 => n4839, B2 => 
                           n6603, ZN => n1844);
   U1987 : OAI22_X1 port map( A1 => n6532, A2 => n6602, B1 => n4840, B2 => 
                           n6603, ZN => n1843);
   U1988 : OAI22_X1 port map( A1 => n6533, A2 => n6602, B1 => n4841, B2 => 
                           n6603, ZN => n1842);
   U1989 : OAI22_X1 port map( A1 => n6534, A2 => n6602, B1 => n4842, B2 => 
                           n6603, ZN => n1841);
   U1990 : OAI22_X1 port map( A1 => n6535, A2 => n6602, B1 => n4843, B2 => 
                           n6603, ZN => n1840);
   U1991 : OAI22_X1 port map( A1 => n6536, A2 => n6602, B1 => n4844, B2 => 
                           n6603, ZN => n1839);
   U1992 : OAI22_X1 port map( A1 => n6537, A2 => n6602, B1 => n4845, B2 => 
                           n6603, ZN => n1838);
   U1993 : OAI22_X1 port map( A1 => n6538, A2 => n6602, B1 => n4846, B2 => 
                           n6603, ZN => n1837);
   U1994 : OAI22_X1 port map( A1 => n6539, A2 => n6602, B1 => n4847, B2 => 
                           n6603, ZN => n1836);
   U1995 : OAI22_X1 port map( A1 => n6540, A2 => n6602, B1 => n4848, B2 => 
                           n6603, ZN => n1835);
   U1996 : OAI22_X1 port map( A1 => n6541, A2 => n6602, B1 => n4849, B2 => 
                           n6603, ZN => n1834);
   U1997 : OAI22_X1 port map( A1 => n6542, A2 => n6602, B1 => n4850, B2 => 
                           n6603, ZN => n1833);
   U1998 : OAI22_X1 port map( A1 => n6543, A2 => n6602, B1 => n4851, B2 => 
                           n6603, ZN => n1832);
   U1999 : OAI22_X1 port map( A1 => n6544, A2 => n6602, B1 => n4852, B2 => 
                           n6603, ZN => n1831);
   U2000 : OAI22_X1 port map( A1 => n6545, A2 => n6602, B1 => n4853, B2 => 
                           n6603, ZN => n1830);
   U2001 : OAI22_X1 port map( A1 => n6546, A2 => n6602, B1 => n4854, B2 => 
                           n6603, ZN => n1829);
   U2002 : OAI22_X1 port map( A1 => n6547, A2 => n6602, B1 => n4855, B2 => 
                           n6603, ZN => n1828);
   U2003 : OAI22_X1 port map( A1 => n6548, A2 => n6602, B1 => n4856, B2 => 
                           n6603, ZN => n1827);
   U2004 : OAI22_X1 port map( A1 => n6549, A2 => n6602, B1 => n4857, B2 => 
                           n6603, ZN => n1826);
   U2005 : OAI22_X1 port map( A1 => n6550, A2 => n6602, B1 => n4858, B2 => 
                           n6603, ZN => n1825);
   U2006 : OAI22_X1 port map( A1 => n6551, A2 => n6602, B1 => n4859, B2 => 
                           n6603, ZN => n1824);
   U2007 : OAI22_X1 port map( A1 => n6552, A2 => n6602, B1 => n4860, B2 => 
                           n6603, ZN => n1823);
   U2008 : OAI22_X1 port map( A1 => n6553, A2 => n6602, B1 => n4861, B2 => 
                           n6603, ZN => n1822);
   U2009 : OAI22_X1 port map( A1 => n6554, A2 => n6602, B1 => n4862, B2 => 
                           n6603, ZN => n1821);
   U2010 : OAI22_X1 port map( A1 => n6555, A2 => n6602, B1 => n4863, B2 => 
                           n6603, ZN => n1820);
   U2011 : OAI22_X1 port map( A1 => n6556, A2 => n6602, B1 => n4864, B2 => 
                           n6603, ZN => n1819);
   U2012 : OAI22_X1 port map( A1 => n6557, A2 => n6602, B1 => n4865, B2 => 
                           n6603, ZN => n1818);
   U2013 : OAI22_X1 port map( A1 => n6558, A2 => n6602, B1 => n4866, B2 => 
                           n6603, ZN => n1817);
   U2014 : OAI22_X1 port map( A1 => n6559, A2 => n6602, B1 => n4867, B2 => 
                           n6603, ZN => n1816);
   U2015 : OAI22_X1 port map( A1 => n6560, A2 => n6602, B1 => n4868, B2 => 
                           n6603, ZN => n1815);
   U2016 : AND3_X1 port map( A1 => n6586, A2 => n6585, A3 => ADD_WR(3), ZN => 
                           n6589);
   U2017 : INV_X1 port map( A => ADD_WR(4), ZN => n6585);
   U2018 : OAI22_X1 port map( A1 => n6528, A2 => n6604, B1 => n5093, B2 => 
                           n6605, ZN => n1814);
   U2019 : OAI22_X1 port map( A1 => n6530, A2 => n6604, B1 => n5094, B2 => 
                           n6605, ZN => n1813);
   U2020 : OAI22_X1 port map( A1 => n6531, A2 => n6604, B1 => n5095, B2 => 
                           n6605, ZN => n1812);
   U2021 : OAI22_X1 port map( A1 => n6532, A2 => n6604, B1 => n5096, B2 => 
                           n6605, ZN => n1811);
   U2022 : OAI22_X1 port map( A1 => n6533, A2 => n6604, B1 => n5097, B2 => 
                           n6605, ZN => n1810);
   U2023 : OAI22_X1 port map( A1 => n6534, A2 => n6604, B1 => n5098, B2 => 
                           n6605, ZN => n1809);
   U2024 : OAI22_X1 port map( A1 => n6535, A2 => n6604, B1 => n5099, B2 => 
                           n6605, ZN => n1808);
   U2025 : OAI22_X1 port map( A1 => n6536, A2 => n6604, B1 => n5100, B2 => 
                           n6605, ZN => n1807);
   U2026 : OAI22_X1 port map( A1 => n6537, A2 => n6604, B1 => n5101, B2 => 
                           n6605, ZN => n1806);
   U2027 : OAI22_X1 port map( A1 => n6538, A2 => n6604, B1 => n5102, B2 => 
                           n6605, ZN => n1805);
   U2028 : OAI22_X1 port map( A1 => n6539, A2 => n6604, B1 => n5103, B2 => 
                           n6605, ZN => n1804);
   U2029 : OAI22_X1 port map( A1 => n6540, A2 => n6604, B1 => n5104, B2 => 
                           n6605, ZN => n1803);
   U2030 : OAI22_X1 port map( A1 => n6541, A2 => n6604, B1 => n5105, B2 => 
                           n6605, ZN => n1802);
   U2031 : OAI22_X1 port map( A1 => n6542, A2 => n6604, B1 => n5106, B2 => 
                           n6605, ZN => n1801);
   U2032 : OAI22_X1 port map( A1 => n6543, A2 => n6604, B1 => n5107, B2 => 
                           n6605, ZN => n1800);
   U2033 : OAI22_X1 port map( A1 => n6544, A2 => n6604, B1 => n5108, B2 => 
                           n6605, ZN => n1799);
   U2034 : OAI22_X1 port map( A1 => n6545, A2 => n6604, B1 => n5109, B2 => 
                           n6605, ZN => n1798);
   U2035 : OAI22_X1 port map( A1 => n6546, A2 => n6604, B1 => n5110, B2 => 
                           n6605, ZN => n1797);
   U2036 : OAI22_X1 port map( A1 => n6547, A2 => n6604, B1 => n5111, B2 => 
                           n6605, ZN => n1796);
   U2037 : OAI22_X1 port map( A1 => n6548, A2 => n6604, B1 => n5112, B2 => 
                           n6605, ZN => n1795);
   U2038 : OAI22_X1 port map( A1 => n6549, A2 => n6604, B1 => n5113, B2 => 
                           n6605, ZN => n1794);
   U2039 : OAI22_X1 port map( A1 => n6550, A2 => n6604, B1 => n5114, B2 => 
                           n6605, ZN => n1793);
   U2040 : OAI22_X1 port map( A1 => n6551, A2 => n6604, B1 => n5115, B2 => 
                           n6605, ZN => n1792);
   U2041 : OAI22_X1 port map( A1 => n6552, A2 => n6604, B1 => n5116, B2 => 
                           n6605, ZN => n1791);
   U2042 : OAI22_X1 port map( A1 => n6553, A2 => n6604, B1 => n5117, B2 => 
                           n6605, ZN => n1790);
   U2043 : OAI22_X1 port map( A1 => n6554, A2 => n6604, B1 => n5118, B2 => 
                           n6605, ZN => n1789);
   U2044 : OAI22_X1 port map( A1 => n6555, A2 => n6604, B1 => n5119, B2 => 
                           n6605, ZN => n1788);
   U2045 : OAI22_X1 port map( A1 => n6556, A2 => n6604, B1 => n5120, B2 => 
                           n6605, ZN => n1787);
   U2046 : OAI22_X1 port map( A1 => n6557, A2 => n6604, B1 => n5121, B2 => 
                           n6605, ZN => n1786);
   U2047 : OAI22_X1 port map( A1 => n6558, A2 => n6604, B1 => n5122, B2 => 
                           n6605, ZN => n1785);
   U2048 : OAI22_X1 port map( A1 => n6559, A2 => n6604, B1 => n5123, B2 => 
                           n6605, ZN => n1784);
   U2049 : OAI22_X1 port map( A1 => n6560, A2 => n6604, B1 => n5124, B2 => 
                           n6605, ZN => n1783);
   U2050 : OAI22_X1 port map( A1 => n6528, A2 => n6607, B1 => n4517, B2 => 
                           n6608, ZN => n1782);
   U2051 : OAI22_X1 port map( A1 => n6530, A2 => n6607, B1 => n4518, B2 => 
                           n6608, ZN => n1781);
   U2052 : OAI22_X1 port map( A1 => n6531, A2 => n6607, B1 => n4519, B2 => 
                           n6608, ZN => n1780);
   U2053 : OAI22_X1 port map( A1 => n6532, A2 => n6607, B1 => n4520, B2 => 
                           n6608, ZN => n1779);
   U2054 : OAI22_X1 port map( A1 => n6533, A2 => n6607, B1 => n4521, B2 => 
                           n6608, ZN => n1778);
   U2055 : OAI22_X1 port map( A1 => n6534, A2 => n6607, B1 => n4522, B2 => 
                           n6608, ZN => n1777);
   U2056 : OAI22_X1 port map( A1 => n6535, A2 => n6607, B1 => n4523, B2 => 
                           n6608, ZN => n1776);
   U2057 : OAI22_X1 port map( A1 => n6536, A2 => n6607, B1 => n4524, B2 => 
                           n6608, ZN => n1775);
   U2058 : OAI22_X1 port map( A1 => n6537, A2 => n6607, B1 => n4525, B2 => 
                           n6608, ZN => n1774);
   U2059 : OAI22_X1 port map( A1 => n6538, A2 => n6607, B1 => n4526, B2 => 
                           n6608, ZN => n1773);
   U2060 : OAI22_X1 port map( A1 => n6539, A2 => n6607, B1 => n4527, B2 => 
                           n6608, ZN => n1772);
   U2061 : OAI22_X1 port map( A1 => n6540, A2 => n6607, B1 => n4528, B2 => 
                           n6608, ZN => n1771);
   U2062 : OAI22_X1 port map( A1 => n6541, A2 => n6607, B1 => n4529, B2 => 
                           n6608, ZN => n1770);
   U2063 : OAI22_X1 port map( A1 => n6542, A2 => n6607, B1 => n4530, B2 => 
                           n6608, ZN => n1769);
   U2064 : OAI22_X1 port map( A1 => n6543, A2 => n6607, B1 => n4531, B2 => 
                           n6608, ZN => n1768);
   U2065 : OAI22_X1 port map( A1 => n6544, A2 => n6607, B1 => n4532, B2 => 
                           n6608, ZN => n1767);
   U2066 : OAI22_X1 port map( A1 => n6545, A2 => n6607, B1 => n4533, B2 => 
                           n6608, ZN => n1766);
   U2067 : OAI22_X1 port map( A1 => n6546, A2 => n6607, B1 => n4534, B2 => 
                           n6608, ZN => n1765);
   U2068 : OAI22_X1 port map( A1 => n6547, A2 => n6607, B1 => n4535, B2 => 
                           n6608, ZN => n1764);
   U2069 : OAI22_X1 port map( A1 => n6548, A2 => n6607, B1 => n4536, B2 => 
                           n6608, ZN => n1763);
   U2070 : OAI22_X1 port map( A1 => n6549, A2 => n6607, B1 => n4537, B2 => 
                           n6608, ZN => n1762);
   U2071 : OAI22_X1 port map( A1 => n6550, A2 => n6607, B1 => n4538, B2 => 
                           n6608, ZN => n1761);
   U2072 : OAI22_X1 port map( A1 => n6551, A2 => n6607, B1 => n4539, B2 => 
                           n6608, ZN => n1760);
   U2073 : OAI22_X1 port map( A1 => n6552, A2 => n6607, B1 => n4540, B2 => 
                           n6608, ZN => n1759);
   U2074 : OAI22_X1 port map( A1 => n6553, A2 => n6607, B1 => n4541, B2 => 
                           n6608, ZN => n1758);
   U2075 : OAI22_X1 port map( A1 => n6554, A2 => n6607, B1 => n4542, B2 => 
                           n6608, ZN => n1757);
   U2076 : OAI22_X1 port map( A1 => n6555, A2 => n6607, B1 => n4543, B2 => 
                           n6608, ZN => n1756);
   U2077 : OAI22_X1 port map( A1 => n6556, A2 => n6607, B1 => n4544, B2 => 
                           n6608, ZN => n1755);
   U2078 : OAI22_X1 port map( A1 => n6557, A2 => n6607, B1 => n4545, B2 => 
                           n6608, ZN => n1754);
   U2079 : OAI22_X1 port map( A1 => n6558, A2 => n6607, B1 => n4546, B2 => 
                           n6608, ZN => n1753);
   U2080 : OAI22_X1 port map( A1 => n6559, A2 => n6607, B1 => n4547, B2 => 
                           n6608, ZN => n1752);
   U2081 : OAI22_X1 port map( A1 => n6560, A2 => n6607, B1 => n4548, B2 => 
                           n6608, ZN => n1751);
   U2082 : OAI22_X1 port map( A1 => n6528, A2 => n6609, B1 => n5125, B2 => 
                           n6610, ZN => n1750);
   U2083 : OAI22_X1 port map( A1 => n6530, A2 => n6609, B1 => n5126, B2 => 
                           n6610, ZN => n1749);
   U2084 : OAI22_X1 port map( A1 => n6531, A2 => n6609, B1 => n5127, B2 => 
                           n6610, ZN => n1748);
   U2085 : OAI22_X1 port map( A1 => n6532, A2 => n6609, B1 => n5128, B2 => 
                           n6610, ZN => n1747);
   U2086 : OAI22_X1 port map( A1 => n6533, A2 => n6609, B1 => n5129, B2 => 
                           n6610, ZN => n1746);
   U2087 : OAI22_X1 port map( A1 => n6534, A2 => n6609, B1 => n5130, B2 => 
                           n6610, ZN => n1745);
   U2088 : OAI22_X1 port map( A1 => n6535, A2 => n6609, B1 => n5131, B2 => 
                           n6610, ZN => n1744);
   U2089 : OAI22_X1 port map( A1 => n6536, A2 => n6609, B1 => n5132, B2 => 
                           n6610, ZN => n1743);
   U2090 : OAI22_X1 port map( A1 => n6537, A2 => n6609, B1 => n5133, B2 => 
                           n6610, ZN => n1742);
   U2091 : OAI22_X1 port map( A1 => n6538, A2 => n6609, B1 => n5134, B2 => 
                           n6610, ZN => n1741);
   U2092 : OAI22_X1 port map( A1 => n6539, A2 => n6609, B1 => n5135, B2 => 
                           n6610, ZN => n1740);
   U2093 : OAI22_X1 port map( A1 => n6540, A2 => n6609, B1 => n5136, B2 => 
                           n6610, ZN => n1739);
   U2094 : OAI22_X1 port map( A1 => n6541, A2 => n6609, B1 => n5137, B2 => 
                           n6610, ZN => n1738);
   U2095 : OAI22_X1 port map( A1 => n6542, A2 => n6609, B1 => n5138, B2 => 
                           n6610, ZN => n1737);
   U2096 : OAI22_X1 port map( A1 => n6543, A2 => n6609, B1 => n5139, B2 => 
                           n6610, ZN => n1736);
   U2097 : OAI22_X1 port map( A1 => n6544, A2 => n6609, B1 => n5140, B2 => 
                           n6610, ZN => n1735);
   U2098 : OAI22_X1 port map( A1 => n6545, A2 => n6609, B1 => n5141, B2 => 
                           n6610, ZN => n1734);
   U2099 : OAI22_X1 port map( A1 => n6546, A2 => n6609, B1 => n5142, B2 => 
                           n6610, ZN => n1733);
   U2100 : OAI22_X1 port map( A1 => n6547, A2 => n6609, B1 => n5143, B2 => 
                           n6610, ZN => n1732);
   U2101 : OAI22_X1 port map( A1 => n6548, A2 => n6609, B1 => n5144, B2 => 
                           n6610, ZN => n1731);
   U2102 : OAI22_X1 port map( A1 => n6549, A2 => n6609, B1 => n5145, B2 => 
                           n6610, ZN => n1730);
   U2103 : OAI22_X1 port map( A1 => n6550, A2 => n6609, B1 => n5146, B2 => 
                           n6610, ZN => n1729);
   U2104 : OAI22_X1 port map( A1 => n6551, A2 => n6609, B1 => n5147, B2 => 
                           n6610, ZN => n1728);
   U2105 : OAI22_X1 port map( A1 => n6552, A2 => n6609, B1 => n5148, B2 => 
                           n6610, ZN => n1727);
   U2106 : OAI22_X1 port map( A1 => n6553, A2 => n6609, B1 => n5149, B2 => 
                           n6610, ZN => n1726);
   U2107 : OAI22_X1 port map( A1 => n6554, A2 => n6609, B1 => n5150, B2 => 
                           n6610, ZN => n1725);
   U2108 : OAI22_X1 port map( A1 => n6555, A2 => n6609, B1 => n5151, B2 => 
                           n6610, ZN => n1724);
   U2109 : OAI22_X1 port map( A1 => n6556, A2 => n6609, B1 => n5152, B2 => 
                           n6610, ZN => n1723);
   U2110 : OAI22_X1 port map( A1 => n6557, A2 => n6609, B1 => n5153, B2 => 
                           n6610, ZN => n1722);
   U2111 : OAI22_X1 port map( A1 => n6558, A2 => n6609, B1 => n5154, B2 => 
                           n6610, ZN => n1721);
   U2112 : OAI22_X1 port map( A1 => n6559, A2 => n6609, B1 => n5155, B2 => 
                           n6610, ZN => n1720);
   U2113 : OAI22_X1 port map( A1 => n6560, A2 => n6609, B1 => n5156, B2 => 
                           n6610, ZN => n1719);
   U2114 : OAI22_X1 port map( A1 => n6528, A2 => n6611, B1 => n4869, B2 => 
                           n6612, ZN => n1718);
   U2115 : OAI22_X1 port map( A1 => n6530, A2 => n6611, B1 => n4870, B2 => 
                           n6612, ZN => n1717);
   U2116 : OAI22_X1 port map( A1 => n6531, A2 => n6611, B1 => n4871, B2 => 
                           n6612, ZN => n1716);
   U2117 : OAI22_X1 port map( A1 => n6532, A2 => n6611, B1 => n4872, B2 => 
                           n6612, ZN => n1715);
   U2118 : OAI22_X1 port map( A1 => n6533, A2 => n6611, B1 => n4873, B2 => 
                           n6612, ZN => n1714);
   U2119 : OAI22_X1 port map( A1 => n6534, A2 => n6611, B1 => n4874, B2 => 
                           n6612, ZN => n1713);
   U2120 : OAI22_X1 port map( A1 => n6535, A2 => n6611, B1 => n4875, B2 => 
                           n6612, ZN => n1712);
   U2121 : OAI22_X1 port map( A1 => n6536, A2 => n6611, B1 => n4876, B2 => 
                           n6612, ZN => n1711);
   U2122 : OAI22_X1 port map( A1 => n6537, A2 => n6611, B1 => n4877, B2 => 
                           n6612, ZN => n1710);
   U2123 : OAI22_X1 port map( A1 => n6538, A2 => n6611, B1 => n4878, B2 => 
                           n6612, ZN => n1709);
   U2124 : OAI22_X1 port map( A1 => n6539, A2 => n6611, B1 => n4879, B2 => 
                           n6612, ZN => n1708);
   U2125 : OAI22_X1 port map( A1 => n6540, A2 => n6611, B1 => n4880, B2 => 
                           n6612, ZN => n1707);
   U2126 : OAI22_X1 port map( A1 => n6541, A2 => n6611, B1 => n4881, B2 => 
                           n6612, ZN => n1706);
   U2127 : OAI22_X1 port map( A1 => n6542, A2 => n6611, B1 => n4882, B2 => 
                           n6612, ZN => n1705);
   U2128 : OAI22_X1 port map( A1 => n6543, A2 => n6611, B1 => n4883, B2 => 
                           n6612, ZN => n1704);
   U2129 : OAI22_X1 port map( A1 => n6544, A2 => n6611, B1 => n4884, B2 => 
                           n6612, ZN => n1703);
   U2130 : OAI22_X1 port map( A1 => n6545, A2 => n6611, B1 => n4885, B2 => 
                           n6612, ZN => n1702);
   U2131 : OAI22_X1 port map( A1 => n6546, A2 => n6611, B1 => n4886, B2 => 
                           n6612, ZN => n1701);
   U2132 : OAI22_X1 port map( A1 => n6547, A2 => n6611, B1 => n4887, B2 => 
                           n6612, ZN => n1700);
   U2133 : OAI22_X1 port map( A1 => n6548, A2 => n6611, B1 => n4888, B2 => 
                           n6612, ZN => n1699);
   U2134 : OAI22_X1 port map( A1 => n6549, A2 => n6611, B1 => n4889, B2 => 
                           n6612, ZN => n1698);
   U2135 : OAI22_X1 port map( A1 => n6550, A2 => n6611, B1 => n4890, B2 => 
                           n6612, ZN => n1697);
   U2136 : OAI22_X1 port map( A1 => n6551, A2 => n6611, B1 => n4891, B2 => 
                           n6612, ZN => n1696);
   U2137 : OAI22_X1 port map( A1 => n6552, A2 => n6611, B1 => n4892, B2 => 
                           n6612, ZN => n1695);
   U2138 : OAI22_X1 port map( A1 => n6553, A2 => n6611, B1 => n4893, B2 => 
                           n6612, ZN => n1694);
   U2139 : OAI22_X1 port map( A1 => n6554, A2 => n6611, B1 => n4894, B2 => 
                           n6612, ZN => n1693);
   U2140 : OAI22_X1 port map( A1 => n6555, A2 => n6611, B1 => n4895, B2 => 
                           n6612, ZN => n1692);
   U2141 : OAI22_X1 port map( A1 => n6556, A2 => n6611, B1 => n4896, B2 => 
                           n6612, ZN => n1691);
   U2142 : OAI22_X1 port map( A1 => n6557, A2 => n6611, B1 => n4897, B2 => 
                           n6612, ZN => n1690);
   U2143 : OAI22_X1 port map( A1 => n6558, A2 => n6611, B1 => n4898, B2 => 
                           n6612, ZN => n1689);
   U2144 : OAI22_X1 port map( A1 => n6559, A2 => n6611, B1 => n4899, B2 => 
                           n6612, ZN => n1688);
   U2145 : OAI22_X1 port map( A1 => n6560, A2 => n6611, B1 => n4900, B2 => 
                           n6612, ZN => n1687);
   U2146 : OAI22_X1 port map( A1 => n6528, A2 => n6613, B1 => n4259, B2 => 
                           n6614, ZN => n1686);
   U2147 : OAI22_X1 port map( A1 => n6530, A2 => n6613, B1 => n4260, B2 => 
                           n6614, ZN => n1685);
   U2148 : OAI22_X1 port map( A1 => n6531, A2 => n6613, B1 => n4261, B2 => 
                           n6614, ZN => n1684);
   U2149 : OAI22_X1 port map( A1 => n6532, A2 => n6613, B1 => n4262, B2 => 
                           n6614, ZN => n1683);
   U2150 : OAI22_X1 port map( A1 => n6533, A2 => n6613, B1 => n4263, B2 => 
                           n6614, ZN => n1682);
   U2151 : OAI22_X1 port map( A1 => n6534, A2 => n6613, B1 => n4264, B2 => 
                           n6614, ZN => n1681);
   U2152 : OAI22_X1 port map( A1 => n6535, A2 => n6613, B1 => n4265, B2 => 
                           n6614, ZN => n1680);
   U2153 : OAI22_X1 port map( A1 => n6536, A2 => n6613, B1 => n4266, B2 => 
                           n6614, ZN => n1679);
   U2154 : OAI22_X1 port map( A1 => n6537, A2 => n6613, B1 => n4267, B2 => 
                           n6614, ZN => n1678);
   U2155 : OAI22_X1 port map( A1 => n6538, A2 => n6613, B1 => n4268, B2 => 
                           n6614, ZN => n1677);
   U2156 : OAI22_X1 port map( A1 => n6539, A2 => n6613, B1 => n4269, B2 => 
                           n6614, ZN => n1676);
   U2157 : OAI22_X1 port map( A1 => n6540, A2 => n6613, B1 => n4270, B2 => 
                           n6614, ZN => n1675);
   U2158 : OAI22_X1 port map( A1 => n6541, A2 => n6613, B1 => n4271, B2 => 
                           n6614, ZN => n1674);
   U2159 : OAI22_X1 port map( A1 => n6542, A2 => n6613, B1 => n4272, B2 => 
                           n6614, ZN => n1673);
   U2160 : OAI22_X1 port map( A1 => n6543, A2 => n6613, B1 => n4273, B2 => 
                           n6614, ZN => n1672);
   U2161 : OAI22_X1 port map( A1 => n6544, A2 => n6613, B1 => n4274, B2 => 
                           n6614, ZN => n1671);
   U2162 : OAI22_X1 port map( A1 => n6545, A2 => n6613, B1 => n4275, B2 => 
                           n6614, ZN => n1670);
   U2163 : OAI22_X1 port map( A1 => n6546, A2 => n6613, B1 => n4276, B2 => 
                           n6614, ZN => n1669);
   U2164 : OAI22_X1 port map( A1 => n6547, A2 => n6613, B1 => n4277, B2 => 
                           n6614, ZN => n1668);
   U2165 : OAI22_X1 port map( A1 => n6548, A2 => n6613, B1 => n4278, B2 => 
                           n6614, ZN => n1667);
   U2166 : OAI22_X1 port map( A1 => n6549, A2 => n6613, B1 => n4279, B2 => 
                           n6614, ZN => n1666);
   U2167 : OAI22_X1 port map( A1 => n6550, A2 => n6613, B1 => n4280, B2 => 
                           n6614, ZN => n1665);
   U2168 : OAI22_X1 port map( A1 => n6551, A2 => n6613, B1 => n4281, B2 => 
                           n6614, ZN => n1664);
   U2169 : OAI22_X1 port map( A1 => n6552, A2 => n6613, B1 => n4282, B2 => 
                           n6614, ZN => n1663);
   U2170 : OAI22_X1 port map( A1 => n6553, A2 => n6613, B1 => n4283, B2 => 
                           n6614, ZN => n1662);
   U2171 : OAI22_X1 port map( A1 => n6554, A2 => n6613, B1 => n4284, B2 => 
                           n6614, ZN => n1661);
   U2172 : OAI22_X1 port map( A1 => n6555, A2 => n6613, B1 => n4285, B2 => 
                           n6614, ZN => n1660);
   U2173 : OAI22_X1 port map( A1 => n6556, A2 => n6613, B1 => n4286, B2 => 
                           n6614, ZN => n1659);
   U2174 : OAI22_X1 port map( A1 => n6557, A2 => n6613, B1 => n4287, B2 => 
                           n6614, ZN => n1658);
   U2175 : OAI22_X1 port map( A1 => n6558, A2 => n6613, B1 => n4288, B2 => 
                           n6614, ZN => n1657);
   U2176 : OAI22_X1 port map( A1 => n6559, A2 => n6613, B1 => n4289, B2 => 
                           n6614, ZN => n1656);
   U2177 : OAI22_X1 port map( A1 => n6560, A2 => n6613, B1 => n4290, B2 => 
                           n6614, ZN => n1655);
   U2178 : OAI22_X1 port map( A1 => n6528, A2 => n6615, B1 => n4291, B2 => 
                           n6616, ZN => n1654);
   U2179 : OAI22_X1 port map( A1 => n6530, A2 => n6615, B1 => n4292, B2 => 
                           n6616, ZN => n1653);
   U2180 : OAI22_X1 port map( A1 => n6531, A2 => n6615, B1 => n4293, B2 => 
                           n6616, ZN => n1652);
   U2181 : OAI22_X1 port map( A1 => n6532, A2 => n6615, B1 => n4294, B2 => 
                           n6616, ZN => n1651);
   U2182 : OAI22_X1 port map( A1 => n6533, A2 => n6615, B1 => n4295, B2 => 
                           n6616, ZN => n1650);
   U2183 : OAI22_X1 port map( A1 => n6534, A2 => n6615, B1 => n4296, B2 => 
                           n6616, ZN => n1649);
   U2184 : OAI22_X1 port map( A1 => n6535, A2 => n6615, B1 => n4297, B2 => 
                           n6616, ZN => n1648);
   U2185 : OAI22_X1 port map( A1 => n6536, A2 => n6615, B1 => n4298, B2 => 
                           n6616, ZN => n1647);
   U2186 : OAI22_X1 port map( A1 => n6537, A2 => n6615, B1 => n4299, B2 => 
                           n6616, ZN => n1646);
   U2187 : OAI22_X1 port map( A1 => n6538, A2 => n6615, B1 => n4300, B2 => 
                           n6616, ZN => n1645);
   U2188 : OAI22_X1 port map( A1 => n6539, A2 => n6615, B1 => n4301, B2 => 
                           n6616, ZN => n1644);
   U2189 : OAI22_X1 port map( A1 => n6540, A2 => n6615, B1 => n4302, B2 => 
                           n6616, ZN => n1643);
   U2190 : OAI22_X1 port map( A1 => n6541, A2 => n6615, B1 => n4303, B2 => 
                           n6616, ZN => n1642);
   U2191 : OAI22_X1 port map( A1 => n6542, A2 => n6615, B1 => n4304, B2 => 
                           n6616, ZN => n1641);
   U2192 : OAI22_X1 port map( A1 => n6543, A2 => n6615, B1 => n4305, B2 => 
                           n6616, ZN => n1640);
   U2193 : OAI22_X1 port map( A1 => n6544, A2 => n6615, B1 => n4306, B2 => 
                           n6616, ZN => n1639);
   U2194 : OAI22_X1 port map( A1 => n6545, A2 => n6615, B1 => n4307, B2 => 
                           n6616, ZN => n1638);
   U2195 : OAI22_X1 port map( A1 => n6546, A2 => n6615, B1 => n4308, B2 => 
                           n6616, ZN => n1637);
   U2196 : OAI22_X1 port map( A1 => n6547, A2 => n6615, B1 => n4309, B2 => 
                           n6616, ZN => n1636);
   U2197 : OAI22_X1 port map( A1 => n6548, A2 => n6615, B1 => n4310, B2 => 
                           n6616, ZN => n1635);
   U2198 : OAI22_X1 port map( A1 => n6549, A2 => n6615, B1 => n4311, B2 => 
                           n6616, ZN => n1634);
   U2199 : OAI22_X1 port map( A1 => n6550, A2 => n6615, B1 => n4312, B2 => 
                           n6616, ZN => n1633);
   U2200 : OAI22_X1 port map( A1 => n6551, A2 => n6615, B1 => n4313, B2 => 
                           n6616, ZN => n1632);
   U2201 : OAI22_X1 port map( A1 => n6552, A2 => n6615, B1 => n4314, B2 => 
                           n6616, ZN => n1631);
   U2202 : OAI22_X1 port map( A1 => n6553, A2 => n6615, B1 => n4315, B2 => 
                           n6616, ZN => n1630);
   U2203 : OAI22_X1 port map( A1 => n6554, A2 => n6615, B1 => n4316, B2 => 
                           n6616, ZN => n1629);
   U2204 : OAI22_X1 port map( A1 => n6555, A2 => n6615, B1 => n4317, B2 => 
                           n6616, ZN => n1628);
   U2205 : OAI22_X1 port map( A1 => n6556, A2 => n6615, B1 => n4318, B2 => 
                           n6616, ZN => n1627);
   U2206 : OAI22_X1 port map( A1 => n6557, A2 => n6615, B1 => n4319, B2 => 
                           n6616, ZN => n1626);
   U2207 : OAI22_X1 port map( A1 => n6558, A2 => n6615, B1 => n4320, B2 => 
                           n6616, ZN => n1625);
   U2208 : OAI22_X1 port map( A1 => n6559, A2 => n6615, B1 => n4321, B2 => 
                           n6616, ZN => n1624);
   U2209 : OAI22_X1 port map( A1 => n6560, A2 => n6615, B1 => n4322, B2 => 
                           n6616, ZN => n1623);
   U2210 : OAI22_X1 port map( A1 => n6528, A2 => n6617, B1 => n4901, B2 => 
                           n6618, ZN => n1622);
   U2211 : OAI22_X1 port map( A1 => n6530, A2 => n6617, B1 => n4902, B2 => 
                           n6618, ZN => n1621);
   U2212 : OAI22_X1 port map( A1 => n6531, A2 => n6617, B1 => n4903, B2 => 
                           n6618, ZN => n1620);
   U2213 : OAI22_X1 port map( A1 => n6532, A2 => n6617, B1 => n4904, B2 => 
                           n6618, ZN => n1619);
   U2214 : OAI22_X1 port map( A1 => n6533, A2 => n6617, B1 => n4905, B2 => 
                           n6618, ZN => n1618);
   U2215 : OAI22_X1 port map( A1 => n6534, A2 => n6617, B1 => n4906, B2 => 
                           n6618, ZN => n1617);
   U2216 : OAI22_X1 port map( A1 => n6535, A2 => n6617, B1 => n4907, B2 => 
                           n6618, ZN => n1616);
   U2217 : OAI22_X1 port map( A1 => n6536, A2 => n6617, B1 => n4908, B2 => 
                           n6618, ZN => n1615);
   U2218 : OAI22_X1 port map( A1 => n6537, A2 => n6617, B1 => n4909, B2 => 
                           n6618, ZN => n1614);
   U2219 : OAI22_X1 port map( A1 => n6538, A2 => n6617, B1 => n4910, B2 => 
                           n6618, ZN => n1613);
   U2220 : OAI22_X1 port map( A1 => n6539, A2 => n6617, B1 => n4911, B2 => 
                           n6618, ZN => n1612);
   U2221 : OAI22_X1 port map( A1 => n6540, A2 => n6617, B1 => n4912, B2 => 
                           n6618, ZN => n1611);
   U2222 : OAI22_X1 port map( A1 => n6541, A2 => n6617, B1 => n4913, B2 => 
                           n6618, ZN => n1610);
   U2223 : OAI22_X1 port map( A1 => n6542, A2 => n6617, B1 => n4914, B2 => 
                           n6618, ZN => n1609);
   U2224 : OAI22_X1 port map( A1 => n6543, A2 => n6617, B1 => n4915, B2 => 
                           n6618, ZN => n1608);
   U2225 : OAI22_X1 port map( A1 => n6544, A2 => n6617, B1 => n4916, B2 => 
                           n6618, ZN => n1607);
   U2226 : OAI22_X1 port map( A1 => n6545, A2 => n6617, B1 => n4917, B2 => 
                           n6618, ZN => n1606);
   U2227 : OAI22_X1 port map( A1 => n6546, A2 => n6617, B1 => n4918, B2 => 
                           n6618, ZN => n1605);
   U2228 : OAI22_X1 port map( A1 => n6547, A2 => n6617, B1 => n4919, B2 => 
                           n6618, ZN => n1604);
   U2229 : OAI22_X1 port map( A1 => n6548, A2 => n6617, B1 => n4920, B2 => 
                           n6618, ZN => n1603);
   U2230 : OAI22_X1 port map( A1 => n6549, A2 => n6617, B1 => n4921, B2 => 
                           n6618, ZN => n1602);
   U2231 : OAI22_X1 port map( A1 => n6550, A2 => n6617, B1 => n4922, B2 => 
                           n6618, ZN => n1601);
   U2232 : OAI22_X1 port map( A1 => n6551, A2 => n6617, B1 => n4923, B2 => 
                           n6618, ZN => n1600);
   U2233 : OAI22_X1 port map( A1 => n6552, A2 => n6617, B1 => n4924, B2 => 
                           n6618, ZN => n1599);
   U2234 : OAI22_X1 port map( A1 => n6553, A2 => n6617, B1 => n4925, B2 => 
                           n6618, ZN => n1598);
   U2235 : OAI22_X1 port map( A1 => n6554, A2 => n6617, B1 => n4926, B2 => 
                           n6618, ZN => n1597);
   U2236 : OAI22_X1 port map( A1 => n6555, A2 => n6617, B1 => n4927, B2 => 
                           n6618, ZN => n1596);
   U2237 : OAI22_X1 port map( A1 => n6556, A2 => n6617, B1 => n4928, B2 => 
                           n6618, ZN => n1595);
   U2238 : OAI22_X1 port map( A1 => n6557, A2 => n6617, B1 => n4929, B2 => 
                           n6618, ZN => n1594);
   U2239 : OAI22_X1 port map( A1 => n6558, A2 => n6617, B1 => n4930, B2 => 
                           n6618, ZN => n1593);
   U2240 : OAI22_X1 port map( A1 => n6559, A2 => n6617, B1 => n4931, B2 => 
                           n6618, ZN => n1592);
   U2241 : OAI22_X1 port map( A1 => n6560, A2 => n6617, B1 => n4932, B2 => 
                           n6618, ZN => n1591);
   U2242 : OAI22_X1 port map( A1 => n6528, A2 => n6619, B1 => n4549, B2 => 
                           n6620, ZN => n1590);
   U2243 : OAI22_X1 port map( A1 => n6530, A2 => n6619, B1 => n4550, B2 => 
                           n6620, ZN => n1589);
   U2244 : OAI22_X1 port map( A1 => n6531, A2 => n6619, B1 => n4551, B2 => 
                           n6620, ZN => n1588);
   U2245 : OAI22_X1 port map( A1 => n6532, A2 => n6619, B1 => n4552, B2 => 
                           n6620, ZN => n1587);
   U2246 : OAI22_X1 port map( A1 => n6533, A2 => n6619, B1 => n4553, B2 => 
                           n6620, ZN => n1586);
   U2247 : OAI22_X1 port map( A1 => n6534, A2 => n6619, B1 => n4554, B2 => 
                           n6620, ZN => n1585);
   U2248 : OAI22_X1 port map( A1 => n6535, A2 => n6619, B1 => n4555, B2 => 
                           n6620, ZN => n1584);
   U2249 : OAI22_X1 port map( A1 => n6536, A2 => n6619, B1 => n4556, B2 => 
                           n6620, ZN => n1583);
   U2250 : OAI22_X1 port map( A1 => n6537, A2 => n6619, B1 => n4557, B2 => 
                           n6620, ZN => n1582);
   U2251 : OAI22_X1 port map( A1 => n6538, A2 => n6619, B1 => n4558, B2 => 
                           n6620, ZN => n1581);
   U2252 : OAI22_X1 port map( A1 => n6539, A2 => n6619, B1 => n4559, B2 => 
                           n6620, ZN => n1580);
   U2253 : OAI22_X1 port map( A1 => n6540, A2 => n6619, B1 => n4560, B2 => 
                           n6620, ZN => n1579);
   U2254 : OAI22_X1 port map( A1 => n6541, A2 => n6619, B1 => n4561, B2 => 
                           n6620, ZN => n1578);
   U2255 : OAI22_X1 port map( A1 => n6542, A2 => n6619, B1 => n4562, B2 => 
                           n6620, ZN => n1577);
   U2256 : OAI22_X1 port map( A1 => n6543, A2 => n6619, B1 => n4563, B2 => 
                           n6620, ZN => n1576);
   U2257 : OAI22_X1 port map( A1 => n6544, A2 => n6619, B1 => n4564, B2 => 
                           n6620, ZN => n1575);
   U2258 : OAI22_X1 port map( A1 => n6545, A2 => n6619, B1 => n4565, B2 => 
                           n6620, ZN => n1574);
   U2259 : OAI22_X1 port map( A1 => n6546, A2 => n6619, B1 => n4566, B2 => 
                           n6620, ZN => n1573);
   U2260 : OAI22_X1 port map( A1 => n6547, A2 => n6619, B1 => n4567, B2 => 
                           n6620, ZN => n1572);
   U2261 : OAI22_X1 port map( A1 => n6548, A2 => n6619, B1 => n4568, B2 => 
                           n6620, ZN => n1571);
   U2262 : OAI22_X1 port map( A1 => n6549, A2 => n6619, B1 => n4569, B2 => 
                           n6620, ZN => n1570);
   U2263 : OAI22_X1 port map( A1 => n6550, A2 => n6619, B1 => n4570, B2 => 
                           n6620, ZN => n1569);
   U2264 : OAI22_X1 port map( A1 => n6551, A2 => n6619, B1 => n4571, B2 => 
                           n6620, ZN => n1568);
   U2265 : OAI22_X1 port map( A1 => n6552, A2 => n6619, B1 => n4572, B2 => 
                           n6620, ZN => n1567);
   U2266 : OAI22_X1 port map( A1 => n6553, A2 => n6619, B1 => n4573, B2 => 
                           n6620, ZN => n1566);
   U2267 : OAI22_X1 port map( A1 => n6554, A2 => n6619, B1 => n4574, B2 => 
                           n6620, ZN => n1565);
   U2268 : OAI22_X1 port map( A1 => n6555, A2 => n6619, B1 => n4575, B2 => 
                           n6620, ZN => n1564);
   U2269 : OAI22_X1 port map( A1 => n6556, A2 => n6619, B1 => n4576, B2 => 
                           n6620, ZN => n1563);
   U2270 : OAI22_X1 port map( A1 => n6557, A2 => n6619, B1 => n4577, B2 => 
                           n6620, ZN => n1562);
   U2271 : OAI22_X1 port map( A1 => n6558, A2 => n6619, B1 => n4578, B2 => 
                           n6620, ZN => n1561);
   U2272 : OAI22_X1 port map( A1 => n6559, A2 => n6619, B1 => n4579, B2 => 
                           n6620, ZN => n1560);
   U2273 : OAI22_X1 port map( A1 => n6560, A2 => n6619, B1 => n4580, B2 => 
                           n6620, ZN => n1559);
   U2274 : AND3_X1 port map( A1 => n6586, A2 => n6584, A3 => ADD_WR(4), ZN => 
                           n6606);
   U2275 : INV_X1 port map( A => ADD_WR(3), ZN => n6584);
   U2276 : OAI22_X1 port map( A1 => n6528, A2 => n6621, B1 => n4581, B2 => 
                           n6622, ZN => n1558);
   U2277 : OAI22_X1 port map( A1 => n6530, A2 => n6621, B1 => n4582, B2 => 
                           n6622, ZN => n1557);
   U2278 : OAI22_X1 port map( A1 => n6531, A2 => n6621, B1 => n4583, B2 => 
                           n6622, ZN => n1556);
   U2279 : OAI22_X1 port map( A1 => n6532, A2 => n6621, B1 => n4584, B2 => 
                           n6622, ZN => n1555);
   U2280 : OAI22_X1 port map( A1 => n6533, A2 => n6621, B1 => n4585, B2 => 
                           n6622, ZN => n1554);
   U2281 : OAI22_X1 port map( A1 => n6534, A2 => n6621, B1 => n4586, B2 => 
                           n6622, ZN => n1553);
   U2282 : OAI22_X1 port map( A1 => n6535, A2 => n6621, B1 => n4587, B2 => 
                           n6622, ZN => n1552);
   U2283 : OAI22_X1 port map( A1 => n6536, A2 => n6621, B1 => n4588, B2 => 
                           n6622, ZN => n1551);
   U2284 : OAI22_X1 port map( A1 => n6537, A2 => n6621, B1 => n4589, B2 => 
                           n6622, ZN => n1550);
   U2285 : OAI22_X1 port map( A1 => n6538, A2 => n6621, B1 => n4590, B2 => 
                           n6622, ZN => n1549);
   U2286 : OAI22_X1 port map( A1 => n6539, A2 => n6621, B1 => n4591, B2 => 
                           n6622, ZN => n1548);
   U2287 : OAI22_X1 port map( A1 => n6540, A2 => n6621, B1 => n4592, B2 => 
                           n6622, ZN => n1547);
   U2288 : OAI22_X1 port map( A1 => n6541, A2 => n6621, B1 => n4593, B2 => 
                           n6622, ZN => n1546);
   U2289 : OAI22_X1 port map( A1 => n6542, A2 => n6621, B1 => n4594, B2 => 
                           n6622, ZN => n1545);
   U2290 : OAI22_X1 port map( A1 => n6543, A2 => n6621, B1 => n4595, B2 => 
                           n6622, ZN => n1544);
   U2291 : OAI22_X1 port map( A1 => n6544, A2 => n6621, B1 => n4596, B2 => 
                           n6622, ZN => n1543);
   U2292 : OAI22_X1 port map( A1 => n6545, A2 => n6621, B1 => n4597, B2 => 
                           n6622, ZN => n1542);
   U2293 : OAI22_X1 port map( A1 => n6546, A2 => n6621, B1 => n4598, B2 => 
                           n6622, ZN => n1541);
   U2294 : OAI22_X1 port map( A1 => n6547, A2 => n6621, B1 => n4599, B2 => 
                           n6622, ZN => n1540);
   U2295 : OAI22_X1 port map( A1 => n6548, A2 => n6621, B1 => n4600, B2 => 
                           n6622, ZN => n1539);
   U2296 : OAI22_X1 port map( A1 => n6549, A2 => n6621, B1 => n4601, B2 => 
                           n6622, ZN => n1538);
   U2297 : OAI22_X1 port map( A1 => n6550, A2 => n6621, B1 => n4602, B2 => 
                           n6622, ZN => n1537);
   U2298 : OAI22_X1 port map( A1 => n6551, A2 => n6621, B1 => n4603, B2 => 
                           n6622, ZN => n1536);
   U2299 : OAI22_X1 port map( A1 => n6552, A2 => n6621, B1 => n4604, B2 => 
                           n6622, ZN => n1535);
   U2300 : OAI22_X1 port map( A1 => n6553, A2 => n6621, B1 => n4605, B2 => 
                           n6622, ZN => n1534);
   U2301 : OAI22_X1 port map( A1 => n6554, A2 => n6621, B1 => n4606, B2 => 
                           n6622, ZN => n1533);
   U2302 : OAI22_X1 port map( A1 => n6555, A2 => n6621, B1 => n4607, B2 => 
                           n6622, ZN => n1532);
   U2303 : OAI22_X1 port map( A1 => n6556, A2 => n6621, B1 => n4608, B2 => 
                           n6622, ZN => n1531);
   U2304 : OAI22_X1 port map( A1 => n6557, A2 => n6621, B1 => n4609, B2 => 
                           n6622, ZN => n1530);
   U2305 : OAI22_X1 port map( A1 => n6558, A2 => n6621, B1 => n4610, B2 => 
                           n6622, ZN => n1529);
   U2306 : OAI22_X1 port map( A1 => n6559, A2 => n6621, B1 => n4611, B2 => 
                           n6622, ZN => n1528);
   U2307 : OAI22_X1 port map( A1 => n6560, A2 => n6621, B1 => n4612, B2 => 
                           n6622, ZN => n1527);
   U2308 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => ADD_WR(0),
                           ZN => n6561);
   U2309 : OAI22_X1 port map( A1 => n6528, A2 => n6624, B1 => n4323, B2 => 
                           n6625, ZN => n1526);
   U2310 : OAI22_X1 port map( A1 => n6530, A2 => n6624, B1 => n4324, B2 => 
                           n6625, ZN => n1525);
   U2311 : OAI22_X1 port map( A1 => n6531, A2 => n6624, B1 => n4325, B2 => 
                           n6625, ZN => n1524);
   U2312 : OAI22_X1 port map( A1 => n6532, A2 => n6624, B1 => n4326, B2 => 
                           n6625, ZN => n1523);
   U2313 : OAI22_X1 port map( A1 => n6533, A2 => n6624, B1 => n4327, B2 => 
                           n6625, ZN => n1522);
   U2314 : OAI22_X1 port map( A1 => n6534, A2 => n6624, B1 => n4328, B2 => 
                           n6625, ZN => n1521);
   U2315 : OAI22_X1 port map( A1 => n6535, A2 => n6624, B1 => n4329, B2 => 
                           n6625, ZN => n1520);
   U2316 : OAI22_X1 port map( A1 => n6536, A2 => n6624, B1 => n4330, B2 => 
                           n6625, ZN => n1519);
   U2317 : OAI22_X1 port map( A1 => n6537, A2 => n6624, B1 => n4331, B2 => 
                           n6625, ZN => n1518);
   U2318 : OAI22_X1 port map( A1 => n6538, A2 => n6624, B1 => n4332, B2 => 
                           n6625, ZN => n1517);
   U2319 : OAI22_X1 port map( A1 => n6539, A2 => n6624, B1 => n4333, B2 => 
                           n6625, ZN => n1516);
   U2320 : OAI22_X1 port map( A1 => n6540, A2 => n6624, B1 => n4334, B2 => 
                           n6625, ZN => n1515);
   U2321 : OAI22_X1 port map( A1 => n6541, A2 => n6624, B1 => n4335, B2 => 
                           n6625, ZN => n1514);
   U2322 : OAI22_X1 port map( A1 => n6542, A2 => n6624, B1 => n4336, B2 => 
                           n6625, ZN => n1513);
   U2323 : OAI22_X1 port map( A1 => n6543, A2 => n6624, B1 => n4337, B2 => 
                           n6625, ZN => n1512);
   U2324 : OAI22_X1 port map( A1 => n6544, A2 => n6624, B1 => n4338, B2 => 
                           n6625, ZN => n1511);
   U2325 : OAI22_X1 port map( A1 => n6545, A2 => n6624, B1 => n4339, B2 => 
                           n6625, ZN => n1510);
   U2326 : OAI22_X1 port map( A1 => n6546, A2 => n6624, B1 => n4340, B2 => 
                           n6625, ZN => n1509);
   U2327 : OAI22_X1 port map( A1 => n6547, A2 => n6624, B1 => n4341, B2 => 
                           n6625, ZN => n1508);
   U2328 : OAI22_X1 port map( A1 => n6548, A2 => n6624, B1 => n4342, B2 => 
                           n6625, ZN => n1507);
   U2329 : OAI22_X1 port map( A1 => n6549, A2 => n6624, B1 => n4343, B2 => 
                           n6625, ZN => n1506);
   U2330 : OAI22_X1 port map( A1 => n6550, A2 => n6624, B1 => n4344, B2 => 
                           n6625, ZN => n1505);
   U2331 : OAI22_X1 port map( A1 => n6551, A2 => n6624, B1 => n4345, B2 => 
                           n6625, ZN => n1504);
   U2332 : OAI22_X1 port map( A1 => n6552, A2 => n6624, B1 => n4346, B2 => 
                           n6625, ZN => n1503);
   U2333 : OAI22_X1 port map( A1 => n6553, A2 => n6624, B1 => n4347, B2 => 
                           n6625, ZN => n1502);
   U2334 : OAI22_X1 port map( A1 => n6554, A2 => n6624, B1 => n4348, B2 => 
                           n6625, ZN => n1501);
   U2335 : OAI22_X1 port map( A1 => n6555, A2 => n6624, B1 => n4349, B2 => 
                           n6625, ZN => n1500);
   U2336 : OAI22_X1 port map( A1 => n6556, A2 => n6624, B1 => n4350, B2 => 
                           n6625, ZN => n1499);
   U2337 : OAI22_X1 port map( A1 => n6557, A2 => n6624, B1 => n4351, B2 => 
                           n6625, ZN => n1498);
   U2338 : OAI22_X1 port map( A1 => n6558, A2 => n6624, B1 => n4352, B2 => 
                           n6625, ZN => n1497);
   U2339 : OAI22_X1 port map( A1 => n6559, A2 => n6624, B1 => n4353, B2 => 
                           n6625, ZN => n1496);
   U2340 : OAI22_X1 port map( A1 => n6560, A2 => n6624, B1 => n4354, B2 => 
                           n6625, ZN => n1495);
   U2341 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n6626, ZN 
                           => n6565);
   U2342 : OAI22_X1 port map( A1 => n6528, A2 => n6627, B1 => n4933, B2 => 
                           n6628, ZN => n1494);
   U2343 : OAI22_X1 port map( A1 => n6530, A2 => n6627, B1 => n4934, B2 => 
                           n6628, ZN => n1493);
   U2344 : OAI22_X1 port map( A1 => n6531, A2 => n6627, B1 => n4935, B2 => 
                           n6628, ZN => n1492);
   U2345 : OAI22_X1 port map( A1 => n6532, A2 => n6627, B1 => n4936, B2 => 
                           n6628, ZN => n1491);
   U2346 : OAI22_X1 port map( A1 => n6533, A2 => n6627, B1 => n4937, B2 => 
                           n6628, ZN => n1490);
   U2347 : OAI22_X1 port map( A1 => n6534, A2 => n6627, B1 => n4938, B2 => 
                           n6628, ZN => n1489);
   U2348 : OAI22_X1 port map( A1 => n6535, A2 => n6627, B1 => n4939, B2 => 
                           n6628, ZN => n1488);
   U2349 : OAI22_X1 port map( A1 => n6536, A2 => n6627, B1 => n4940, B2 => 
                           n6628, ZN => n1487);
   U2350 : OAI22_X1 port map( A1 => n6537, A2 => n6627, B1 => n4941, B2 => 
                           n6628, ZN => n1486);
   U2351 : OAI22_X1 port map( A1 => n6538, A2 => n6627, B1 => n4942, B2 => 
                           n6628, ZN => n1485);
   U2352 : OAI22_X1 port map( A1 => n6539, A2 => n6627, B1 => n4943, B2 => 
                           n6628, ZN => n1484);
   U2353 : OAI22_X1 port map( A1 => n6540, A2 => n6627, B1 => n4944, B2 => 
                           n6628, ZN => n1483);
   U2354 : OAI22_X1 port map( A1 => n6541, A2 => n6627, B1 => n4945, B2 => 
                           n6628, ZN => n1482);
   U2355 : OAI22_X1 port map( A1 => n6542, A2 => n6627, B1 => n4946, B2 => 
                           n6628, ZN => n1481);
   U2356 : OAI22_X1 port map( A1 => n6543, A2 => n6627, B1 => n4947, B2 => 
                           n6628, ZN => n1480);
   U2357 : OAI22_X1 port map( A1 => n6544, A2 => n6627, B1 => n4948, B2 => 
                           n6628, ZN => n1479);
   U2358 : OAI22_X1 port map( A1 => n6545, A2 => n6627, B1 => n4949, B2 => 
                           n6628, ZN => n1478);
   U2359 : OAI22_X1 port map( A1 => n6546, A2 => n6627, B1 => n4950, B2 => 
                           n6628, ZN => n1477);
   U2360 : OAI22_X1 port map( A1 => n6547, A2 => n6627, B1 => n4951, B2 => 
                           n6628, ZN => n1476);
   U2361 : OAI22_X1 port map( A1 => n6548, A2 => n6627, B1 => n4952, B2 => 
                           n6628, ZN => n1475);
   U2362 : OAI22_X1 port map( A1 => n6549, A2 => n6627, B1 => n4953, B2 => 
                           n6628, ZN => n1474);
   U2363 : OAI22_X1 port map( A1 => n6550, A2 => n6627, B1 => n4954, B2 => 
                           n6628, ZN => n1473);
   U2364 : OAI22_X1 port map( A1 => n6551, A2 => n6627, B1 => n4955, B2 => 
                           n6628, ZN => n1472);
   U2365 : OAI22_X1 port map( A1 => n6552, A2 => n6627, B1 => n4956, B2 => 
                           n6628, ZN => n1471);
   U2366 : OAI22_X1 port map( A1 => n6553, A2 => n6627, B1 => n4957, B2 => 
                           n6628, ZN => n1470);
   U2367 : OAI22_X1 port map( A1 => n6554, A2 => n6627, B1 => n4958, B2 => 
                           n6628, ZN => n1469);
   U2368 : OAI22_X1 port map( A1 => n6555, A2 => n6627, B1 => n4959, B2 => 
                           n6628, ZN => n1468);
   U2369 : OAI22_X1 port map( A1 => n6556, A2 => n6627, B1 => n4960, B2 => 
                           n6628, ZN => n1467);
   U2370 : OAI22_X1 port map( A1 => n6557, A2 => n6627, B1 => n4961, B2 => 
                           n6628, ZN => n1466);
   U2371 : OAI22_X1 port map( A1 => n6558, A2 => n6627, B1 => n4962, B2 => 
                           n6628, ZN => n1465);
   U2372 : OAI22_X1 port map( A1 => n6559, A2 => n6627, B1 => n4963, B2 => 
                           n6628, ZN => n1464);
   U2373 : OAI22_X1 port map( A1 => n6560, A2 => n6627, B1 => n4964, B2 => 
                           n6628, ZN => n1463);
   U2374 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n6629, ZN 
                           => n6568);
   U2375 : OAI22_X1 port map( A1 => n6528, A2 => n6630, B1 => n4355, B2 => 
                           n6631, ZN => n1462);
   U2376 : OAI22_X1 port map( A1 => n6530, A2 => n6630, B1 => n4356, B2 => 
                           n6631, ZN => n1461);
   U2377 : OAI22_X1 port map( A1 => n6531, A2 => n6630, B1 => n4357, B2 => 
                           n6631, ZN => n1460);
   U2378 : OAI22_X1 port map( A1 => n6532, A2 => n6630, B1 => n4358, B2 => 
                           n6631, ZN => n1459);
   U2379 : OAI22_X1 port map( A1 => n6533, A2 => n6630, B1 => n4359, B2 => 
                           n6631, ZN => n1458);
   U2380 : OAI22_X1 port map( A1 => n6534, A2 => n6630, B1 => n4360, B2 => 
                           n6631, ZN => n1457);
   U2381 : OAI22_X1 port map( A1 => n6535, A2 => n6630, B1 => n4361, B2 => 
                           n6631, ZN => n1456);
   U2382 : OAI22_X1 port map( A1 => n6536, A2 => n6630, B1 => n4362, B2 => 
                           n6631, ZN => n1455);
   U2383 : OAI22_X1 port map( A1 => n6537, A2 => n6630, B1 => n4363, B2 => 
                           n6631, ZN => n1454);
   U2384 : OAI22_X1 port map( A1 => n6538, A2 => n6630, B1 => n4364, B2 => 
                           n6631, ZN => n1453);
   U2385 : OAI22_X1 port map( A1 => n6539, A2 => n6630, B1 => n4365, B2 => 
                           n6631, ZN => n1452);
   U2386 : OAI22_X1 port map( A1 => n6540, A2 => n6630, B1 => n4366, B2 => 
                           n6631, ZN => n1451);
   U2387 : OAI22_X1 port map( A1 => n6541, A2 => n6630, B1 => n4367, B2 => 
                           n6631, ZN => n1450);
   U2388 : OAI22_X1 port map( A1 => n6542, A2 => n6630, B1 => n4368, B2 => 
                           n6631, ZN => n1449);
   U2389 : OAI22_X1 port map( A1 => n6543, A2 => n6630, B1 => n4369, B2 => 
                           n6631, ZN => n1448);
   U2390 : OAI22_X1 port map( A1 => n6544, A2 => n6630, B1 => n4370, B2 => 
                           n6631, ZN => n1447);
   U2391 : OAI22_X1 port map( A1 => n6545, A2 => n6630, B1 => n4371, B2 => 
                           n6631, ZN => n1446);
   U2392 : OAI22_X1 port map( A1 => n6546, A2 => n6630, B1 => n4372, B2 => 
                           n6631, ZN => n1445);
   U2393 : OAI22_X1 port map( A1 => n6547, A2 => n6630, B1 => n4373, B2 => 
                           n6631, ZN => n1444);
   U2394 : OAI22_X1 port map( A1 => n6548, A2 => n6630, B1 => n4374, B2 => 
                           n6631, ZN => n1443);
   U2395 : OAI22_X1 port map( A1 => n6549, A2 => n6630, B1 => n4375, B2 => 
                           n6631, ZN => n1442);
   U2396 : OAI22_X1 port map( A1 => n6550, A2 => n6630, B1 => n4376, B2 => 
                           n6631, ZN => n1441);
   U2397 : OAI22_X1 port map( A1 => n6551, A2 => n6630, B1 => n4377, B2 => 
                           n6631, ZN => n1440);
   U2398 : OAI22_X1 port map( A1 => n6552, A2 => n6630, B1 => n4378, B2 => 
                           n6631, ZN => n1439);
   U2399 : OAI22_X1 port map( A1 => n6553, A2 => n6630, B1 => n4379, B2 => 
                           n6631, ZN => n1438);
   U2400 : OAI22_X1 port map( A1 => n6554, A2 => n6630, B1 => n4380, B2 => 
                           n6631, ZN => n1437);
   U2401 : OAI22_X1 port map( A1 => n6555, A2 => n6630, B1 => n4381, B2 => 
                           n6631, ZN => n1436);
   U2402 : OAI22_X1 port map( A1 => n6556, A2 => n6630, B1 => n4382, B2 => 
                           n6631, ZN => n1435);
   U2403 : OAI22_X1 port map( A1 => n6557, A2 => n6630, B1 => n4383, B2 => 
                           n6631, ZN => n1434);
   U2404 : OAI22_X1 port map( A1 => n6558, A2 => n6630, B1 => n4384, B2 => 
                           n6631, ZN => n1433);
   U2405 : OAI22_X1 port map( A1 => n6559, A2 => n6630, B1 => n4385, B2 => 
                           n6631, ZN => n1432);
   U2406 : OAI22_X1 port map( A1 => n6560, A2 => n6630, B1 => n4386, B2 => 
                           n6631, ZN => n1431);
   U2407 : NOR3_X1 port map( A1 => n6626, A2 => ADD_WR(2), A3 => n6629, ZN => 
                           n6571);
   U2408 : OAI22_X1 port map( A1 => n6528, A2 => n6632, B1 => n4613, B2 => 
                           n6633, ZN => n1430);
   U2409 : OAI22_X1 port map( A1 => n6530, A2 => n6632, B1 => n4614, B2 => 
                           n6633, ZN => n1429);
   U2410 : OAI22_X1 port map( A1 => n6531, A2 => n6632, B1 => n4615, B2 => 
                           n6633, ZN => n1428);
   U2411 : OAI22_X1 port map( A1 => n6532, A2 => n6632, B1 => n4616, B2 => 
                           n6633, ZN => n1427);
   U2412 : OAI22_X1 port map( A1 => n6533, A2 => n6632, B1 => n4617, B2 => 
                           n6633, ZN => n1426);
   U2413 : OAI22_X1 port map( A1 => n6534, A2 => n6632, B1 => n4618, B2 => 
                           n6633, ZN => n1425);
   U2414 : OAI22_X1 port map( A1 => n6535, A2 => n6632, B1 => n4619, B2 => 
                           n6633, ZN => n1424);
   U2415 : OAI22_X1 port map( A1 => n6536, A2 => n6632, B1 => n4620, B2 => 
                           n6633, ZN => n1423);
   U2416 : OAI22_X1 port map( A1 => n6537, A2 => n6632, B1 => n4621, B2 => 
                           n6633, ZN => n1422);
   U2417 : OAI22_X1 port map( A1 => n6538, A2 => n6632, B1 => n4622, B2 => 
                           n6633, ZN => n1421);
   U2418 : OAI22_X1 port map( A1 => n6539, A2 => n6632, B1 => n4623, B2 => 
                           n6633, ZN => n1420);
   U2419 : OAI22_X1 port map( A1 => n6540, A2 => n6632, B1 => n4624, B2 => 
                           n6633, ZN => n1419);
   U2420 : OAI22_X1 port map( A1 => n6541, A2 => n6632, B1 => n4625, B2 => 
                           n6633, ZN => n1418);
   U2421 : OAI22_X1 port map( A1 => n6542, A2 => n6632, B1 => n4626, B2 => 
                           n6633, ZN => n1417);
   U2422 : OAI22_X1 port map( A1 => n6543, A2 => n6632, B1 => n4627, B2 => 
                           n6633, ZN => n1416);
   U2423 : OAI22_X1 port map( A1 => n6544, A2 => n6632, B1 => n4628, B2 => 
                           n6633, ZN => n1415);
   U2424 : OAI22_X1 port map( A1 => n6545, A2 => n6632, B1 => n4629, B2 => 
                           n6633, ZN => n1414);
   U2425 : OAI22_X1 port map( A1 => n6546, A2 => n6632, B1 => n4630, B2 => 
                           n6633, ZN => n1413);
   U2426 : OAI22_X1 port map( A1 => n6547, A2 => n6632, B1 => n4631, B2 => 
                           n6633, ZN => n1412);
   U2427 : OAI22_X1 port map( A1 => n6548, A2 => n6632, B1 => n4632, B2 => 
                           n6633, ZN => n1411);
   U2428 : OAI22_X1 port map( A1 => n6549, A2 => n6632, B1 => n4633, B2 => 
                           n6633, ZN => n1410);
   U2429 : OAI22_X1 port map( A1 => n6550, A2 => n6632, B1 => n4634, B2 => 
                           n6633, ZN => n1409);
   U2430 : OAI22_X1 port map( A1 => n6551, A2 => n6632, B1 => n4635, B2 => 
                           n6633, ZN => n1408);
   U2431 : OAI22_X1 port map( A1 => n6552, A2 => n6632, B1 => n4636, B2 => 
                           n6633, ZN => n1407);
   U2432 : OAI22_X1 port map( A1 => n6553, A2 => n6632, B1 => n4637, B2 => 
                           n6633, ZN => n1406);
   U2433 : OAI22_X1 port map( A1 => n6554, A2 => n6632, B1 => n4638, B2 => 
                           n6633, ZN => n1405);
   U2434 : OAI22_X1 port map( A1 => n6555, A2 => n6632, B1 => n4639, B2 => 
                           n6633, ZN => n1404);
   U2435 : OAI22_X1 port map( A1 => n6556, A2 => n6632, B1 => n4640, B2 => 
                           n6633, ZN => n1403);
   U2436 : OAI22_X1 port map( A1 => n6557, A2 => n6632, B1 => n4641, B2 => 
                           n6633, ZN => n1402);
   U2437 : OAI22_X1 port map( A1 => n6558, A2 => n6632, B1 => n4642, B2 => 
                           n6633, ZN => n1401);
   U2438 : OAI22_X1 port map( A1 => n6559, A2 => n6632, B1 => n4643, B2 => 
                           n6633, ZN => n1400);
   U2439 : OAI22_X1 port map( A1 => n6560, A2 => n6632, B1 => n4644, B2 => 
                           n6633, ZN => n1399);
   U2440 : AND3_X1 port map( A1 => n6626, A2 => n6629, A3 => ADD_WR(2), ZN => 
                           n6574);
   U2441 : OAI22_X1 port map( A1 => n6528, A2 => n6634, B1 => n4387, B2 => 
                           n6635, ZN => n1398);
   U2442 : OAI22_X1 port map( A1 => n6530, A2 => n6634, B1 => n4388, B2 => 
                           n6635, ZN => n1397);
   U2443 : OAI22_X1 port map( A1 => n6531, A2 => n6634, B1 => n4389, B2 => 
                           n6635, ZN => n1396);
   U2444 : OAI22_X1 port map( A1 => n6532, A2 => n6634, B1 => n4390, B2 => 
                           n6635, ZN => n1395);
   U2445 : OAI22_X1 port map( A1 => n6533, A2 => n6634, B1 => n4391, B2 => 
                           n6635, ZN => n1394);
   U2446 : OAI22_X1 port map( A1 => n6534, A2 => n6634, B1 => n4392, B2 => 
                           n6635, ZN => n1393);
   U2447 : OAI22_X1 port map( A1 => n6535, A2 => n6634, B1 => n4393, B2 => 
                           n6635, ZN => n1392);
   U2448 : OAI22_X1 port map( A1 => n6536, A2 => n6634, B1 => n4394, B2 => 
                           n6635, ZN => n1391);
   U2449 : OAI22_X1 port map( A1 => n6537, A2 => n6634, B1 => n4395, B2 => 
                           n6635, ZN => n1390);
   U2450 : OAI22_X1 port map( A1 => n6538, A2 => n6634, B1 => n4396, B2 => 
                           n6635, ZN => n1389);
   U2451 : OAI22_X1 port map( A1 => n6539, A2 => n6634, B1 => n4397, B2 => 
                           n6635, ZN => n1388);
   U2452 : OAI22_X1 port map( A1 => n6540, A2 => n6634, B1 => n4398, B2 => 
                           n6635, ZN => n1387);
   U2453 : OAI22_X1 port map( A1 => n6541, A2 => n6634, B1 => n4399, B2 => 
                           n6635, ZN => n1386);
   U2454 : OAI22_X1 port map( A1 => n6542, A2 => n6634, B1 => n4400, B2 => 
                           n6635, ZN => n1385);
   U2455 : OAI22_X1 port map( A1 => n6543, A2 => n6634, B1 => n4401, B2 => 
                           n6635, ZN => n1384);
   U2456 : OAI22_X1 port map( A1 => n6544, A2 => n6634, B1 => n4402, B2 => 
                           n6635, ZN => n1383);
   U2457 : OAI22_X1 port map( A1 => n6545, A2 => n6634, B1 => n4403, B2 => 
                           n6635, ZN => n1382);
   U2458 : OAI22_X1 port map( A1 => n6546, A2 => n6634, B1 => n4404, B2 => 
                           n6635, ZN => n1381);
   U2459 : OAI22_X1 port map( A1 => n6547, A2 => n6634, B1 => n4405, B2 => 
                           n6635, ZN => n1380);
   U2460 : OAI22_X1 port map( A1 => n6548, A2 => n6634, B1 => n4406, B2 => 
                           n6635, ZN => n1379);
   U2461 : OAI22_X1 port map( A1 => n6549, A2 => n6634, B1 => n4407, B2 => 
                           n6635, ZN => n1378);
   U2462 : OAI22_X1 port map( A1 => n6550, A2 => n6634, B1 => n4408, B2 => 
                           n6635, ZN => n1377);
   U2463 : OAI22_X1 port map( A1 => n6551, A2 => n6634, B1 => n4409, B2 => 
                           n6635, ZN => n1376);
   U2464 : OAI22_X1 port map( A1 => n6552, A2 => n6634, B1 => n4410, B2 => 
                           n6635, ZN => n1375);
   U2465 : OAI22_X1 port map( A1 => n6553, A2 => n6634, B1 => n4411, B2 => 
                           n6635, ZN => n1374);
   U2466 : OAI22_X1 port map( A1 => n6554, A2 => n6634, B1 => n4412, B2 => 
                           n6635, ZN => n1373);
   U2467 : OAI22_X1 port map( A1 => n6555, A2 => n6634, B1 => n4413, B2 => 
                           n6635, ZN => n1372);
   U2468 : OAI22_X1 port map( A1 => n6556, A2 => n6634, B1 => n4414, B2 => 
                           n6635, ZN => n1371);
   U2469 : OAI22_X1 port map( A1 => n6557, A2 => n6634, B1 => n4415, B2 => 
                           n6635, ZN => n1370);
   U2470 : OAI22_X1 port map( A1 => n6558, A2 => n6634, B1 => n4416, B2 => 
                           n6635, ZN => n1369);
   U2471 : OAI22_X1 port map( A1 => n6559, A2 => n6634, B1 => n4417, B2 => 
                           n6635, ZN => n1368);
   U2472 : OAI22_X1 port map( A1 => n6560, A2 => n6634, B1 => n4418, B2 => 
                           n6635, ZN => n1367);
   U2473 : AND3_X1 port map( A1 => ADD_WR(0), A2 => n6629, A3 => ADD_WR(2), ZN 
                           => n6577);
   U2474 : INV_X1 port map( A => ADD_WR(1), ZN => n6629);
   U2475 : OAI22_X1 port map( A1 => n6528, A2 => n6636, B1 => n5157, B2 => 
                           n6637, ZN => n1366);
   U2476 : OAI22_X1 port map( A1 => n6530, A2 => n6636, B1 => n5158, B2 => 
                           n6637, ZN => n1365);
   U2477 : OAI22_X1 port map( A1 => n6531, A2 => n6636, B1 => n5159, B2 => 
                           n6637, ZN => n1364);
   U2478 : OAI22_X1 port map( A1 => n6532, A2 => n6636, B1 => n5160, B2 => 
                           n6637, ZN => n1363);
   U2479 : OAI22_X1 port map( A1 => n6533, A2 => n6636, B1 => n5161, B2 => 
                           n6637, ZN => n1362);
   U2480 : OAI22_X1 port map( A1 => n6534, A2 => n6636, B1 => n5162, B2 => 
                           n6637, ZN => n1361);
   U2481 : OAI22_X1 port map( A1 => n6535, A2 => n6636, B1 => n5163, B2 => 
                           n6637, ZN => n1360);
   U2482 : OAI22_X1 port map( A1 => n6536, A2 => n6636, B1 => n5164, B2 => 
                           n6637, ZN => n1359);
   U2483 : OAI22_X1 port map( A1 => n6537, A2 => n6636, B1 => n5165, B2 => 
                           n6637, ZN => n1358);
   U2484 : OAI22_X1 port map( A1 => n6538, A2 => n6636, B1 => n5166, B2 => 
                           n6637, ZN => n1357);
   U2485 : OAI22_X1 port map( A1 => n6539, A2 => n6636, B1 => n5167, B2 => 
                           n6637, ZN => n1356);
   U2486 : OAI22_X1 port map( A1 => n6540, A2 => n6636, B1 => n5168, B2 => 
                           n6637, ZN => n1355);
   U2487 : OAI22_X1 port map( A1 => n6541, A2 => n6636, B1 => n5169, B2 => 
                           n6637, ZN => n1354);
   U2488 : OAI22_X1 port map( A1 => n6542, A2 => n6636, B1 => n5170, B2 => 
                           n6637, ZN => n1353);
   U2489 : OAI22_X1 port map( A1 => n6543, A2 => n6636, B1 => n5171, B2 => 
                           n6637, ZN => n1352);
   U2490 : OAI22_X1 port map( A1 => n6544, A2 => n6636, B1 => n5172, B2 => 
                           n6637, ZN => n1351);
   U2491 : OAI22_X1 port map( A1 => n6545, A2 => n6636, B1 => n5173, B2 => 
                           n6637, ZN => n1350);
   U2492 : OAI22_X1 port map( A1 => n6546, A2 => n6636, B1 => n5174, B2 => 
                           n6637, ZN => n1349);
   U2493 : OAI22_X1 port map( A1 => n6547, A2 => n6636, B1 => n5175, B2 => 
                           n6637, ZN => n1348);
   U2494 : OAI22_X1 port map( A1 => n6548, A2 => n6636, B1 => n5176, B2 => 
                           n6637, ZN => n1347);
   U2495 : OAI22_X1 port map( A1 => n6549, A2 => n6636, B1 => n5177, B2 => 
                           n6637, ZN => n1346);
   U2496 : OAI22_X1 port map( A1 => n6550, A2 => n6636, B1 => n5178, B2 => 
                           n6637, ZN => n1345);
   U2497 : OAI22_X1 port map( A1 => n6551, A2 => n6636, B1 => n5179, B2 => 
                           n6637, ZN => n1344);
   U2498 : OAI22_X1 port map( A1 => n6552, A2 => n6636, B1 => n5180, B2 => 
                           n6637, ZN => n1343);
   U2499 : OAI22_X1 port map( A1 => n6553, A2 => n6636, B1 => n5181, B2 => 
                           n6637, ZN => n1342);
   U2500 : OAI22_X1 port map( A1 => n6554, A2 => n6636, B1 => n5182, B2 => 
                           n6637, ZN => n1341);
   U2501 : OAI22_X1 port map( A1 => n6555, A2 => n6636, B1 => n5183, B2 => 
                           n6637, ZN => n1340);
   U2502 : OAI22_X1 port map( A1 => n6556, A2 => n6636, B1 => n5184, B2 => 
                           n6637, ZN => n1339);
   U2503 : OAI22_X1 port map( A1 => n6557, A2 => n6636, B1 => n5185, B2 => 
                           n6637, ZN => n1338);
   U2504 : OAI22_X1 port map( A1 => n6558, A2 => n6636, B1 => n5186, B2 => 
                           n6637, ZN => n1337);
   U2505 : OAI22_X1 port map( A1 => n6559, A2 => n6636, B1 => n5187, B2 => 
                           n6637, ZN => n1336);
   U2506 : OAI22_X1 port map( A1 => n6560, A2 => n6636, B1 => n5188, B2 => 
                           n6637, ZN => n1335);
   U2507 : AND3_X1 port map( A1 => ADD_WR(1), A2 => n6626, A3 => ADD_WR(2), ZN 
                           => n6580);
   U2508 : INV_X1 port map( A => ADD_WR(0), ZN => n6626);
   U2509 : OAI22_X1 port map( A1 => n6528, A2 => n6638, B1 => n4645, B2 => 
                           n6639, ZN => n1334);
   U2510 : OAI22_X1 port map( A1 => n6530, A2 => n6638, B1 => n4646, B2 => 
                           n6639, ZN => n1333);
   U2511 : OAI22_X1 port map( A1 => n6531, A2 => n6638, B1 => n4647, B2 => 
                           n6639, ZN => n1332);
   U2512 : OAI22_X1 port map( A1 => n6532, A2 => n6638, B1 => n4648, B2 => 
                           n6639, ZN => n1331);
   U2513 : OAI22_X1 port map( A1 => n6533, A2 => n6638, B1 => n4649, B2 => 
                           n6639, ZN => n1330);
   U2514 : OAI22_X1 port map( A1 => n6534, A2 => n6638, B1 => n4650, B2 => 
                           n6639, ZN => n1329);
   U2515 : OAI22_X1 port map( A1 => n6535, A2 => n6638, B1 => n4651, B2 => 
                           n6639, ZN => n1328);
   U2516 : OAI22_X1 port map( A1 => n6536, A2 => n6638, B1 => n4652, B2 => 
                           n6639, ZN => n1327);
   U2517 : OAI22_X1 port map( A1 => n6537, A2 => n6638, B1 => n4653, B2 => 
                           n6639, ZN => n1326);
   U2518 : OAI22_X1 port map( A1 => n6538, A2 => n6638, B1 => n4654, B2 => 
                           n6639, ZN => n1325);
   U2519 : OAI22_X1 port map( A1 => n6539, A2 => n6638, B1 => n4655, B2 => 
                           n6639, ZN => n1324);
   U2520 : OAI22_X1 port map( A1 => n6540, A2 => n6638, B1 => n4656, B2 => 
                           n6639, ZN => n1323);
   U2521 : OAI22_X1 port map( A1 => n6541, A2 => n6638, B1 => n4657, B2 => 
                           n6639, ZN => n1322);
   U2522 : OAI22_X1 port map( A1 => n6542, A2 => n6638, B1 => n4658, B2 => 
                           n6639, ZN => n1321);
   U2523 : OAI22_X1 port map( A1 => n6543, A2 => n6638, B1 => n4659, B2 => 
                           n6639, ZN => n1320);
   U2524 : OAI22_X1 port map( A1 => n6544, A2 => n6638, B1 => n4660, B2 => 
                           n6639, ZN => n1319);
   U2525 : OAI22_X1 port map( A1 => n6545, A2 => n6638, B1 => n4661, B2 => 
                           n6639, ZN => n1318);
   U2526 : OAI22_X1 port map( A1 => n6546, A2 => n6638, B1 => n4662, B2 => 
                           n6639, ZN => n1317);
   U2527 : OAI22_X1 port map( A1 => n6547, A2 => n6638, B1 => n4663, B2 => 
                           n6639, ZN => n1316);
   U2528 : OAI22_X1 port map( A1 => n6548, A2 => n6638, B1 => n4664, B2 => 
                           n6639, ZN => n1315);
   U2529 : OAI22_X1 port map( A1 => n6549, A2 => n6638, B1 => n4665, B2 => 
                           n6639, ZN => n1314);
   U2530 : OAI22_X1 port map( A1 => n6550, A2 => n6638, B1 => n4666, B2 => 
                           n6639, ZN => n1313);
   U2531 : OAI22_X1 port map( A1 => n6551, A2 => n6638, B1 => n4667, B2 => 
                           n6639, ZN => n1312);
   U2532 : OAI22_X1 port map( A1 => n6552, A2 => n6638, B1 => n4668, B2 => 
                           n6639, ZN => n1311);
   U2533 : OAI22_X1 port map( A1 => n6553, A2 => n6638, B1 => n4669, B2 => 
                           n6639, ZN => n1310);
   U2534 : OAI22_X1 port map( A1 => n6554, A2 => n6638, B1 => n4670, B2 => 
                           n6639, ZN => n1309);
   U2535 : OAI22_X1 port map( A1 => n6555, A2 => n6638, B1 => n4671, B2 => 
                           n6639, ZN => n1308);
   U2536 : OAI22_X1 port map( A1 => n6556, A2 => n6638, B1 => n4672, B2 => 
                           n6639, ZN => n1307);
   U2537 : OAI22_X1 port map( A1 => n6557, A2 => n6638, B1 => n4673, B2 => 
                           n6639, ZN => n1306);
   U2538 : OAI22_X1 port map( A1 => n6558, A2 => n6638, B1 => n4674, B2 => 
                           n6639, ZN => n1305);
   U2539 : OAI22_X1 port map( A1 => n6559, A2 => n6638, B1 => n4675, B2 => 
                           n6639, ZN => n1304);
   U2540 : OAI22_X1 port map( A1 => n6560, A2 => n6638, B1 => n4676, B2 => 
                           n6639, ZN => n1303);
   U2541 : AND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2),
                           ZN => n6583);
   U2542 : AND3_X1 port map( A1 => ADD_WR(3), A2 => n6586, A3 => ADD_WR(4), ZN 
                           => n6623);
   U2543 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n6586);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity SIGN_EXT_bits16 is

   port( inputt : in std_logic_vector (15 downto 0);  outputt : out 
         std_logic_vector (31 downto 0));

end SIGN_EXT_bits16;

architecture SYN_BEHAVIORAL of SIGN_EXT_bits16 is

begin
   outputt <= ( inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), 
      inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), 
      inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), inputt(15), 
      inputt(14), inputt(13), inputt(12), inputt(11), inputt(10), inputt(9), 
      inputt(8), inputt(7), inputt(6), inputt(5), inputt(4), inputt(3), 
      inputt(2), inputt(1), inputt(0) );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity RCA_NBITS32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end RCA_NBITS32;

architecture SYN_BEHAVIORAL of RCA_NBITS32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346 : std_logic;

begin
   
   U2 : INV_X1 port map( A => n175, ZN => Co);
   U3 : AOI22_X1 port map( A1 => n176, A2 => A(31), B1 => n177, B2 => B(31), ZN
                           => n175);
   U4 : OR2_X1 port map( A1 => A(31), A2 => n176, ZN => n177);
   U5 : XOR2_X1 port map( A => n178, B => n179, Z => S(9));
   U6 : XOR2_X1 port map( A => n180, B => A(9), Z => n179);
   U7 : XNOR2_X1 port map( A => B(9), B => Ci, ZN => n178);
   U8 : XOR2_X1 port map( A => n181, B => n182, Z => S(8));
   U9 : XOR2_X1 port map( A => Ci, B => B(8), Z => n182);
   U10 : XOR2_X1 port map( A => A(8), B => n183, Z => n181);
   U11 : XOR2_X1 port map( A => n184, B => n185, Z => S(7));
   U12 : XOR2_X1 port map( A => n186, B => A(7), Z => n185);
   U13 : XNOR2_X1 port map( A => B(7), B => Ci, ZN => n184);
   U14 : XOR2_X1 port map( A => n187, B => n188, Z => S(6));
   U15 : XOR2_X1 port map( A => Ci, B => B(6), Z => n188);
   U16 : XOR2_X1 port map( A => A(6), B => n189, Z => n187);
   U17 : XOR2_X1 port map( A => n190, B => n191, Z => S(5));
   U18 : XNOR2_X1 port map( A => n192, B => A(5), ZN => n191);
   U19 : XNOR2_X1 port map( A => B(5), B => Ci, ZN => n190);
   U20 : XOR2_X1 port map( A => n193, B => n194, Z => S(4));
   U21 : XOR2_X1 port map( A => n195, B => A(4), Z => n194);
   U22 : XNOR2_X1 port map( A => B(4), B => Ci, ZN => n193);
   U23 : XOR2_X1 port map( A => n196, B => n197, Z => S(3));
   U24 : XOR2_X1 port map( A => n198, B => A(3), Z => n197);
   U25 : XNOR2_X1 port map( A => B(3), B => Ci, ZN => n196);
   U26 : XOR2_X1 port map( A => n199, B => n200, Z => S(31));
   U27 : XOR2_X1 port map( A => Ci, B => B(31), Z => n200);
   U28 : XOR2_X1 port map( A => n176, B => A(31), Z => n199);
   U29 : INV_X1 port map( A => n201, ZN => n176);
   U30 : AOI22_X1 port map( A1 => n202, A2 => A(30), B1 => n203, B2 => B(30), 
                           ZN => n201);
   U31 : OR2_X1 port map( A1 => n202, A2 => A(30), ZN => n203);
   U32 : XOR2_X1 port map( A => n204, B => n205, Z => S(30));
   U33 : XOR2_X1 port map( A => A(30), B => n202, Z => n205);
   U34 : AOI21_X1 port map( B1 => n206, B2 => n207, A => n208, ZN => n202);
   U35 : AOI21_X1 port map( B1 => n209, B2 => A(29), A => B(29), ZN => n208);
   U36 : INV_X1 port map( A => n209, ZN => n207);
   U37 : INV_X1 port map( A => A(29), ZN => n206);
   U38 : XOR2_X1 port map( A => Ci, B => B(30), Z => n204);
   U39 : XOR2_X1 port map( A => n210, B => n211, Z => S(2));
   U40 : XOR2_X1 port map( A => n212, B => A(2), Z => n211);
   U41 : XNOR2_X1 port map( A => B(2), B => Ci, ZN => n210);
   U42 : XOR2_X1 port map( A => n213, B => n214, Z => S(29));
   U43 : XOR2_X1 port map( A => Ci, B => B(29), Z => n214);
   U44 : XOR2_X1 port map( A => n209, B => A(29), Z => n213);
   U45 : OAI21_X1 port map( B1 => n215, B2 => n216, A => n217, ZN => n209);
   U46 : OAI21_X1 port map( B1 => A(28), B2 => n218, A => B(28), ZN => n217);
   U47 : INV_X1 port map( A => A(28), ZN => n216);
   U48 : INV_X1 port map( A => n218, ZN => n215);
   U49 : XOR2_X1 port map( A => n219, B => n220, Z => S(28));
   U50 : XOR2_X1 port map( A => Ci, B => B(28), Z => n220);
   U51 : XOR2_X1 port map( A => n218, B => A(28), Z => n219);
   U52 : OAI21_X1 port map( B1 => n221, B2 => n222, A => n223, ZN => n218);
   U53 : OAI21_X1 port map( B1 => A(27), B2 => n224, A => B(27), ZN => n223);
   U54 : INV_X1 port map( A => A(27), ZN => n222);
   U55 : INV_X1 port map( A => n224, ZN => n221);
   U56 : XOR2_X1 port map( A => n225, B => n226, Z => S(27));
   U57 : XOR2_X1 port map( A => Ci, B => B(27), Z => n226);
   U58 : XOR2_X1 port map( A => n224, B => A(27), Z => n225);
   U59 : OAI21_X1 port map( B1 => n227, B2 => n228, A => n229, ZN => n224);
   U60 : OAI21_X1 port map( B1 => A(26), B2 => n230, A => B(26), ZN => n229);
   U61 : INV_X1 port map( A => A(26), ZN => n228);
   U62 : INV_X1 port map( A => n230, ZN => n227);
   U63 : XOR2_X1 port map( A => n231, B => n232, Z => S(26));
   U64 : XOR2_X1 port map( A => Ci, B => B(26), Z => n232);
   U65 : XOR2_X1 port map( A => n230, B => A(26), Z => n231);
   U66 : OAI21_X1 port map( B1 => n233, B2 => n234, A => n235, ZN => n230);
   U67 : OAI21_X1 port map( B1 => A(25), B2 => n236, A => B(25), ZN => n235);
   U68 : INV_X1 port map( A => A(25), ZN => n234);
   U69 : XOR2_X1 port map( A => n237, B => n238, Z => S(25));
   U70 : XOR2_X1 port map( A => Ci, B => B(25), Z => n238);
   U71 : XOR2_X1 port map( A => n236, B => A(25), Z => n237);
   U72 : INV_X1 port map( A => n233, ZN => n236);
   U73 : AOI22_X1 port map( A1 => n239, A2 => A(24), B1 => n240, B2 => B(24), 
                           ZN => n233);
   U74 : OR2_X1 port map( A1 => A(24), A2 => n239, ZN => n240);
   U75 : XOR2_X1 port map( A => n241, B => n242, Z => S(24));
   U76 : XOR2_X1 port map( A => Ci, B => B(24), Z => n242);
   U77 : XOR2_X1 port map( A => n239, B => A(24), Z => n241);
   U78 : INV_X1 port map( A => n243, ZN => n239);
   U79 : AOI22_X1 port map( A1 => n244, A2 => A(23), B1 => n245, B2 => B(23), 
                           ZN => n243);
   U80 : OR2_X1 port map( A1 => A(23), A2 => n244, ZN => n245);
   U81 : XOR2_X1 port map( A => n246, B => n247, Z => S(23));
   U82 : XOR2_X1 port map( A => Ci, B => B(23), Z => n247);
   U83 : XOR2_X1 port map( A => n244, B => A(23), Z => n246);
   U84 : OAI21_X1 port map( B1 => n248, B2 => n249, A => n250, ZN => n244);
   U85 : OAI21_X1 port map( B1 => A(22), B2 => n251, A => B(22), ZN => n250);
   U86 : XOR2_X1 port map( A => n252, B => n253, Z => S(22));
   U87 : XOR2_X1 port map( A => n249, B => n251, Z => n253);
   U88 : INV_X1 port map( A => n248, ZN => n251);
   U89 : AOI21_X1 port map( B1 => n254, B2 => A(21), A => n255, ZN => n248);
   U90 : INV_X1 port map( A => n256, ZN => n255);
   U91 : OAI21_X1 port map( B1 => n254, B2 => A(21), A => B(21), ZN => n256);
   U92 : INV_X1 port map( A => A(22), ZN => n249);
   U93 : XNOR2_X1 port map( A => B(22), B => Ci, ZN => n252);
   U94 : XOR2_X1 port map( A => n257, B => n258, Z => S(21));
   U95 : XNOR2_X1 port map( A => n254, B => A(21), ZN => n258);
   U96 : AOI21_X1 port map( B1 => n259, B2 => n260, A => n261, ZN => n254);
   U97 : AOI21_X1 port map( B1 => n262, B2 => A(20), A => B(20), ZN => n261);
   U98 : XNOR2_X1 port map( A => B(21), B => Ci, ZN => n257);
   U99 : XOR2_X1 port map( A => n263, B => n264, Z => S(20));
   U100 : XOR2_X1 port map( A => n259, B => n262, Z => n264);
   U101 : INV_X1 port map( A => n260, ZN => n262);
   U102 : AOI21_X1 port map( B1 => n265, B2 => A(19), A => n266, ZN => n260);
   U103 : INV_X1 port map( A => n267, ZN => n266);
   U104 : OAI21_X1 port map( B1 => n265, B2 => A(19), A => B(19), ZN => n267);
   U105 : INV_X1 port map( A => A(20), ZN => n259);
   U106 : XNOR2_X1 port map( A => B(20), B => Ci, ZN => n263);
   U107 : XOR2_X1 port map( A => n268, B => n269, Z => S(1));
   U108 : XOR2_X1 port map( A => n270, B => A(1), Z => n269);
   U109 : XNOR2_X1 port map( A => B(1), B => Ci, ZN => n268);
   U110 : XOR2_X1 port map( A => n271, B => n272, Z => S(19));
   U111 : XNOR2_X1 port map( A => n265, B => A(19), ZN => n272);
   U112 : AOI21_X1 port map( B1 => n273, B2 => n274, A => n275, ZN => n265);
   U113 : AOI21_X1 port map( B1 => n276, B2 => A(18), A => B(18), ZN => n275);
   U114 : XNOR2_X1 port map( A => B(19), B => Ci, ZN => n271);
   U115 : XOR2_X1 port map( A => n277, B => n278, Z => S(18));
   U116 : XOR2_X1 port map( A => n273, B => n276, Z => n278);
   U117 : INV_X1 port map( A => n274, ZN => n276);
   U118 : AOI21_X1 port map( B1 => n279, B2 => A(17), A => n280, ZN => n274);
   U119 : INV_X1 port map( A => n281, ZN => n280);
   U120 : OAI21_X1 port map( B1 => A(17), B2 => n279, A => B(17), ZN => n281);
   U121 : INV_X1 port map( A => A(18), ZN => n273);
   U122 : XNOR2_X1 port map( A => B(18), B => Ci, ZN => n277);
   U123 : XOR2_X1 port map( A => n282, B => n283, Z => S(17));
   U124 : XOR2_X1 port map( A => Ci, B => B(17), Z => n283);
   U125 : XOR2_X1 port map( A => A(17), B => n279, Z => n282);
   U126 : OAI21_X1 port map( B1 => n284, B2 => n285, A => n286, ZN => n279);
   U127 : OAI21_X1 port map( B1 => n287, B2 => A(16), A => B(16), ZN => n286);
   U128 : INV_X1 port map( A => n284, ZN => n287);
   U129 : INV_X1 port map( A => A(16), ZN => n285);
   U130 : XOR2_X1 port map( A => n288, B => n289, Z => S(16));
   U131 : XOR2_X1 port map( A => n284, B => A(16), Z => n289);
   U132 : OAI21_X1 port map( B1 => A(15), B2 => n290, A => n291, ZN => n284);
   U133 : INV_X1 port map( A => n292, ZN => n291);
   U134 : AOI21_X1 port map( B1 => n290, B2 => A(15), A => B(15), ZN => n292);
   U135 : XNOR2_X1 port map( A => B(16), B => Ci, ZN => n288);
   U136 : XOR2_X1 port map( A => n293, B => n294, Z => S(15));
   U137 : XNOR2_X1 port map( A => n290, B => A(15), ZN => n294);
   U138 : AOI21_X1 port map( B1 => n295, B2 => n296, A => n297, ZN => n290);
   U139 : AOI21_X1 port map( B1 => n298, B2 => A(14), A => B(14), ZN => n297);
   U140 : INV_X1 port map( A => n296, ZN => n298);
   U141 : INV_X1 port map( A => A(14), ZN => n295);
   U142 : XNOR2_X1 port map( A => B(15), B => Ci, ZN => n293);
   U143 : XOR2_X1 port map( A => n299, B => n300, Z => S(14));
   U144 : XOR2_X1 port map( A => A(14), B => n296, Z => n300);
   U145 : AOI21_X1 port map( B1 => n301, B2 => A(13), A => n302, ZN => n296);
   U146 : INV_X1 port map( A => n303, ZN => n302);
   U147 : OAI21_X1 port map( B1 => n301, B2 => A(13), A => B(13), ZN => n303);
   U148 : XNOR2_X1 port map( A => B(14), B => Ci, ZN => n299);
   U149 : XOR2_X1 port map( A => n304, B => n305, Z => S(13));
   U150 : XNOR2_X1 port map( A => n301, B => A(13), ZN => n305);
   U151 : AOI21_X1 port map( B1 => n306, B2 => n307, A => n308, ZN => n301);
   U152 : AOI21_X1 port map( B1 => n309, B2 => A(12), A => B(12), ZN => n308);
   U153 : INV_X1 port map( A => A(12), ZN => n306);
   U154 : XNOR2_X1 port map( A => B(13), B => Ci, ZN => n304);
   U155 : XOR2_X1 port map( A => n310, B => n311, Z => S(12));
   U156 : XOR2_X1 port map( A => A(12), B => n307, Z => n311);
   U157 : INV_X1 port map( A => n309, ZN => n307);
   U158 : OAI21_X1 port map( B1 => n312, B2 => n313, A => n314, ZN => n309);
   U159 : OAI21_X1 port map( B1 => n315, B2 => A(11), A => B(11), ZN => n314);
   U160 : INV_X1 port map( A => n312, ZN => n315);
   U161 : INV_X1 port map( A => A(11), ZN => n313);
   U162 : XNOR2_X1 port map( A => B(12), B => Ci, ZN => n310);
   U163 : XOR2_X1 port map( A => n316, B => n317, Z => S(11));
   U164 : XOR2_X1 port map( A => n312, B => A(11), Z => n317);
   U165 : OAI22_X1 port map( A1 => A(10), A2 => n318, B1 => B(10), B2 => n319, 
                           ZN => n312);
   U166 : AND2_X1 port map( A1 => n318, A2 => A(10), ZN => n319);
   U167 : XNOR2_X1 port map( A => B(11), B => Ci, ZN => n316);
   U168 : XOR2_X1 port map( A => n320, B => n321, Z => S(10));
   U169 : XOR2_X1 port map( A => Ci, B => B(10), Z => n321);
   U170 : XOR2_X1 port map( A => A(10), B => n318, Z => n320);
   U171 : OAI21_X1 port map( B1 => n180, B2 => n322, A => n323, ZN => n318);
   U172 : OAI21_X1 port map( B1 => n324, B2 => A(9), A => B(9), ZN => n323);
   U173 : INV_X1 port map( A => n180, ZN => n324);
   U174 : INV_X1 port map( A => A(9), ZN => n322);
   U175 : OAI22_X1 port map( A1 => A(8), A2 => n183, B1 => B(8), B2 => n325, ZN
                           => n180);
   U176 : AND2_X1 port map( A1 => n183, A2 => A(8), ZN => n325);
   U177 : OAI21_X1 port map( B1 => n186, B2 => n326, A => n327, ZN => n183);
   U178 : OAI21_X1 port map( B1 => n328, B2 => A(7), A => B(7), ZN => n327);
   U179 : INV_X1 port map( A => n186, ZN => n328);
   U180 : INV_X1 port map( A => A(7), ZN => n326);
   U181 : OAI22_X1 port map( A1 => A(6), A2 => n189, B1 => B(6), B2 => n329, ZN
                           => n186);
   U182 : AND2_X1 port map( A1 => n189, A2 => A(6), ZN => n329);
   U183 : OAI21_X1 port map( B1 => n330, B2 => n331, A => n332, ZN => n189);
   U184 : OAI21_X1 port map( B1 => n192, B2 => A(5), A => B(5), ZN => n332);
   U185 : INV_X1 port map( A => n330, ZN => n192);
   U186 : INV_X1 port map( A => A(5), ZN => n331);
   U187 : OAI21_X1 port map( B1 => A(4), B2 => n333, A => n334, ZN => n330);
   U188 : INV_X1 port map( A => n335, ZN => n334);
   U189 : AOI21_X1 port map( B1 => n333, B2 => A(4), A => B(4), ZN => n335);
   U190 : INV_X1 port map( A => n195, ZN => n333);
   U191 : OAI21_X1 port map( B1 => A(3), B2 => n336, A => n337, ZN => n195);
   U192 : INV_X1 port map( A => n338, ZN => n337);
   U193 : AOI21_X1 port map( B1 => n336, B2 => A(3), A => B(3), ZN => n338);
   U194 : INV_X1 port map( A => n198, ZN => n336);
   U195 : OAI21_X1 port map( B1 => A(2), B2 => n339, A => n340, ZN => n198);
   U196 : INV_X1 port map( A => n341, ZN => n340);
   U197 : AOI21_X1 port map( B1 => n339, B2 => A(2), A => B(2), ZN => n341);
   U198 : INV_X1 port map( A => n212, ZN => n339);
   U199 : OAI21_X1 port map( B1 => A(1), B2 => n342, A => n343, ZN => n212);
   U200 : INV_X1 port map( A => n344, ZN => n343);
   U201 : AOI21_X1 port map( B1 => n342, B2 => A(1), A => B(1), ZN => n344);
   U202 : INV_X1 port map( A => n270, ZN => n342);
   U203 : MUX2_X1 port map( A => n345, B => n346, S => Ci, Z => S(0));
   U204 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n270, ZN => n346);
   U205 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n270);
   U206 : XOR2_X1 port map( A => B(0), B => A(0), Z => n345);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity writeBack_nbits32 is

   port( LMD_OUT, ALUREG_OUTPUT : in std_logic_vector (31 downto 0);  
         WB_MUX_SEL : in std_logic;  DATAIN_RF : out std_logic_vector (31 
         downto 0));

end writeBack_nbits32;

architecture SYN_STRUCTURAL of writeBack_nbits32 is

   component MUX21_GENERIC_bits32_1
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;

begin
   
   MUXWB : MUX21_GENERIC_bits32_1 port map( A(31) => ALUREG_OUTPUT(31), A(30) 
                           => ALUREG_OUTPUT(30), A(29) => ALUREG_OUTPUT(29), 
                           A(28) => ALUREG_OUTPUT(28), A(27) => 
                           ALUREG_OUTPUT(27), A(26) => ALUREG_OUTPUT(26), A(25)
                           => ALUREG_OUTPUT(25), A(24) => ALUREG_OUTPUT(24), 
                           A(23) => ALUREG_OUTPUT(23), A(22) => 
                           ALUREG_OUTPUT(22), A(21) => ALUREG_OUTPUT(21), A(20)
                           => ALUREG_OUTPUT(20), A(19) => ALUREG_OUTPUT(19), 
                           A(18) => ALUREG_OUTPUT(18), A(17) => 
                           ALUREG_OUTPUT(17), A(16) => ALUREG_OUTPUT(16), A(15)
                           => ALUREG_OUTPUT(15), A(14) => ALUREG_OUTPUT(14), 
                           A(13) => ALUREG_OUTPUT(13), A(12) => 
                           ALUREG_OUTPUT(12), A(11) => ALUREG_OUTPUT(11), A(10)
                           => ALUREG_OUTPUT(10), A(9) => ALUREG_OUTPUT(9), A(8)
                           => ALUREG_OUTPUT(8), A(7) => ALUREG_OUTPUT(7), A(6) 
                           => ALUREG_OUTPUT(6), A(5) => ALUREG_OUTPUT(5), A(4) 
                           => ALUREG_OUTPUT(4), A(3) => ALUREG_OUTPUT(3), A(2) 
                           => ALUREG_OUTPUT(2), A(1) => ALUREG_OUTPUT(1), A(0) 
                           => ALUREG_OUTPUT(0), B(31) => LMD_OUT(31), B(30) => 
                           LMD_OUT(30), B(29) => LMD_OUT(29), B(28) => 
                           LMD_OUT(28), B(27) => LMD_OUT(27), B(26) => 
                           LMD_OUT(26), B(25) => LMD_OUT(25), B(24) => 
                           LMD_OUT(24), B(23) => LMD_OUT(23), B(22) => 
                           LMD_OUT(22), B(21) => LMD_OUT(21), B(20) => 
                           LMD_OUT(20), B(19) => LMD_OUT(19), B(18) => 
                           LMD_OUT(18), B(17) => LMD_OUT(17), B(16) => 
                           LMD_OUT(16), B(15) => LMD_OUT(15), B(14) => 
                           LMD_OUT(14), B(13) => LMD_OUT(13), B(12) => 
                           LMD_OUT(12), B(11) => LMD_OUT(11), B(10) => 
                           LMD_OUT(10), B(9) => LMD_OUT(9), B(8) => LMD_OUT(8),
                           B(7) => LMD_OUT(7), B(6) => LMD_OUT(6), B(5) => 
                           LMD_OUT(5), B(4) => LMD_OUT(4), B(3) => LMD_OUT(3), 
                           B(2) => LMD_OUT(2), B(1) => LMD_OUT(1), B(0) => 
                           LMD_OUT(0), S => WB_MUX_SEL, Y(31) => DATAIN_RF(31),
                           Y(30) => DATAIN_RF(30), Y(29) => DATAIN_RF(29), 
                           Y(28) => DATAIN_RF(28), Y(27) => DATAIN_RF(27), 
                           Y(26) => DATAIN_RF(26), Y(25) => DATAIN_RF(25), 
                           Y(24) => DATAIN_RF(24), Y(23) => DATAIN_RF(23), 
                           Y(22) => DATAIN_RF(22), Y(21) => DATAIN_RF(21), 
                           Y(20) => DATAIN_RF(20), Y(19) => DATAIN_RF(19), 
                           Y(18) => DATAIN_RF(18), Y(17) => DATAIN_RF(17), 
                           Y(16) => DATAIN_RF(16), Y(15) => DATAIN_RF(15), 
                           Y(14) => DATAIN_RF(14), Y(13) => DATAIN_RF(13), 
                           Y(12) => DATAIN_RF(12), Y(11) => DATAIN_RF(11), 
                           Y(10) => DATAIN_RF(10), Y(9) => DATAIN_RF(9), Y(8) 
                           => DATAIN_RF(8), Y(7) => DATAIN_RF(7), Y(6) => 
                           DATAIN_RF(6), Y(5) => DATAIN_RF(5), Y(4) => 
                           DATAIN_RF(4), Y(3) => DATAIN_RF(3), Y(2) => 
                           DATAIN_RF(2), Y(1) => DATAIN_RF(1), Y(0) => 
                           DATAIN_RF(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity memoryUnit_nbits32 is

   port( clk, rst, LMD_LATCH_EN, JUMP_EN : in std_logic;  DRAM_DATA, 
         ALUREG_OUTPUT, NPC_OUT : in std_logic_vector (31 downto 0);  COND_OUT 
         : in std_logic;  DRAM_DATAout, TO_PC_OUT, ALU_OUT2 : out 
         std_logic_vector (31 downto 0);  IR_IN4 : in std_logic_vector (31 
         downto 0);  IR_OUT4 : out std_logic_vector (31 downto 0));

end memoryUnit_nbits32;

architecture SYN_STRUCTURAL of memoryUnit_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component register_generic_nbits32_1
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_2
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_bits32_2
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, muxjmp_to_mux, n3, n4 : std_logic;

begin
   DRAM_DATAout <= ( DRAM_DATA(31), DRAM_DATA(30), DRAM_DATA(29), DRAM_DATA(28)
      , DRAM_DATA(27), DRAM_DATA(26), DRAM_DATA(25), DRAM_DATA(24), 
      DRAM_DATA(23), DRAM_DATA(22), DRAM_DATA(21), DRAM_DATA(20), DRAM_DATA(19)
      , DRAM_DATA(18), DRAM_DATA(17), DRAM_DATA(16), DRAM_DATA(15), 
      DRAM_DATA(14), DRAM_DATA(13), DRAM_DATA(12), DRAM_DATA(11), DRAM_DATA(10)
      , DRAM_DATA(9), DRAM_DATA(8), DRAM_DATA(7), DRAM_DATA(6), DRAM_DATA(5), 
      DRAM_DATA(4), DRAM_DATA(3), DRAM_DATA(2), DRAM_DATA(1), DRAM_DATA(0) );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   JUMPMUX : MUX21 port map( A => COND_OUT, B => X_Logic0_port, S => JUMP_EN, Y
                           => muxjmp_to_mux);
   MUX_PC : MUX21_GENERIC_bits32_2 port map( A(31) => ALUREG_OUTPUT(31), A(30) 
                           => ALUREG_OUTPUT(30), A(29) => ALUREG_OUTPUT(29), 
                           A(28) => ALUREG_OUTPUT(28), A(27) => 
                           ALUREG_OUTPUT(27), A(26) => ALUREG_OUTPUT(26), A(25)
                           => ALUREG_OUTPUT(25), A(24) => ALUREG_OUTPUT(24), 
                           A(23) => ALUREG_OUTPUT(23), A(22) => 
                           ALUREG_OUTPUT(22), A(21) => ALUREG_OUTPUT(21), A(20)
                           => ALUREG_OUTPUT(20), A(19) => ALUREG_OUTPUT(19), 
                           A(18) => ALUREG_OUTPUT(18), A(17) => 
                           ALUREG_OUTPUT(17), A(16) => ALUREG_OUTPUT(16), A(15)
                           => ALUREG_OUTPUT(15), A(14) => ALUREG_OUTPUT(14), 
                           A(13) => ALUREG_OUTPUT(13), A(12) => 
                           ALUREG_OUTPUT(12), A(11) => ALUREG_OUTPUT(11), A(10)
                           => ALUREG_OUTPUT(10), A(9) => ALUREG_OUTPUT(9), A(8)
                           => ALUREG_OUTPUT(8), A(7) => ALUREG_OUTPUT(7), A(6) 
                           => ALUREG_OUTPUT(6), A(5) => ALUREG_OUTPUT(5), A(4) 
                           => ALUREG_OUTPUT(4), A(3) => ALUREG_OUTPUT(3), A(2) 
                           => ALUREG_OUTPUT(2), A(1) => ALUREG_OUTPUT(1), A(0) 
                           => ALUREG_OUTPUT(0), B(31) => NPC_OUT(31), B(30) => 
                           NPC_OUT(30), B(29) => NPC_OUT(29), B(28) => 
                           NPC_OUT(28), B(27) => NPC_OUT(27), B(26) => 
                           NPC_OUT(26), B(25) => NPC_OUT(25), B(24) => 
                           NPC_OUT(24), B(23) => NPC_OUT(23), B(22) => 
                           NPC_OUT(22), B(21) => NPC_OUT(21), B(20) => 
                           NPC_OUT(20), B(19) => NPC_OUT(19), B(18) => 
                           NPC_OUT(18), B(17) => NPC_OUT(17), B(16) => 
                           NPC_OUT(16), B(15) => NPC_OUT(15), B(14) => 
                           NPC_OUT(14), B(13) => NPC_OUT(13), B(12) => 
                           NPC_OUT(12), B(11) => NPC_OUT(11), B(10) => 
                           NPC_OUT(10), B(9) => NPC_OUT(9), B(8) => NPC_OUT(8),
                           B(7) => NPC_OUT(7), B(6) => NPC_OUT(6), B(5) => 
                           NPC_OUT(5), B(4) => NPC_OUT(4), B(3) => NPC_OUT(3), 
                           B(2) => NPC_OUT(2), B(1) => NPC_OUT(1), B(0) => 
                           NPC_OUT(0), S => muxjmp_to_mux, Y(31) => 
                           TO_PC_OUT(31), Y(30) => TO_PC_OUT(30), Y(29) => 
                           TO_PC_OUT(29), Y(28) => TO_PC_OUT(28), Y(27) => 
                           TO_PC_OUT(27), Y(26) => TO_PC_OUT(26), Y(25) => 
                           TO_PC_OUT(25), Y(24) => TO_PC_OUT(24), Y(23) => 
                           TO_PC_OUT(23), Y(22) => TO_PC_OUT(22), Y(21) => 
                           TO_PC_OUT(21), Y(20) => TO_PC_OUT(20), Y(19) => 
                           TO_PC_OUT(19), Y(18) => TO_PC_OUT(18), Y(17) => 
                           TO_PC_OUT(17), Y(16) => TO_PC_OUT(16), Y(15) => 
                           TO_PC_OUT(15), Y(14) => TO_PC_OUT(14), Y(13) => 
                           TO_PC_OUT(13), Y(12) => TO_PC_OUT(12), Y(11) => 
                           TO_PC_OUT(11), Y(10) => TO_PC_OUT(10), Y(9) => 
                           TO_PC_OUT(9), Y(8) => TO_PC_OUT(8), Y(7) => 
                           TO_PC_OUT(7), Y(6) => TO_PC_OUT(6), Y(5) => 
                           TO_PC_OUT(5), Y(4) => TO_PC_OUT(4), Y(3) => 
                           TO_PC_OUT(3), Y(2) => TO_PC_OUT(2), Y(1) => 
                           TO_PC_OUT(1), Y(0) => TO_PC_OUT(0));
   ALU_OUT2r : register_generic_nbits32_2 port map( data_in(31) => 
                           ALUREG_OUTPUT(31), data_in(30) => ALUREG_OUTPUT(30),
                           data_in(29) => ALUREG_OUTPUT(29), data_in(28) => 
                           ALUREG_OUTPUT(28), data_in(27) => ALUREG_OUTPUT(27),
                           data_in(26) => ALUREG_OUTPUT(26), data_in(25) => 
                           ALUREG_OUTPUT(25), data_in(24) => ALUREG_OUTPUT(24),
                           data_in(23) => ALUREG_OUTPUT(23), data_in(22) => 
                           ALUREG_OUTPUT(22), data_in(21) => ALUREG_OUTPUT(21),
                           data_in(20) => ALUREG_OUTPUT(20), data_in(19) => 
                           ALUREG_OUTPUT(19), data_in(18) => ALUREG_OUTPUT(18),
                           data_in(17) => ALUREG_OUTPUT(17), data_in(16) => 
                           ALUREG_OUTPUT(16), data_in(15) => ALUREG_OUTPUT(15),
                           data_in(14) => ALUREG_OUTPUT(14), data_in(13) => 
                           ALUREG_OUTPUT(13), data_in(12) => ALUREG_OUTPUT(12),
                           data_in(11) => ALUREG_OUTPUT(11), data_in(10) => 
                           ALUREG_OUTPUT(10), data_in(9) => ALUREG_OUTPUT(9), 
                           data_in(8) => ALUREG_OUTPUT(8), data_in(7) => 
                           ALUREG_OUTPUT(7), data_in(6) => ALUREG_OUTPUT(6), 
                           data_in(5) => ALUREG_OUTPUT(5), data_in(4) => 
                           ALUREG_OUTPUT(4), data_in(3) => ALUREG_OUTPUT(3), 
                           data_in(2) => ALUREG_OUTPUT(2), data_in(1) => 
                           ALUREG_OUTPUT(1), data_in(0) => ALUREG_OUTPUT(0), CK
                           => n4, RESET => n3, ENABLE => X_Logic1_port, 
                           data_out(31) => ALU_OUT2(31), data_out(30) => 
                           ALU_OUT2(30), data_out(29) => ALU_OUT2(29), 
                           data_out(28) => ALU_OUT2(28), data_out(27) => 
                           ALU_OUT2(27), data_out(26) => ALU_OUT2(26), 
                           data_out(25) => ALU_OUT2(25), data_out(24) => 
                           ALU_OUT2(24), data_out(23) => ALU_OUT2(23), 
                           data_out(22) => ALU_OUT2(22), data_out(21) => 
                           ALU_OUT2(21), data_out(20) => ALU_OUT2(20), 
                           data_out(19) => ALU_OUT2(19), data_out(18) => 
                           ALU_OUT2(18), data_out(17) => ALU_OUT2(17), 
                           data_out(16) => ALU_OUT2(16), data_out(15) => 
                           ALU_OUT2(15), data_out(14) => ALU_OUT2(14), 
                           data_out(13) => ALU_OUT2(13), data_out(12) => 
                           ALU_OUT2(12), data_out(11) => ALU_OUT2(11), 
                           data_out(10) => ALU_OUT2(10), data_out(9) => 
                           ALU_OUT2(9), data_out(8) => ALU_OUT2(8), data_out(7)
                           => ALU_OUT2(7), data_out(6) => ALU_OUT2(6), 
                           data_out(5) => ALU_OUT2(5), data_out(4) => 
                           ALU_OUT2(4), data_out(3) => ALU_OUT2(3), data_out(2)
                           => ALU_OUT2(2), data_out(1) => ALU_OUT2(1), 
                           data_out(0) => ALU_OUT2(0));
   IR4 : register_generic_nbits32_1 port map( data_in(31) => IR_IN4(31), 
                           data_in(30) => IR_IN4(30), data_in(29) => IR_IN4(29)
                           , data_in(28) => IR_IN4(28), data_in(27) => 
                           IR_IN4(27), data_in(26) => IR_IN4(26), data_in(25) 
                           => IR_IN4(25), data_in(24) => IR_IN4(24), 
                           data_in(23) => IR_IN4(23), data_in(22) => IR_IN4(22)
                           , data_in(21) => IR_IN4(21), data_in(20) => 
                           IR_IN4(20), data_in(19) => IR_IN4(19), data_in(18) 
                           => IR_IN4(18), data_in(17) => IR_IN4(17), 
                           data_in(16) => IR_IN4(16), data_in(15) => IR_IN4(15)
                           , data_in(14) => IR_IN4(14), data_in(13) => 
                           IR_IN4(13), data_in(12) => IR_IN4(12), data_in(11) 
                           => IR_IN4(11), data_in(10) => IR_IN4(10), data_in(9)
                           => IR_IN4(9), data_in(8) => IR_IN4(8), data_in(7) =>
                           IR_IN4(7), data_in(6) => IR_IN4(6), data_in(5) => 
                           IR_IN4(5), data_in(4) => IR_IN4(4), data_in(3) => 
                           IR_IN4(3), data_in(2) => IR_IN4(2), data_in(1) => 
                           IR_IN4(1), data_in(0) => IR_IN4(0), CK => n4, RESET 
                           => n3, ENABLE => X_Logic1_port, data_out(31) => 
                           IR_OUT4(31), data_out(30) => IR_OUT4(30), 
                           data_out(29) => IR_OUT4(29), data_out(28) => 
                           IR_OUT4(28), data_out(27) => IR_OUT4(27), 
                           data_out(26) => IR_OUT4(26), data_out(25) => 
                           IR_OUT4(25), data_out(24) => IR_OUT4(24), 
                           data_out(23) => IR_OUT4(23), data_out(22) => 
                           IR_OUT4(22), data_out(21) => IR_OUT4(21), 
                           data_out(20) => IR_OUT4(20), data_out(19) => 
                           IR_OUT4(19), data_out(18) => IR_OUT4(18), 
                           data_out(17) => IR_OUT4(17), data_out(16) => 
                           IR_OUT4(16), data_out(15) => IR_OUT4(15), 
                           data_out(14) => IR_OUT4(14), data_out(13) => 
                           IR_OUT4(13), data_out(12) => IR_OUT4(12), 
                           data_out(11) => IR_OUT4(11), data_out(10) => 
                           IR_OUT4(10), data_out(9) => IR_OUT4(9), data_out(8) 
                           => IR_OUT4(8), data_out(7) => IR_OUT4(7), 
                           data_out(6) => IR_OUT4(6), data_out(5) => IR_OUT4(5)
                           , data_out(4) => IR_OUT4(4), data_out(3) => 
                           IR_OUT4(3), data_out(2) => IR_OUT4(2), data_out(1) 
                           => IR_OUT4(1), data_out(0) => IR_OUT4(0));
   U3 : BUF_X1 port map( A => rst, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity executionUnit_nbits32 is

   port( clk, rst, ALU_OUTREG_ENABLE, MUXA_SEL, MUXB_SEL, COND_ENABLE : in 
         std_logic;  ALU_BITS : in std_logic_vector (0 to 3);  NPC_OUT, A_out, 
         B_out, Imm_out : in std_logic_vector (31 downto 0);  ALUREG_OUTPUT : 
         out std_logic_vector (31 downto 0);  COND_OUT : out std_logic;  IR_IN3
         : in std_logic_vector (31 downto 0);  IR_OUT3, B_outreg : out 
         std_logic_vector (31 downto 0));

end executionUnit_nbits32;

architecture SYN_STRUCTURAL of executionUnit_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_0
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component XNOR_logic
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component alu_nbits32
      port( FUNC : in std_logic_vector (0 to 3);  A, B : in std_logic_vector 
            (31 downto 0);  OUTALU : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_3
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_4
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_5
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_bits32_3
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_bits32_0
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component ZERO_DEC_bits32
      port( data : in std_logic_vector (31 downto 0);  zero_detect : out 
            std_logic);
   end component;
   
   signal X_Logic1_port, ZERO_DEC_OUT, MUX1_OUT_31_port, MUX1_OUT_30_port, 
      MUX1_OUT_29_port, MUX1_OUT_28_port, MUX1_OUT_27_port, MUX1_OUT_26_port, 
      MUX1_OUT_25_port, MUX1_OUT_24_port, MUX1_OUT_23_port, MUX1_OUT_22_port, 
      MUX1_OUT_21_port, MUX1_OUT_20_port, MUX1_OUT_19_port, MUX1_OUT_18_port, 
      MUX1_OUT_17_port, MUX1_OUT_16_port, MUX1_OUT_15_port, MUX1_OUT_14_port, 
      MUX1_OUT_13_port, MUX1_OUT_12_port, MUX1_OUT_11_port, MUX1_OUT_10_port, 
      MUX1_OUT_9_port, MUX1_OUT_8_port, MUX1_OUT_7_port, MUX1_OUT_6_port, 
      MUX1_OUT_5_port, MUX1_OUT_4_port, MUX1_OUT_3_port, MUX1_OUT_2_port, 
      MUX1_OUT_1_port, MUX1_OUT_0_port, MUX2_OUT_31_port, MUX2_OUT_30_port, 
      MUX2_OUT_29_port, MUX2_OUT_28_port, MUX2_OUT_27_port, MUX2_OUT_26_port, 
      MUX2_OUT_25_port, MUX2_OUT_24_port, MUX2_OUT_23_port, MUX2_OUT_22_port, 
      MUX2_OUT_21_port, MUX2_OUT_20_port, MUX2_OUT_19_port, MUX2_OUT_18_port, 
      MUX2_OUT_17_port, MUX2_OUT_16_port, MUX2_OUT_15_port, MUX2_OUT_14_port, 
      MUX2_OUT_13_port, MUX2_OUT_12_port, MUX2_OUT_11_port, MUX2_OUT_10_port, 
      MUX2_OUT_9_port, MUX2_OUT_8_port, MUX2_OUT_7_port, MUX2_OUT_6_port, 
      MUX2_OUT_5_port, MUX2_OUT_4_port, MUX2_OUT_3_port, MUX2_OUT_2_port, 
      MUX2_OUT_1_port, MUX2_OUT_0_port, ALU_output_31_port, ALU_output_30_port,
      ALU_output_29_port, ALU_output_28_port, ALU_output_27_port, 
      ALU_output_26_port, ALU_output_25_port, ALU_output_24_port, 
      ALU_output_23_port, ALU_output_22_port, ALU_output_21_port, 
      ALU_output_20_port, ALU_output_19_port, ALU_output_18_port, 
      ALU_output_17_port, ALU_output_16_port, ALU_output_15_port, 
      ALU_output_14_port, ALU_output_13_port, ALU_output_12_port, 
      ALU_output_11_port, ALU_output_10_port, ALU_output_9_port, 
      ALU_output_8_port, ALU_output_7_port, ALU_output_6_port, 
      ALU_output_5_port, ALU_output_4_port, ALU_output_3_port, 
      ALU_output_2_port, ALU_output_1_port, ALU_output_0_port, XNOR_OUT, n3, n4
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   zerodec : ZERO_DEC_bits32 port map( data(31) => A_out(31), data(30) => 
                           A_out(30), data(29) => A_out(29), data(28) => 
                           A_out(28), data(27) => A_out(27), data(26) => 
                           A_out(26), data(25) => A_out(25), data(24) => 
                           A_out(24), data(23) => A_out(23), data(22) => 
                           A_out(22), data(21) => A_out(21), data(20) => 
                           A_out(20), data(19) => A_out(19), data(18) => 
                           A_out(18), data(17) => A_out(17), data(16) => 
                           A_out(16), data(15) => A_out(15), data(14) => 
                           A_out(14), data(13) => A_out(13), data(12) => 
                           A_out(12), data(11) => A_out(11), data(10) => 
                           A_out(10), data(9) => A_out(9), data(8) => A_out(8),
                           data(7) => A_out(7), data(6) => A_out(6), data(5) =>
                           A_out(5), data(4) => A_out(4), data(3) => A_out(3), 
                           data(2) => A_out(2), data(1) => A_out(1), data(0) =>
                           A_out(0), zero_detect => ZERO_DEC_OUT);
   mux1 : MUX21_GENERIC_bits32_0 port map( A(31) => A_out(31), A(30) => 
                           A_out(30), A(29) => A_out(29), A(28) => A_out(28), 
                           A(27) => A_out(27), A(26) => A_out(26), A(25) => 
                           A_out(25), A(24) => A_out(24), A(23) => A_out(23), 
                           A(22) => A_out(22), A(21) => A_out(21), A(20) => 
                           A_out(20), A(19) => A_out(19), A(18) => A_out(18), 
                           A(17) => A_out(17), A(16) => A_out(16), A(15) => 
                           A_out(15), A(14) => A_out(14), A(13) => A_out(13), 
                           A(12) => A_out(12), A(11) => A_out(11), A(10) => 
                           A_out(10), A(9) => A_out(9), A(8) => A_out(8), A(7) 
                           => A_out(7), A(6) => A_out(6), A(5) => A_out(5), 
                           A(4) => A_out(4), A(3) => A_out(3), A(2) => A_out(2)
                           , A(1) => A_out(1), A(0) => A_out(0), B(31) => 
                           NPC_OUT(31), B(30) => NPC_OUT(30), B(29) => 
                           NPC_OUT(29), B(28) => NPC_OUT(28), B(27) => 
                           NPC_OUT(27), B(26) => NPC_OUT(26), B(25) => 
                           NPC_OUT(25), B(24) => NPC_OUT(24), B(23) => 
                           NPC_OUT(23), B(22) => NPC_OUT(22), B(21) => 
                           NPC_OUT(21), B(20) => NPC_OUT(20), B(19) => 
                           NPC_OUT(19), B(18) => NPC_OUT(18), B(17) => 
                           NPC_OUT(17), B(16) => NPC_OUT(16), B(15) => 
                           NPC_OUT(15), B(14) => NPC_OUT(14), B(13) => 
                           NPC_OUT(13), B(12) => NPC_OUT(12), B(11) => 
                           NPC_OUT(11), B(10) => NPC_OUT(10), B(9) => 
                           NPC_OUT(9), B(8) => NPC_OUT(8), B(7) => NPC_OUT(7), 
                           B(6) => NPC_OUT(6), B(5) => NPC_OUT(5), B(4) => 
                           NPC_OUT(4), B(3) => NPC_OUT(3), B(2) => NPC_OUT(2), 
                           B(1) => NPC_OUT(1), B(0) => NPC_OUT(0), S => 
                           MUXA_SEL, Y(31) => MUX1_OUT_31_port, Y(30) => 
                           MUX1_OUT_30_port, Y(29) => MUX1_OUT_29_port, Y(28) 
                           => MUX1_OUT_28_port, Y(27) => MUX1_OUT_27_port, 
                           Y(26) => MUX1_OUT_26_port, Y(25) => MUX1_OUT_25_port
                           , Y(24) => MUX1_OUT_24_port, Y(23) => 
                           MUX1_OUT_23_port, Y(22) => MUX1_OUT_22_port, Y(21) 
                           => MUX1_OUT_21_port, Y(20) => MUX1_OUT_20_port, 
                           Y(19) => MUX1_OUT_19_port, Y(18) => MUX1_OUT_18_port
                           , Y(17) => MUX1_OUT_17_port, Y(16) => 
                           MUX1_OUT_16_port, Y(15) => MUX1_OUT_15_port, Y(14) 
                           => MUX1_OUT_14_port, Y(13) => MUX1_OUT_13_port, 
                           Y(12) => MUX1_OUT_12_port, Y(11) => MUX1_OUT_11_port
                           , Y(10) => MUX1_OUT_10_port, Y(9) => MUX1_OUT_9_port
                           , Y(8) => MUX1_OUT_8_port, Y(7) => MUX1_OUT_7_port, 
                           Y(6) => MUX1_OUT_6_port, Y(5) => MUX1_OUT_5_port, 
                           Y(4) => MUX1_OUT_4_port, Y(3) => MUX1_OUT_3_port, 
                           Y(2) => MUX1_OUT_2_port, Y(1) => MUX1_OUT_1_port, 
                           Y(0) => MUX1_OUT_0_port);
   mux2 : MUX21_GENERIC_bits32_3 port map( A(31) => Imm_out(31), A(30) => 
                           Imm_out(30), A(29) => Imm_out(29), A(28) => 
                           Imm_out(28), A(27) => Imm_out(27), A(26) => 
                           Imm_out(26), A(25) => Imm_out(25), A(24) => 
                           Imm_out(24), A(23) => Imm_out(23), A(22) => 
                           Imm_out(22), A(21) => Imm_out(21), A(20) => 
                           Imm_out(20), A(19) => Imm_out(19), A(18) => 
                           Imm_out(18), A(17) => Imm_out(17), A(16) => 
                           Imm_out(16), A(15) => Imm_out(15), A(14) => 
                           Imm_out(14), A(13) => Imm_out(13), A(12) => 
                           Imm_out(12), A(11) => Imm_out(11), A(10) => 
                           Imm_out(10), A(9) => Imm_out(9), A(8) => Imm_out(8),
                           A(7) => Imm_out(7), A(6) => Imm_out(6), A(5) => 
                           Imm_out(5), A(4) => Imm_out(4), A(3) => Imm_out(3), 
                           A(2) => Imm_out(2), A(1) => Imm_out(1), A(0) => 
                           Imm_out(0), B(31) => B_out(31), B(30) => B_out(30), 
                           B(29) => B_out(29), B(28) => B_out(28), B(27) => 
                           B_out(27), B(26) => B_out(26), B(25) => B_out(25), 
                           B(24) => B_out(24), B(23) => B_out(23), B(22) => 
                           B_out(22), B(21) => B_out(21), B(20) => B_out(20), 
                           B(19) => B_out(19), B(18) => B_out(18), B(17) => 
                           B_out(17), B(16) => B_out(16), B(15) => B_out(15), 
                           B(14) => B_out(14), B(13) => B_out(13), B(12) => 
                           B_out(12), B(11) => B_out(11), B(10) => B_out(10), 
                           B(9) => B_out(9), B(8) => B_out(8), B(7) => B_out(7)
                           , B(6) => B_out(6), B(5) => B_out(5), B(4) => 
                           B_out(4), B(3) => B_out(3), B(2) => B_out(2), B(1) 
                           => B_out(1), B(0) => B_out(0), S => MUXB_SEL, Y(31) 
                           => MUX2_OUT_31_port, Y(30) => MUX2_OUT_30_port, 
                           Y(29) => MUX2_OUT_29_port, Y(28) => MUX2_OUT_28_port
                           , Y(27) => MUX2_OUT_27_port, Y(26) => 
                           MUX2_OUT_26_port, Y(25) => MUX2_OUT_25_port, Y(24) 
                           => MUX2_OUT_24_port, Y(23) => MUX2_OUT_23_port, 
                           Y(22) => MUX2_OUT_22_port, Y(21) => MUX2_OUT_21_port
                           , Y(20) => MUX2_OUT_20_port, Y(19) => 
                           MUX2_OUT_19_port, Y(18) => MUX2_OUT_18_port, Y(17) 
                           => MUX2_OUT_17_port, Y(16) => MUX2_OUT_16_port, 
                           Y(15) => MUX2_OUT_15_port, Y(14) => MUX2_OUT_14_port
                           , Y(13) => MUX2_OUT_13_port, Y(12) => 
                           MUX2_OUT_12_port, Y(11) => MUX2_OUT_11_port, Y(10) 
                           => MUX2_OUT_10_port, Y(9) => MUX2_OUT_9_port, Y(8) 
                           => MUX2_OUT_8_port, Y(7) => MUX2_OUT_7_port, Y(6) =>
                           MUX2_OUT_6_port, Y(5) => MUX2_OUT_5_port, Y(4) => 
                           MUX2_OUT_4_port, Y(3) => MUX2_OUT_3_port, Y(2) => 
                           MUX2_OUT_2_port, Y(1) => MUX2_OUT_1_port, Y(0) => 
                           MUX2_OUT_0_port);
   ALUoutput : register_generic_nbits32_5 port map( data_in(31) => 
                           ALU_output_31_port, data_in(30) => 
                           ALU_output_30_port, data_in(29) => 
                           ALU_output_29_port, data_in(28) => 
                           ALU_output_28_port, data_in(27) => 
                           ALU_output_27_port, data_in(26) => 
                           ALU_output_26_port, data_in(25) => 
                           ALU_output_25_port, data_in(24) => 
                           ALU_output_24_port, data_in(23) => 
                           ALU_output_23_port, data_in(22) => 
                           ALU_output_22_port, data_in(21) => 
                           ALU_output_21_port, data_in(20) => 
                           ALU_output_20_port, data_in(19) => 
                           ALU_output_19_port, data_in(18) => 
                           ALU_output_18_port, data_in(17) => 
                           ALU_output_17_port, data_in(16) => 
                           ALU_output_16_port, data_in(15) => 
                           ALU_output_15_port, data_in(14) => 
                           ALU_output_14_port, data_in(13) => 
                           ALU_output_13_port, data_in(12) => 
                           ALU_output_12_port, data_in(11) => 
                           ALU_output_11_port, data_in(10) => 
                           ALU_output_10_port, data_in(9) => ALU_output_9_port,
                           data_in(8) => ALU_output_8_port, data_in(7) => 
                           ALU_output_7_port, data_in(6) => ALU_output_6_port, 
                           data_in(5) => ALU_output_5_port, data_in(4) => 
                           ALU_output_4_port, data_in(3) => ALU_output_3_port, 
                           data_in(2) => ALU_output_2_port, data_in(1) => 
                           ALU_output_1_port, data_in(0) => ALU_output_0_port, 
                           CK => n4, RESET => n3, ENABLE => ALU_OUTREG_ENABLE, 
                           data_out(31) => ALUREG_OUTPUT(31), data_out(30) => 
                           ALUREG_OUTPUT(30), data_out(29) => ALUREG_OUTPUT(29)
                           , data_out(28) => ALUREG_OUTPUT(28), data_out(27) =>
                           ALUREG_OUTPUT(27), data_out(26) => ALUREG_OUTPUT(26)
                           , data_out(25) => ALUREG_OUTPUT(25), data_out(24) =>
                           ALUREG_OUTPUT(24), data_out(23) => ALUREG_OUTPUT(23)
                           , data_out(22) => ALUREG_OUTPUT(22), data_out(21) =>
                           ALUREG_OUTPUT(21), data_out(20) => ALUREG_OUTPUT(20)
                           , data_out(19) => ALUREG_OUTPUT(19), data_out(18) =>
                           ALUREG_OUTPUT(18), data_out(17) => ALUREG_OUTPUT(17)
                           , data_out(16) => ALUREG_OUTPUT(16), data_out(15) =>
                           ALUREG_OUTPUT(15), data_out(14) => ALUREG_OUTPUT(14)
                           , data_out(13) => ALUREG_OUTPUT(13), data_out(12) =>
                           ALUREG_OUTPUT(12), data_out(11) => ALUREG_OUTPUT(11)
                           , data_out(10) => ALUREG_OUTPUT(10), data_out(9) => 
                           ALUREG_OUTPUT(9), data_out(8) => ALUREG_OUTPUT(8), 
                           data_out(7) => ALUREG_OUTPUT(7), data_out(6) => 
                           ALUREG_OUTPUT(6), data_out(5) => ALUREG_OUTPUT(5), 
                           data_out(4) => ALUREG_OUTPUT(4), data_out(3) => 
                           ALUREG_OUTPUT(3), data_out(2) => ALUREG_OUTPUT(2), 
                           data_out(1) => ALUREG_OUTPUT(1), data_out(0) => 
                           ALUREG_OUTPUT(0));
   IR3 : register_generic_nbits32_4 port map( data_in(31) => IR_IN3(31), 
                           data_in(30) => IR_IN3(30), data_in(29) => IR_IN3(29)
                           , data_in(28) => IR_IN3(28), data_in(27) => 
                           IR_IN3(27), data_in(26) => IR_IN3(26), data_in(25) 
                           => IR_IN3(25), data_in(24) => IR_IN3(24), 
                           data_in(23) => IR_IN3(23), data_in(22) => IR_IN3(22)
                           , data_in(21) => IR_IN3(21), data_in(20) => 
                           IR_IN3(20), data_in(19) => IR_IN3(19), data_in(18) 
                           => IR_IN3(18), data_in(17) => IR_IN3(17), 
                           data_in(16) => IR_IN3(16), data_in(15) => IR_IN3(15)
                           , data_in(14) => IR_IN3(14), data_in(13) => 
                           IR_IN3(13), data_in(12) => IR_IN3(12), data_in(11) 
                           => IR_IN3(11), data_in(10) => IR_IN3(10), data_in(9)
                           => IR_IN3(9), data_in(8) => IR_IN3(8), data_in(7) =>
                           IR_IN3(7), data_in(6) => IR_IN3(6), data_in(5) => 
                           IR_IN3(5), data_in(4) => IR_IN3(4), data_in(3) => 
                           IR_IN3(3), data_in(2) => IR_IN3(2), data_in(1) => 
                           IR_IN3(1), data_in(0) => IR_IN3(0), CK => n4, RESET 
                           => n3, ENABLE => X_Logic1_port, data_out(31) => 
                           IR_OUT3(31), data_out(30) => IR_OUT3(30), 
                           data_out(29) => IR_OUT3(29), data_out(28) => 
                           IR_OUT3(28), data_out(27) => IR_OUT3(27), 
                           data_out(26) => IR_OUT3(26), data_out(25) => 
                           IR_OUT3(25), data_out(24) => IR_OUT3(24), 
                           data_out(23) => IR_OUT3(23), data_out(22) => 
                           IR_OUT3(22), data_out(21) => IR_OUT3(21), 
                           data_out(20) => IR_OUT3(20), data_out(19) => 
                           IR_OUT3(19), data_out(18) => IR_OUT3(18), 
                           data_out(17) => IR_OUT3(17), data_out(16) => 
                           IR_OUT3(16), data_out(15) => IR_OUT3(15), 
                           data_out(14) => IR_OUT3(14), data_out(13) => 
                           IR_OUT3(13), data_out(12) => IR_OUT3(12), 
                           data_out(11) => IR_OUT3(11), data_out(10) => 
                           IR_OUT3(10), data_out(9) => IR_OUT3(9), data_out(8) 
                           => IR_OUT3(8), data_out(7) => IR_OUT3(7), 
                           data_out(6) => IR_OUT3(6), data_out(5) => IR_OUT3(5)
                           , data_out(4) => IR_OUT3(4), data_out(3) => 
                           IR_OUT3(3), data_out(2) => IR_OUT3(2), data_out(1) 
                           => IR_OUT3(1), data_out(0) => IR_OUT3(0));
   B_outregister : register_generic_nbits32_3 port map( data_in(31) => 
                           B_out(31), data_in(30) => B_out(30), data_in(29) => 
                           B_out(29), data_in(28) => B_out(28), data_in(27) => 
                           B_out(27), data_in(26) => B_out(26), data_in(25) => 
                           B_out(25), data_in(24) => B_out(24), data_in(23) => 
                           B_out(23), data_in(22) => B_out(22), data_in(21) => 
                           B_out(21), data_in(20) => B_out(20), data_in(19) => 
                           B_out(19), data_in(18) => B_out(18), data_in(17) => 
                           B_out(17), data_in(16) => B_out(16), data_in(15) => 
                           B_out(15), data_in(14) => B_out(14), data_in(13) => 
                           B_out(13), data_in(12) => B_out(12), data_in(11) => 
                           B_out(11), data_in(10) => B_out(10), data_in(9) => 
                           B_out(9), data_in(8) => B_out(8), data_in(7) => 
                           B_out(7), data_in(6) => B_out(6), data_in(5) => 
                           B_out(5), data_in(4) => B_out(4), data_in(3) => 
                           B_out(3), data_in(2) => B_out(2), data_in(1) => 
                           B_out(1), data_in(0) => B_out(0), CK => n4, RESET =>
                           n3, ENABLE => X_Logic1_port, data_out(31) => 
                           B_outreg(31), data_out(30) => B_outreg(30), 
                           data_out(29) => B_outreg(29), data_out(28) => 
                           B_outreg(28), data_out(27) => B_outreg(27), 
                           data_out(26) => B_outreg(26), data_out(25) => 
                           B_outreg(25), data_out(24) => B_outreg(24), 
                           data_out(23) => B_outreg(23), data_out(22) => 
                           B_outreg(22), data_out(21) => B_outreg(21), 
                           data_out(20) => B_outreg(20), data_out(19) => 
                           B_outreg(19), data_out(18) => B_outreg(18), 
                           data_out(17) => B_outreg(17), data_out(16) => 
                           B_outreg(16), data_out(15) => B_outreg(15), 
                           data_out(14) => B_outreg(14), data_out(13) => 
                           B_outreg(13), data_out(12) => B_outreg(12), 
                           data_out(11) => B_outreg(11), data_out(10) => 
                           B_outreg(10), data_out(9) => B_outreg(9), 
                           data_out(8) => B_outreg(8), data_out(7) => 
                           B_outreg(7), data_out(6) => B_outreg(6), data_out(5)
                           => B_outreg(5), data_out(4) => B_outreg(4), 
                           data_out(3) => B_outreg(3), data_out(2) => 
                           B_outreg(2), data_out(1) => B_outreg(1), data_out(0)
                           => B_outreg(0));
   alu1 : alu_nbits32 port map( FUNC(0) => ALU_BITS(0), FUNC(1) => ALU_BITS(1),
                           FUNC(2) => ALU_BITS(2), FUNC(3) => ALU_BITS(3), 
                           A(31) => MUX1_OUT_31_port, A(30) => MUX1_OUT_30_port
                           , A(29) => MUX1_OUT_29_port, A(28) => 
                           MUX1_OUT_28_port, A(27) => MUX1_OUT_27_port, A(26) 
                           => MUX1_OUT_26_port, A(25) => MUX1_OUT_25_port, 
                           A(24) => MUX1_OUT_24_port, A(23) => MUX1_OUT_23_port
                           , A(22) => MUX1_OUT_22_port, A(21) => 
                           MUX1_OUT_21_port, A(20) => MUX1_OUT_20_port, A(19) 
                           => MUX1_OUT_19_port, A(18) => MUX1_OUT_18_port, 
                           A(17) => MUX1_OUT_17_port, A(16) => MUX1_OUT_16_port
                           , A(15) => MUX1_OUT_15_port, A(14) => 
                           MUX1_OUT_14_port, A(13) => MUX1_OUT_13_port, A(12) 
                           => MUX1_OUT_12_port, A(11) => MUX1_OUT_11_port, 
                           A(10) => MUX1_OUT_10_port, A(9) => MUX1_OUT_9_port, 
                           A(8) => MUX1_OUT_8_port, A(7) => MUX1_OUT_7_port, 
                           A(6) => MUX1_OUT_6_port, A(5) => MUX1_OUT_5_port, 
                           A(4) => MUX1_OUT_4_port, A(3) => MUX1_OUT_3_port, 
                           A(2) => MUX1_OUT_2_port, A(1) => MUX1_OUT_1_port, 
                           A(0) => MUX1_OUT_0_port, B(31) => MUX2_OUT_31_port, 
                           B(30) => MUX2_OUT_30_port, B(29) => MUX2_OUT_29_port
                           , B(28) => MUX2_OUT_28_port, B(27) => 
                           MUX2_OUT_27_port, B(26) => MUX2_OUT_26_port, B(25) 
                           => MUX2_OUT_25_port, B(24) => MUX2_OUT_24_port, 
                           B(23) => MUX2_OUT_23_port, B(22) => MUX2_OUT_22_port
                           , B(21) => MUX2_OUT_21_port, B(20) => 
                           MUX2_OUT_20_port, B(19) => MUX2_OUT_19_port, B(18) 
                           => MUX2_OUT_18_port, B(17) => MUX2_OUT_17_port, 
                           B(16) => MUX2_OUT_16_port, B(15) => MUX2_OUT_15_port
                           , B(14) => MUX2_OUT_14_port, B(13) => 
                           MUX2_OUT_13_port, B(12) => MUX2_OUT_12_port, B(11) 
                           => MUX2_OUT_11_port, B(10) => MUX2_OUT_10_port, B(9)
                           => MUX2_OUT_9_port, B(8) => MUX2_OUT_8_port, B(7) =>
                           MUX2_OUT_7_port, B(6) => MUX2_OUT_6_port, B(5) => 
                           MUX2_OUT_5_port, B(4) => MUX2_OUT_4_port, B(3) => 
                           MUX2_OUT_3_port, B(2) => MUX2_OUT_2_port, B(1) => 
                           MUX2_OUT_1_port, B(0) => MUX2_OUT_0_port, OUTALU(31)
                           => ALU_output_31_port, OUTALU(30) => 
                           ALU_output_30_port, OUTALU(29) => ALU_output_29_port
                           , OUTALU(28) => ALU_output_28_port, OUTALU(27) => 
                           ALU_output_27_port, OUTALU(26) => ALU_output_26_port
                           , OUTALU(25) => ALU_output_25_port, OUTALU(24) => 
                           ALU_output_24_port, OUTALU(23) => ALU_output_23_port
                           , OUTALU(22) => ALU_output_22_port, OUTALU(21) => 
                           ALU_output_21_port, OUTALU(20) => ALU_output_20_port
                           , OUTALU(19) => ALU_output_19_port, OUTALU(18) => 
                           ALU_output_18_port, OUTALU(17) => ALU_output_17_port
                           , OUTALU(16) => ALU_output_16_port, OUTALU(15) => 
                           ALU_output_15_port, OUTALU(14) => ALU_output_14_port
                           , OUTALU(13) => ALU_output_13_port, OUTALU(12) => 
                           ALU_output_12_port, OUTALU(11) => ALU_output_11_port
                           , OUTALU(10) => ALU_output_10_port, OUTALU(9) => 
                           ALU_output_9_port, OUTALU(8) => ALU_output_8_port, 
                           OUTALU(7) => ALU_output_7_port, OUTALU(6) => 
                           ALU_output_6_port, OUTALU(5) => ALU_output_5_port, 
                           OUTALU(4) => ALU_output_4_port, OUTALU(3) => 
                           ALU_output_3_port, OUTALU(2) => ALU_output_2_port, 
                           OUTALU(1) => ALU_output_1_port, OUTALU(0) => 
                           ALU_output_0_port);
   XNOR_2 : XNOR_logic port map( A => ZERO_DEC_OUT, B => COND_ENABLE, Y => 
                           XNOR_OUT);
   COND : FD_0 port map( D => XNOR_OUT, CK => n4, RESET => n3, ENABLE => 
                           X_Logic1_port, Q => COND_OUT);
   U2 : BUF_X1 port map( A => rst, Z => n3);
   U3 : BUF_X1 port map( A => clk, Z => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity decodeUnit_nbits32 is

   port( clk, rst, RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE : in 
         std_logic;  DATAIN, IR_OUT : in std_logic_vector (31 downto 0);  A_out
         , B_out, Imm_out : out std_logic_vector (31 downto 0);  IR_IN2 : in 
         std_logic_vector (31 downto 0);  IR_OUT2 : out std_logic_vector (31 
         downto 0);  NPC_IN : in std_logic_vector (31 downto 0);  NPC2_OUT : 
         out std_logic_vector (31 downto 0));

end decodeUnit_nbits32;

architecture SYN_STRUCTURAL of decodeUnit_nbits32 is

   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component REGISTER_FILE_NBITS32_NREGISTERS32
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component SIGN_EXT_bits16
      port( inputt : in std_logic_vector (15 downto 0);  outputt : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_6
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_7
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_8
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, signExtOut_31_port, signExtOut_30_port, 
      signExtOut_29_port, signExtOut_28_port, signExtOut_27_port, 
      signExtOut_26_port, signExtOut_25_port, signExtOut_24_port, 
      signExtOut_23_port, signExtOut_22_port, signExtOut_21_port, 
      signExtOut_20_port, signExtOut_19_port, signExtOut_18_port, 
      signExtOut_17_port, signExtOut_16_port, signExtOut_15_port, 
      signExtOut_14_port, signExtOut_13_port, signExtOut_12_port, 
      signExtOut_11_port, signExtOut_10_port, signExtOut_9_port, 
      signExtOut_8_port, signExtOut_7_port, signExtOut_6_port, 
      signExtOut_5_port, signExtOut_4_port, signExtOut_3_port, 
      signExtOut_2_port, signExtOut_1_port, signExtOut_0_port, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18 : std_logic;

begin
   
   X_Logic1_port <= '1';
   NPC2 : register_generic_nbits32_8 port map( data_in(31) => NPC_IN(31), 
                           data_in(30) => NPC_IN(30), data_in(29) => NPC_IN(29)
                           , data_in(28) => NPC_IN(28), data_in(27) => 
                           NPC_IN(27), data_in(26) => NPC_IN(26), data_in(25) 
                           => NPC_IN(25), data_in(24) => NPC_IN(24), 
                           data_in(23) => NPC_IN(23), data_in(22) => NPC_IN(22)
                           , data_in(21) => NPC_IN(21), data_in(20) => 
                           NPC_IN(20), data_in(19) => NPC_IN(19), data_in(18) 
                           => NPC_IN(18), data_in(17) => NPC_IN(17), 
                           data_in(16) => NPC_IN(16), data_in(15) => NPC_IN(15)
                           , data_in(14) => NPC_IN(14), data_in(13) => 
                           NPC_IN(13), data_in(12) => NPC_IN(12), data_in(11) 
                           => NPC_IN(11), data_in(10) => NPC_IN(10), data_in(9)
                           => NPC_IN(9), data_in(8) => NPC_IN(8), data_in(7) =>
                           NPC_IN(7), data_in(6) => NPC_IN(6), data_in(5) => 
                           NPC_IN(5), data_in(4) => NPC_IN(4), data_in(3) => 
                           NPC_IN(3), data_in(2) => NPC_IN(2), data_in(1) => 
                           NPC_IN(1), data_in(0) => NPC_IN(0), CK => n11, RESET
                           => n10, ENABLE => X_Logic1_port, data_out(31) => 
                           NPC2_OUT(31), data_out(30) => NPC2_OUT(30), 
                           data_out(29) => NPC2_OUT(29), data_out(28) => 
                           NPC2_OUT(28), data_out(27) => NPC2_OUT(27), 
                           data_out(26) => NPC2_OUT(26), data_out(25) => 
                           NPC2_OUT(25), data_out(24) => NPC2_OUT(24), 
                           data_out(23) => NPC2_OUT(23), data_out(22) => 
                           NPC2_OUT(22), data_out(21) => NPC2_OUT(21), 
                           data_out(20) => NPC2_OUT(20), data_out(19) => 
                           NPC2_OUT(19), data_out(18) => NPC2_OUT(18), 
                           data_out(17) => NPC2_OUT(17), data_out(16) => 
                           NPC2_OUT(16), data_out(15) => NPC2_OUT(15), 
                           data_out(14) => NPC2_OUT(14), data_out(13) => 
                           NPC2_OUT(13), data_out(12) => NPC2_OUT(12), 
                           data_out(11) => NPC2_OUT(11), data_out(10) => 
                           NPC2_OUT(10), data_out(9) => NPC2_OUT(9), 
                           data_out(8) => NPC2_OUT(8), data_out(7) => 
                           NPC2_OUT(7), data_out(6) => NPC2_OUT(6), data_out(5)
                           => NPC2_OUT(5), data_out(4) => NPC2_OUT(4), 
                           data_out(3) => NPC2_OUT(3), data_out(2) => 
                           NPC2_OUT(2), data_out(1) => NPC2_OUT(1), data_out(0)
                           => NPC2_OUT(0));
   Imm : register_generic_nbits32_7 port map( data_in(31) => signExtOut_31_port
                           , data_in(30) => signExtOut_30_port, data_in(29) => 
                           signExtOut_29_port, data_in(28) => 
                           signExtOut_28_port, data_in(27) => 
                           signExtOut_27_port, data_in(26) => 
                           signExtOut_26_port, data_in(25) => 
                           signExtOut_25_port, data_in(24) => 
                           signExtOut_24_port, data_in(23) => 
                           signExtOut_23_port, data_in(22) => 
                           signExtOut_22_port, data_in(21) => 
                           signExtOut_21_port, data_in(20) => 
                           signExtOut_20_port, data_in(19) => 
                           signExtOut_19_port, data_in(18) => 
                           signExtOut_18_port, data_in(17) => 
                           signExtOut_17_port, data_in(16) => 
                           signExtOut_16_port, data_in(15) => 
                           signExtOut_15_port, data_in(14) => 
                           signExtOut_14_port, data_in(13) => 
                           signExtOut_13_port, data_in(12) => 
                           signExtOut_12_port, data_in(11) => 
                           signExtOut_11_port, data_in(10) => 
                           signExtOut_10_port, data_in(9) => signExtOut_9_port,
                           data_in(8) => signExtOut_8_port, data_in(7) => 
                           signExtOut_7_port, data_in(6) => signExtOut_6_port, 
                           data_in(5) => signExtOut_5_port, data_in(4) => 
                           signExtOut_4_port, data_in(3) => signExtOut_3_port, 
                           data_in(2) => signExtOut_2_port, data_in(1) => 
                           signExtOut_1_port, data_in(0) => signExtOut_0_port, 
                           CK => n11, RESET => n10, ENABLE => RegIMM_LATCH_EN, 
                           data_out(31) => Imm_out(31), data_out(30) => 
                           Imm_out(30), data_out(29) => Imm_out(29), 
                           data_out(28) => Imm_out(28), data_out(27) => 
                           Imm_out(27), data_out(26) => Imm_out(26), 
                           data_out(25) => Imm_out(25), data_out(24) => 
                           Imm_out(24), data_out(23) => Imm_out(23), 
                           data_out(22) => Imm_out(22), data_out(21) => 
                           Imm_out(21), data_out(20) => Imm_out(20), 
                           data_out(19) => Imm_out(19), data_out(18) => 
                           Imm_out(18), data_out(17) => Imm_out(17), 
                           data_out(16) => Imm_out(16), data_out(15) => 
                           Imm_out(15), data_out(14) => Imm_out(14), 
                           data_out(13) => Imm_out(13), data_out(12) => 
                           Imm_out(12), data_out(11) => Imm_out(11), 
                           data_out(10) => Imm_out(10), data_out(9) => 
                           Imm_out(9), data_out(8) => Imm_out(8), data_out(7) 
                           => Imm_out(7), data_out(6) => Imm_out(6), 
                           data_out(5) => Imm_out(5), data_out(4) => Imm_out(4)
                           , data_out(3) => Imm_out(3), data_out(2) => 
                           Imm_out(2), data_out(1) => Imm_out(1), data_out(0) 
                           => Imm_out(0));
   IR2 : register_generic_nbits32_6 port map( data_in(31) => IR_OUT(31), 
                           data_in(30) => IR_OUT(30), data_in(29) => IR_OUT(29)
                           , data_in(28) => IR_OUT(28), data_in(27) => 
                           IR_OUT(27), data_in(26) => IR_OUT(26), data_in(25) 
                           => IR_OUT(25), data_in(24) => IR_OUT(24), 
                           data_in(23) => IR_OUT(23), data_in(22) => IR_OUT(22)
                           , data_in(21) => IR_OUT(21), data_in(20) => 
                           IR_OUT(20), data_in(19) => IR_OUT(19), data_in(18) 
                           => IR_OUT(18), data_in(17) => IR_OUT(17), 
                           data_in(16) => IR_OUT(16), data_in(15) => IR_OUT(15)
                           , data_in(14) => IR_OUT(14), data_in(13) => 
                           IR_OUT(13), data_in(12) => IR_OUT(12), data_in(11) 
                           => IR_OUT(11), data_in(10) => IR_OUT(10), data_in(9)
                           => IR_OUT(9), data_in(8) => IR_OUT(8), data_in(7) =>
                           IR_OUT(7), data_in(6) => IR_OUT(6), data_in(5) => 
                           IR_OUT(5), data_in(4) => IR_OUT(4), data_in(3) => 
                           IR_OUT(3), data_in(2) => IR_OUT(2), data_in(1) => 
                           IR_OUT(1), data_in(0) => IR_OUT(0), CK => n11, RESET
                           => n10, ENABLE => X_Logic1_port, data_out(31) => 
                           IR_OUT2(31), data_out(30) => IR_OUT2(30), 
                           data_out(29) => IR_OUT2(29), data_out(28) => 
                           IR_OUT2(28), data_out(27) => IR_OUT2(27), 
                           data_out(26) => IR_OUT2(26), data_out(25) => 
                           IR_OUT2(25), data_out(24) => IR_OUT2(24), 
                           data_out(23) => IR_OUT2(23), data_out(22) => 
                           IR_OUT2(22), data_out(21) => IR_OUT2(21), 
                           data_out(20) => IR_OUT2(20), data_out(19) => 
                           IR_OUT2(19), data_out(18) => IR_OUT2(18), 
                           data_out(17) => IR_OUT2(17), data_out(16) => 
                           IR_OUT2(16), data_out(15) => IR_OUT2(15), 
                           data_out(14) => IR_OUT2(14), data_out(13) => 
                           IR_OUT2(13), data_out(12) => IR_OUT2(12), 
                           data_out(11) => IR_OUT2(11), data_out(10) => 
                           IR_OUT2(10), data_out(9) => IR_OUT2(9), data_out(8) 
                           => IR_OUT2(8), data_out(7) => IR_OUT2(7), 
                           data_out(6) => IR_OUT2(6), data_out(5) => IR_OUT2(5)
                           , data_out(4) => IR_OUT2(4), data_out(3) => 
                           IR_OUT2(3), data_out(2) => IR_OUT2(2), data_out(1) 
                           => IR_OUT2(1), data_out(0) => IR_OUT2(0));
   Signext : SIGN_EXT_bits16 port map( inputt(15) => IR_OUT(15), inputt(14) => 
                           IR_OUT(14), inputt(13) => IR_OUT(13), inputt(12) => 
                           IR_OUT(12), inputt(11) => IR_OUT(11), inputt(10) => 
                           IR_OUT(10), inputt(9) => IR_OUT(9), inputt(8) => 
                           IR_OUT(8), inputt(7) => IR_OUT(7), inputt(6) => 
                           IR_OUT(6), inputt(5) => IR_OUT(5), inputt(4) => 
                           IR_OUT(4), inputt(3) => IR_OUT(3), inputt(2) => 
                           IR_OUT(2), inputt(1) => IR_OUT(1), inputt(0) => 
                           IR_OUT(0), outputt(31) => signExtOut_31_port, 
                           outputt(30) => signExtOut_30_port, outputt(29) => 
                           signExtOut_29_port, outputt(28) => 
                           signExtOut_28_port, outputt(27) => 
                           signExtOut_27_port, outputt(26) => 
                           signExtOut_26_port, outputt(25) => 
                           signExtOut_25_port, outputt(24) => 
                           signExtOut_24_port, outputt(23) => 
                           signExtOut_23_port, outputt(22) => 
                           signExtOut_22_port, outputt(21) => 
                           signExtOut_21_port, outputt(20) => 
                           signExtOut_20_port, outputt(19) => 
                           signExtOut_19_port, outputt(18) => 
                           signExtOut_18_port, outputt(17) => 
                           signExtOut_17_port, outputt(16) => 
                           signExtOut_16_port, outputt(15) => 
                           signExtOut_15_port, outputt(14) => 
                           signExtOut_14_port, outputt(13) => 
                           signExtOut_13_port, outputt(12) => 
                           signExtOut_12_port, outputt(11) => 
                           signExtOut_11_port, outputt(10) => 
                           signExtOut_10_port, outputt(9) => signExtOut_9_port,
                           outputt(8) => signExtOut_8_port, outputt(7) => 
                           signExtOut_7_port, outputt(6) => signExtOut_6_port, 
                           outputt(5) => signExtOut_5_port, outputt(4) => 
                           signExtOut_4_port, outputt(3) => signExtOut_3_port, 
                           outputt(2) => signExtOut_2_port, outputt(1) => 
                           signExtOut_1_port, outputt(0) => signExtOut_0_port);
   RF : REGISTER_FILE_NBITS32_NREGISTERS32 port map( CLK => n11, RESET => n10, 
                           ENABLE => X_Logic1_port, RD1 => X_Logic1_port, RD2 
                           => X_Logic1_port, WR => RF_WE, ADD_WR(4) => n18, 
                           ADD_WR(3) => n17, ADD_WR(2) => n16, ADD_WR(1) => n15
                           , ADD_WR(0) => n14, ADD_RD1(4) => IR_OUT(25), 
                           ADD_RD1(3) => IR_OUT(24), ADD_RD1(2) => IR_OUT(23), 
                           ADD_RD1(1) => IR_OUT(22), ADD_RD1(0) => IR_OUT(21), 
                           ADD_RD2(4) => IR_OUT(20), ADD_RD2(3) => IR_OUT(19), 
                           ADD_RD2(2) => IR_OUT(18), ADD_RD2(1) => IR_OUT(17), 
                           ADD_RD2(0) => IR_OUT(16), DATAIN(31) => DATAIN(31), 
                           DATAIN(30) => DATAIN(30), DATAIN(29) => DATAIN(29), 
                           DATAIN(28) => DATAIN(28), DATAIN(27) => DATAIN(27), 
                           DATAIN(26) => DATAIN(26), DATAIN(25) => DATAIN(25), 
                           DATAIN(24) => DATAIN(24), DATAIN(23) => DATAIN(23), 
                           DATAIN(22) => DATAIN(22), DATAIN(21) => DATAIN(21), 
                           DATAIN(20) => DATAIN(20), DATAIN(19) => DATAIN(19), 
                           DATAIN(18) => DATAIN(18), DATAIN(17) => DATAIN(17), 
                           DATAIN(16) => DATAIN(16), DATAIN(15) => DATAIN(15), 
                           DATAIN(14) => DATAIN(14), DATAIN(13) => DATAIN(13), 
                           DATAIN(12) => DATAIN(12), DATAIN(11) => DATAIN(11), 
                           DATAIN(10) => DATAIN(10), DATAIN(9) => DATAIN(9), 
                           DATAIN(8) => DATAIN(8), DATAIN(7) => DATAIN(7), 
                           DATAIN(6) => DATAIN(6), DATAIN(5) => DATAIN(5), 
                           DATAIN(4) => DATAIN(4), DATAIN(3) => DATAIN(3), 
                           DATAIN(2) => DATAIN(2), DATAIN(1) => DATAIN(1), 
                           DATAIN(0) => DATAIN(0), OUT1(31) => A_out(31), 
                           OUT1(30) => A_out(30), OUT1(29) => A_out(29), 
                           OUT1(28) => A_out(28), OUT1(27) => A_out(27), 
                           OUT1(26) => A_out(26), OUT1(25) => A_out(25), 
                           OUT1(24) => A_out(24), OUT1(23) => A_out(23), 
                           OUT1(22) => A_out(22), OUT1(21) => A_out(21), 
                           OUT1(20) => A_out(20), OUT1(19) => A_out(19), 
                           OUT1(18) => A_out(18), OUT1(17) => A_out(17), 
                           OUT1(16) => A_out(16), OUT1(15) => A_out(15), 
                           OUT1(14) => A_out(14), OUT1(13) => A_out(13), 
                           OUT1(12) => A_out(12), OUT1(11) => A_out(11), 
                           OUT1(10) => A_out(10), OUT1(9) => A_out(9), OUT1(8) 
                           => A_out(8), OUT1(7) => A_out(7), OUT1(6) => 
                           A_out(6), OUT1(5) => A_out(5), OUT1(4) => A_out(4), 
                           OUT1(3) => A_out(3), OUT1(2) => A_out(2), OUT1(1) =>
                           A_out(1), OUT1(0) => A_out(0), OUT2(31) => B_out(31)
                           , OUT2(30) => B_out(30), OUT2(29) => B_out(29), 
                           OUT2(28) => B_out(28), OUT2(27) => B_out(27), 
                           OUT2(26) => B_out(26), OUT2(25) => B_out(25), 
                           OUT2(24) => B_out(24), OUT2(23) => B_out(23), 
                           OUT2(22) => B_out(22), OUT2(21) => B_out(21), 
                           OUT2(20) => B_out(20), OUT2(19) => B_out(19), 
                           OUT2(18) => B_out(18), OUT2(17) => B_out(17), 
                           OUT2(16) => B_out(16), OUT2(15) => B_out(15), 
                           OUT2(14) => B_out(14), OUT2(13) => B_out(13), 
                           OUT2(12) => B_out(12), OUT2(11) => B_out(11), 
                           OUT2(10) => B_out(10), OUT2(9) => B_out(9), OUT2(8) 
                           => B_out(8), OUT2(7) => B_out(7), OUT2(6) => 
                           B_out(6), OUT2(5) => B_out(5), OUT2(4) => B_out(4), 
                           OUT2(3) => B_out(3), OUT2(2) => B_out(2), OUT2(1) =>
                           B_out(1), OUT2(0) => B_out(0));
   U2 : NOR4_X2 port map( A1 => IR_IN2(28), A2 => IR_IN2(27), A3 => IR_IN2(26),
                           A4 => n13, ZN => n12);
   U3 : BUF_X1 port map( A => clk, Z => n11);
   U4 : BUF_X1 port map( A => rst, Z => n10);
   U5 : MUX2_X1 port map( A => IR_IN2(16), B => IR_IN2(11), S => n12, Z => n14)
                           ;
   U6 : MUX2_X1 port map( A => IR_IN2(17), B => IR_IN2(12), S => n12, Z => n15)
                           ;
   U7 : MUX2_X1 port map( A => IR_IN2(18), B => IR_IN2(13), S => n12, Z => n16)
                           ;
   U8 : MUX2_X1 port map( A => IR_IN2(19), B => IR_IN2(14), S => n12, Z => n17)
                           ;
   U9 : MUX2_X1 port map( A => IR_IN2(20), B => IR_IN2(15), S => n12, Z => n18)
                           ;
   U10 : OR3_X1 port map( A1 => IR_IN2(31), A2 => IR_IN2(30), A3 => IR_IN2(29),
                           ZN => n13);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity fetchUnit_nbits32 is

   port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 downto 
         0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN : in std_logic;  PC_IN : 
         in std_logic_vector (31 downto 0);  ADDRESS_IRAM, NPC_OUT, IR_OUT, 
         ADDERPC_OUT : out std_logic_vector (31 downto 0));

end fetchUnit_nbits32;

architecture SYN_STRUCTURAL of fetchUnit_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component register_generic_nbits32_9
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_10
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component register_generic_nbits32_0
      port( data_in : in std_logic_vector (31 downto 0);  CK, RESET, ENABLE : 
            in std_logic;  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component RCA_NBITS32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ADDRESS_IRAM_31_port, 
      ADDRESS_IRAM_30_port, ADDRESS_IRAM_29_port, ADDRESS_IRAM_28_port, 
      ADDRESS_IRAM_27_port, ADDRESS_IRAM_26_port, ADDRESS_IRAM_25_port, 
      ADDRESS_IRAM_24_port, ADDRESS_IRAM_23_port, ADDRESS_IRAM_22_port, 
      ADDRESS_IRAM_21_port, ADDRESS_IRAM_20_port, ADDRESS_IRAM_19_port, 
      ADDRESS_IRAM_18_port, ADDRESS_IRAM_17_port, ADDRESS_IRAM_16_port, 
      ADDRESS_IRAM_15_port, ADDRESS_IRAM_14_port, ADDRESS_IRAM_13_port, 
      ADDRESS_IRAM_12_port, ADDRESS_IRAM_11_port, ADDRESS_IRAM_10_port, 
      ADDRESS_IRAM_9_port, ADDRESS_IRAM_8_port, ADDRESS_IRAM_7_port, 
      ADDRESS_IRAM_6_port, ADDRESS_IRAM_5_port, ADDRESS_IRAM_4_port, 
      ADDRESS_IRAM_3_port, ADDRESS_IRAM_2_port, ADDRESS_IRAM_1_port, 
      ADDRESS_IRAM_0_port, ADDERPC_OUT_31_port, ADDERPC_OUT_30_port, 
      ADDERPC_OUT_29_port, ADDERPC_OUT_28_port, ADDERPC_OUT_27_port, 
      ADDERPC_OUT_26_port, ADDERPC_OUT_25_port, ADDERPC_OUT_24_port, 
      ADDERPC_OUT_23_port, ADDERPC_OUT_22_port, ADDERPC_OUT_21_port, 
      ADDERPC_OUT_20_port, ADDERPC_OUT_19_port, ADDERPC_OUT_18_port, 
      ADDERPC_OUT_17_port, ADDERPC_OUT_16_port, ADDERPC_OUT_15_port, 
      ADDERPC_OUT_14_port, ADDERPC_OUT_13_port, ADDERPC_OUT_12_port, 
      ADDERPC_OUT_11_port, ADDERPC_OUT_10_port, ADDERPC_OUT_9_port, 
      ADDERPC_OUT_8_port, ADDERPC_OUT_7_port, ADDERPC_OUT_6_port, 
      ADDERPC_OUT_5_port, ADDERPC_OUT_4_port, ADDERPC_OUT_3_port, 
      ADDERPC_OUT_2_port, ADDERPC_OUT_1_port, ADDERPC_OUT_0_port, n3, n4, 
      n_2044 : std_logic;

begin
   ADDRESS_IRAM <= ( ADDRESS_IRAM_31_port, ADDRESS_IRAM_30_port, 
      ADDRESS_IRAM_29_port, ADDRESS_IRAM_28_port, ADDRESS_IRAM_27_port, 
      ADDRESS_IRAM_26_port, ADDRESS_IRAM_25_port, ADDRESS_IRAM_24_port, 
      ADDRESS_IRAM_23_port, ADDRESS_IRAM_22_port, ADDRESS_IRAM_21_port, 
      ADDRESS_IRAM_20_port, ADDRESS_IRAM_19_port, ADDRESS_IRAM_18_port, 
      ADDRESS_IRAM_17_port, ADDRESS_IRAM_16_port, ADDRESS_IRAM_15_port, 
      ADDRESS_IRAM_14_port, ADDRESS_IRAM_13_port, ADDRESS_IRAM_12_port, 
      ADDRESS_IRAM_11_port, ADDRESS_IRAM_10_port, ADDRESS_IRAM_9_port, 
      ADDRESS_IRAM_8_port, ADDRESS_IRAM_7_port, ADDRESS_IRAM_6_port, 
      ADDRESS_IRAM_5_port, ADDRESS_IRAM_4_port, ADDRESS_IRAM_3_port, 
      ADDRESS_IRAM_2_port, ADDRESS_IRAM_1_port, ADDRESS_IRAM_0_port );
   ADDERPC_OUT <= ( ADDERPC_OUT_31_port, ADDERPC_OUT_30_port, 
      ADDERPC_OUT_29_port, ADDERPC_OUT_28_port, ADDERPC_OUT_27_port, 
      ADDERPC_OUT_26_port, ADDERPC_OUT_25_port, ADDERPC_OUT_24_port, 
      ADDERPC_OUT_23_port, ADDERPC_OUT_22_port, ADDERPC_OUT_21_port, 
      ADDERPC_OUT_20_port, ADDERPC_OUT_19_port, ADDERPC_OUT_18_port, 
      ADDERPC_OUT_17_port, ADDERPC_OUT_16_port, ADDERPC_OUT_15_port, 
      ADDERPC_OUT_14_port, ADDERPC_OUT_13_port, ADDERPC_OUT_12_port, 
      ADDERPC_OUT_11_port, ADDERPC_OUT_10_port, ADDERPC_OUT_9_port, 
      ADDERPC_OUT_8_port, ADDERPC_OUT_7_port, ADDERPC_OUT_6_port, 
      ADDERPC_OUT_5_port, ADDERPC_OUT_4_port, ADDERPC_OUT_3_port, 
      ADDERPC_OUT_2_port, ADDERPC_OUT_1_port, ADDERPC_OUT_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADD : RCA_NBITS32 port map( A(31) => ADDRESS_IRAM_31_port, A(30) => 
                           ADDRESS_IRAM_30_port, A(29) => ADDRESS_IRAM_29_port,
                           A(28) => ADDRESS_IRAM_28_port, A(27) => 
                           ADDRESS_IRAM_27_port, A(26) => ADDRESS_IRAM_26_port,
                           A(25) => ADDRESS_IRAM_25_port, A(24) => 
                           ADDRESS_IRAM_24_port, A(23) => ADDRESS_IRAM_23_port,
                           A(22) => ADDRESS_IRAM_22_port, A(21) => 
                           ADDRESS_IRAM_21_port, A(20) => ADDRESS_IRAM_20_port,
                           A(19) => ADDRESS_IRAM_19_port, A(18) => 
                           ADDRESS_IRAM_18_port, A(17) => ADDRESS_IRAM_17_port,
                           A(16) => ADDRESS_IRAM_16_port, A(15) => 
                           ADDRESS_IRAM_15_port, A(14) => ADDRESS_IRAM_14_port,
                           A(13) => ADDRESS_IRAM_13_port, A(12) => 
                           ADDRESS_IRAM_12_port, A(11) => ADDRESS_IRAM_11_port,
                           A(10) => ADDRESS_IRAM_10_port, A(9) => 
                           ADDRESS_IRAM_9_port, A(8) => ADDRESS_IRAM_8_port, 
                           A(7) => ADDRESS_IRAM_7_port, A(6) => 
                           ADDRESS_IRAM_6_port, A(5) => ADDRESS_IRAM_5_port, 
                           A(4) => ADDRESS_IRAM_4_port, A(3) => 
                           ADDRESS_IRAM_3_port, A(2) => ADDRESS_IRAM_2_port, 
                           A(1) => ADDRESS_IRAM_1_port, A(0) => 
                           ADDRESS_IRAM_0_port, B(31) => X_Logic0_port, B(30) 
                           => X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic1_port, Ci => X_Logic0_port, S(31) => 
                           ADDERPC_OUT_31_port, S(30) => ADDERPC_OUT_30_port, 
                           S(29) => ADDERPC_OUT_29_port, S(28) => 
                           ADDERPC_OUT_28_port, S(27) => ADDERPC_OUT_27_port, 
                           S(26) => ADDERPC_OUT_26_port, S(25) => 
                           ADDERPC_OUT_25_port, S(24) => ADDERPC_OUT_24_port, 
                           S(23) => ADDERPC_OUT_23_port, S(22) => 
                           ADDERPC_OUT_22_port, S(21) => ADDERPC_OUT_21_port, 
                           S(20) => ADDERPC_OUT_20_port, S(19) => 
                           ADDERPC_OUT_19_port, S(18) => ADDERPC_OUT_18_port, 
                           S(17) => ADDERPC_OUT_17_port, S(16) => 
                           ADDERPC_OUT_16_port, S(15) => ADDERPC_OUT_15_port, 
                           S(14) => ADDERPC_OUT_14_port, S(13) => 
                           ADDERPC_OUT_13_port, S(12) => ADDERPC_OUT_12_port, 
                           S(11) => ADDERPC_OUT_11_port, S(10) => 
                           ADDERPC_OUT_10_port, S(9) => ADDERPC_OUT_9_port, 
                           S(8) => ADDERPC_OUT_8_port, S(7) => 
                           ADDERPC_OUT_7_port, S(6) => ADDERPC_OUT_6_port, S(5)
                           => ADDERPC_OUT_5_port, S(4) => ADDERPC_OUT_4_port, 
                           S(3) => ADDERPC_OUT_3_port, S(2) => 
                           ADDERPC_OUT_2_port, S(1) => ADDERPC_OUT_1_port, S(0)
                           => ADDERPC_OUT_0_port, Co => n_2044);
   PC : register_generic_nbits32_0 port map( data_in(31) => PC_IN(31), 
                           data_in(30) => PC_IN(30), data_in(29) => PC_IN(29), 
                           data_in(28) => PC_IN(28), data_in(27) => PC_IN(27), 
                           data_in(26) => PC_IN(26), data_in(25) => PC_IN(25), 
                           data_in(24) => PC_IN(24), data_in(23) => PC_IN(23), 
                           data_in(22) => PC_IN(22), data_in(21) => PC_IN(21), 
                           data_in(20) => PC_IN(20), data_in(19) => PC_IN(19), 
                           data_in(18) => PC_IN(18), data_in(17) => PC_IN(17), 
                           data_in(16) => PC_IN(16), data_in(15) => PC_IN(15), 
                           data_in(14) => PC_IN(14), data_in(13) => PC_IN(13), 
                           data_in(12) => PC_IN(12), data_in(11) => PC_IN(11), 
                           data_in(10) => PC_IN(10), data_in(9) => PC_IN(9), 
                           data_in(8) => PC_IN(8), data_in(7) => PC_IN(7), 
                           data_in(6) => PC_IN(6), data_in(5) => PC_IN(5), 
                           data_in(4) => PC_IN(4), data_in(3) => PC_IN(3), 
                           data_in(2) => PC_IN(2), data_in(1) => PC_IN(1), 
                           data_in(0) => PC_IN(0), CK => n4, RESET => n3, 
                           ENABLE => PC_LATCH_EN, data_out(31) => 
                           ADDRESS_IRAM_31_port, data_out(30) => 
                           ADDRESS_IRAM_30_port, data_out(29) => 
                           ADDRESS_IRAM_29_port, data_out(28) => 
                           ADDRESS_IRAM_28_port, data_out(27) => 
                           ADDRESS_IRAM_27_port, data_out(26) => 
                           ADDRESS_IRAM_26_port, data_out(25) => 
                           ADDRESS_IRAM_25_port, data_out(24) => 
                           ADDRESS_IRAM_24_port, data_out(23) => 
                           ADDRESS_IRAM_23_port, data_out(22) => 
                           ADDRESS_IRAM_22_port, data_out(21) => 
                           ADDRESS_IRAM_21_port, data_out(20) => 
                           ADDRESS_IRAM_20_port, data_out(19) => 
                           ADDRESS_IRAM_19_port, data_out(18) => 
                           ADDRESS_IRAM_18_port, data_out(17) => 
                           ADDRESS_IRAM_17_port, data_out(16) => 
                           ADDRESS_IRAM_16_port, data_out(15) => 
                           ADDRESS_IRAM_15_port, data_out(14) => 
                           ADDRESS_IRAM_14_port, data_out(13) => 
                           ADDRESS_IRAM_13_port, data_out(12) => 
                           ADDRESS_IRAM_12_port, data_out(11) => 
                           ADDRESS_IRAM_11_port, data_out(10) => 
                           ADDRESS_IRAM_10_port, data_out(9) => 
                           ADDRESS_IRAM_9_port, data_out(8) => 
                           ADDRESS_IRAM_8_port, data_out(7) => 
                           ADDRESS_IRAM_7_port, data_out(6) => 
                           ADDRESS_IRAM_6_port, data_out(5) => 
                           ADDRESS_IRAM_5_port, data_out(4) => 
                           ADDRESS_IRAM_4_port, data_out(3) => 
                           ADDRESS_IRAM_3_port, data_out(2) => 
                           ADDRESS_IRAM_2_port, data_out(1) => 
                           ADDRESS_IRAM_1_port, data_out(0) => 
                           ADDRESS_IRAM_0_port);
   IR : register_generic_nbits32_10 port map( data_in(31) => DATA_IRAM(31), 
                           data_in(30) => DATA_IRAM(30), data_in(29) => 
                           DATA_IRAM(29), data_in(28) => DATA_IRAM(28), 
                           data_in(27) => DATA_IRAM(27), data_in(26) => 
                           DATA_IRAM(26), data_in(25) => DATA_IRAM(25), 
                           data_in(24) => DATA_IRAM(24), data_in(23) => 
                           DATA_IRAM(23), data_in(22) => DATA_IRAM(22), 
                           data_in(21) => DATA_IRAM(21), data_in(20) => 
                           DATA_IRAM(20), data_in(19) => DATA_IRAM(19), 
                           data_in(18) => DATA_IRAM(18), data_in(17) => 
                           DATA_IRAM(17), data_in(16) => DATA_IRAM(16), 
                           data_in(15) => DATA_IRAM(15), data_in(14) => 
                           DATA_IRAM(14), data_in(13) => DATA_IRAM(13), 
                           data_in(12) => DATA_IRAM(12), data_in(11) => 
                           DATA_IRAM(11), data_in(10) => DATA_IRAM(10), 
                           data_in(9) => DATA_IRAM(9), data_in(8) => 
                           DATA_IRAM(8), data_in(7) => DATA_IRAM(7), data_in(6)
                           => DATA_IRAM(6), data_in(5) => DATA_IRAM(5), 
                           data_in(4) => DATA_IRAM(4), data_in(3) => 
                           DATA_IRAM(3), data_in(2) => DATA_IRAM(2), data_in(1)
                           => DATA_IRAM(1), data_in(0) => DATA_IRAM(0), CK => 
                           n4, RESET => n3, ENABLE => IR_LATCH_EN, data_out(31)
                           => IR_OUT(31), data_out(30) => IR_OUT(30), 
                           data_out(29) => IR_OUT(29), data_out(28) => 
                           IR_OUT(28), data_out(27) => IR_OUT(27), data_out(26)
                           => IR_OUT(26), data_out(25) => IR_OUT(25), 
                           data_out(24) => IR_OUT(24), data_out(23) => 
                           IR_OUT(23), data_out(22) => IR_OUT(22), data_out(21)
                           => IR_OUT(21), data_out(20) => IR_OUT(20), 
                           data_out(19) => IR_OUT(19), data_out(18) => 
                           IR_OUT(18), data_out(17) => IR_OUT(17), data_out(16)
                           => IR_OUT(16), data_out(15) => IR_OUT(15), 
                           data_out(14) => IR_OUT(14), data_out(13) => 
                           IR_OUT(13), data_out(12) => IR_OUT(12), data_out(11)
                           => IR_OUT(11), data_out(10) => IR_OUT(10), 
                           data_out(9) => IR_OUT(9), data_out(8) => IR_OUT(8), 
                           data_out(7) => IR_OUT(7), data_out(6) => IR_OUT(6), 
                           data_out(5) => IR_OUT(5), data_out(4) => IR_OUT(4), 
                           data_out(3) => IR_OUT(3), data_out(2) => IR_OUT(2), 
                           data_out(1) => IR_OUT(1), data_out(0) => IR_OUT(0));
   NPC : register_generic_nbits32_9 port map( data_in(31) => 
                           ADDERPC_OUT_31_port, data_in(30) => 
                           ADDERPC_OUT_30_port, data_in(29) => 
                           ADDERPC_OUT_29_port, data_in(28) => 
                           ADDERPC_OUT_28_port, data_in(27) => 
                           ADDERPC_OUT_27_port, data_in(26) => 
                           ADDERPC_OUT_26_port, data_in(25) => 
                           ADDERPC_OUT_25_port, data_in(24) => 
                           ADDERPC_OUT_24_port, data_in(23) => 
                           ADDERPC_OUT_23_port, data_in(22) => 
                           ADDERPC_OUT_22_port, data_in(21) => 
                           ADDERPC_OUT_21_port, data_in(20) => 
                           ADDERPC_OUT_20_port, data_in(19) => 
                           ADDERPC_OUT_19_port, data_in(18) => 
                           ADDERPC_OUT_18_port, data_in(17) => 
                           ADDERPC_OUT_17_port, data_in(16) => 
                           ADDERPC_OUT_16_port, data_in(15) => 
                           ADDERPC_OUT_15_port, data_in(14) => 
                           ADDERPC_OUT_14_port, data_in(13) => 
                           ADDERPC_OUT_13_port, data_in(12) => 
                           ADDERPC_OUT_12_port, data_in(11) => 
                           ADDERPC_OUT_11_port, data_in(10) => 
                           ADDERPC_OUT_10_port, data_in(9) => 
                           ADDERPC_OUT_9_port, data_in(8) => ADDERPC_OUT_8_port
                           , data_in(7) => ADDERPC_OUT_7_port, data_in(6) => 
                           ADDERPC_OUT_6_port, data_in(5) => ADDERPC_OUT_5_port
                           , data_in(4) => ADDERPC_OUT_4_port, data_in(3) => 
                           ADDERPC_OUT_3_port, data_in(2) => ADDERPC_OUT_2_port
                           , data_in(1) => ADDERPC_OUT_1_port, data_in(0) => 
                           ADDERPC_OUT_0_port, CK => n4, RESET => n3, ENABLE =>
                           NPC_LATCH_EN, data_out(31) => NPC_OUT(31), 
                           data_out(30) => NPC_OUT(30), data_out(29) => 
                           NPC_OUT(29), data_out(28) => NPC_OUT(28), 
                           data_out(27) => NPC_OUT(27), data_out(26) => 
                           NPC_OUT(26), data_out(25) => NPC_OUT(25), 
                           data_out(24) => NPC_OUT(24), data_out(23) => 
                           NPC_OUT(23), data_out(22) => NPC_OUT(22), 
                           data_out(21) => NPC_OUT(21), data_out(20) => 
                           NPC_OUT(20), data_out(19) => NPC_OUT(19), 
                           data_out(18) => NPC_OUT(18), data_out(17) => 
                           NPC_OUT(17), data_out(16) => NPC_OUT(16), 
                           data_out(15) => NPC_OUT(15), data_out(14) => 
                           NPC_OUT(14), data_out(13) => NPC_OUT(13), 
                           data_out(12) => NPC_OUT(12), data_out(11) => 
                           NPC_OUT(11), data_out(10) => NPC_OUT(10), 
                           data_out(9) => NPC_OUT(9), data_out(8) => NPC_OUT(8)
                           , data_out(7) => NPC_OUT(7), data_out(6) => 
                           NPC_OUT(6), data_out(5) => NPC_OUT(5), data_out(4) 
                           => NPC_OUT(4), data_out(3) => NPC_OUT(3), 
                           data_out(2) => NPC_OUT(2), data_out(1) => NPC_OUT(1)
                           , data_out(0) => NPC_OUT(0));
   U3 : BUF_X1 port map( A => rst, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity datapath_nbits32 is

   port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 downto 
         0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN, RegA_LATCH_EN, 
         RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE, MUXA_SEL, MUXB_SEL, 
         ALU_OUTREG_EN, EQ_COND : in std_logic;  ALU_OPCODE : in 
         std_logic_vector (0 to 3);  DRAM_DATA : in std_logic_vector (31 downto
         0);  LMD_LATCH_EN, JUMP_EN, WB_MUX_SEL : in std_logic;  B, ALU_OUT, 
         ADDRESS_IRAM, IR_OUT : out std_logic_vector (31 downto 0));

end datapath_nbits32;

architecture SYN_STRUCTURAL of datapath_nbits32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component writeBack_nbits32
      port( LMD_OUT, ALUREG_OUTPUT : in std_logic_vector (31 downto 0);  
            WB_MUX_SEL : in std_logic;  DATAIN_RF : out std_logic_vector (31 
            downto 0));
   end component;
   
   component memoryUnit_nbits32
      port( clk, rst, LMD_LATCH_EN, JUMP_EN : in std_logic;  DRAM_DATA, 
            ALUREG_OUTPUT, NPC_OUT : in std_logic_vector (31 downto 0);  
            COND_OUT : in std_logic;  DRAM_DATAout, TO_PC_OUT, ALU_OUT2 : out 
            std_logic_vector (31 downto 0);  IR_IN4 : in std_logic_vector (31 
            downto 0);  IR_OUT4 : out std_logic_vector (31 downto 0));
   end component;
   
   component executionUnit_nbits32
      port( clk, rst, ALU_OUTREG_ENABLE, MUXA_SEL, MUXB_SEL, COND_ENABLE : in 
            std_logic;  ALU_BITS : in std_logic_vector (0 to 3);  NPC_OUT, 
            A_out, B_out, Imm_out : in std_logic_vector (31 downto 0);  
            ALUREG_OUTPUT : out std_logic_vector (31 downto 0);  COND_OUT : out
            std_logic;  IR_IN3 : in std_logic_vector (31 downto 0);  IR_OUT3, 
            B_outreg : out std_logic_vector (31 downto 0));
   end component;
   
   component decodeUnit_nbits32
      port( clk, rst, RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE : in
            std_logic;  DATAIN, IR_OUT : in std_logic_vector (31 downto 0);  
            A_out, B_out, Imm_out : out std_logic_vector (31 downto 0);  IR_IN2
            : in std_logic_vector (31 downto 0);  IR_OUT2 : out 
            std_logic_vector (31 downto 0);  NPC_IN : in std_logic_vector (31 
            downto 0);  NPC2_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component fetchUnit_nbits32
      port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 
            downto 0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN : in std_logic; 
            PC_IN : in std_logic_vector (31 downto 0);  ADDRESS_IRAM, NPC_OUT, 
            IR_OUT, ADDERPC_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal ALU_OUT_31_port, ALU_OUT_30_port, ALU_OUT_29_port, ALU_OUT_28_port, 
      ALU_OUT_27_port, ALU_OUT_26_port, ALU_OUT_25_port, ALU_OUT_24_port, 
      ALU_OUT_23_port, ALU_OUT_22_port, ALU_OUT_21_port, ALU_OUT_20_port, 
      ALU_OUT_19_port, ALU_OUT_18_port, ALU_OUT_17_port, ALU_OUT_16_port, 
      ALU_OUT_15_port, ALU_OUT_14_port, ALU_OUT_13_port, ALU_OUT_12_port, 
      ALU_OUT_11_port, ALU_OUT_10_port, ALU_OUT_9_port, ALU_OUT_8_port, 
      ALU_OUT_7_port, ALU_OUT_6_port, ALU_OUT_5_port, ALU_OUT_4_port, 
      ALU_OUT_3_port, ALU_OUT_2_port, ALU_OUT_1_port, ALU_OUT_0_port, 
      IR_OUT_31_port, IR_OUT_30_port, IR_OUT_29_port, IR_OUT_28_port, 
      IR_OUT_27_port, IR_OUT_26_port, IR_OUT_25_port, IR_OUT_24_port, 
      IR_OUT_23_port, IR_OUT_22_port, IR_OUT_21_port, IR_OUT_20_port, 
      IR_OUT_19_port, IR_OUT_18_port, IR_OUT_17_port, IR_OUT_16_port, 
      IR_OUT_15_port, IR_OUT_14_port, IR_OUT_13_port, IR_OUT_12_port, 
      IR_OUT_11_port, IR_OUT_10_port, IR_OUT_9_port, IR_OUT_8_port, 
      IR_OUT_7_port, IR_OUT_6_port, IR_OUT_5_port, IR_OUT_4_port, IR_OUT_3_port
      , IR_OUT_2_port, IR_OUT_1_port, IR_OUT_0_port, TO_PC_OUTs_31_port, 
      TO_PC_OUTs_30_port, TO_PC_OUTs_29_port, TO_PC_OUTs_28_port, 
      TO_PC_OUTs_27_port, TO_PC_OUTs_26_port, TO_PC_OUTs_25_port, 
      TO_PC_OUTs_24_port, TO_PC_OUTs_23_port, TO_PC_OUTs_22_port, 
      TO_PC_OUTs_21_port, TO_PC_OUTs_20_port, TO_PC_OUTs_19_port, 
      TO_PC_OUTs_18_port, TO_PC_OUTs_17_port, TO_PC_OUTs_16_port, 
      TO_PC_OUTs_15_port, TO_PC_OUTs_14_port, TO_PC_OUTs_13_port, 
      TO_PC_OUTs_12_port, TO_PC_OUTs_11_port, TO_PC_OUTs_10_port, 
      TO_PC_OUTs_9_port, TO_PC_OUTs_8_port, TO_PC_OUTs_7_port, 
      TO_PC_OUTs_6_port, TO_PC_OUTs_5_port, TO_PC_OUTs_4_port, 
      TO_PC_OUTs_3_port, TO_PC_OUTs_2_port, TO_PC_OUTs_1_port, 
      TO_PC_OUTs_0_port, NPC_OUTs_31_port, NPC_OUTs_30_port, NPC_OUTs_29_port, 
      NPC_OUTs_28_port, NPC_OUTs_27_port, NPC_OUTs_26_port, NPC_OUTs_25_port, 
      NPC_OUTs_24_port, NPC_OUTs_23_port, NPC_OUTs_22_port, NPC_OUTs_21_port, 
      NPC_OUTs_20_port, NPC_OUTs_19_port, NPC_OUTs_18_port, NPC_OUTs_17_port, 
      NPC_OUTs_16_port, NPC_OUTs_15_port, NPC_OUTs_14_port, NPC_OUTs_13_port, 
      NPC_OUTs_12_port, NPC_OUTs_11_port, NPC_OUTs_10_port, NPC_OUTs_9_port, 
      NPC_OUTs_8_port, NPC_OUTs_7_port, NPC_OUTs_6_port, NPC_OUTs_5_port, 
      NPC_OUTs_4_port, NPC_OUTs_3_port, NPC_OUTs_2_port, NPC_OUTs_1_port, 
      NPC_OUTs_0_port, ADDERPC_OUTs_31_port, ADDERPC_OUTs_30_port, 
      ADDERPC_OUTs_29_port, ADDERPC_OUTs_28_port, ADDERPC_OUTs_27_port, 
      ADDERPC_OUTs_26_port, ADDERPC_OUTs_25_port, ADDERPC_OUTs_24_port, 
      ADDERPC_OUTs_23_port, ADDERPC_OUTs_22_port, ADDERPC_OUTs_21_port, 
      ADDERPC_OUTs_20_port, ADDERPC_OUTs_19_port, ADDERPC_OUTs_18_port, 
      ADDERPC_OUTs_17_port, ADDERPC_OUTs_16_port, ADDERPC_OUTs_15_port, 
      ADDERPC_OUTs_14_port, ADDERPC_OUTs_13_port, ADDERPC_OUTs_12_port, 
      ADDERPC_OUTs_11_port, ADDERPC_OUTs_10_port, ADDERPC_OUTs_9_port, 
      ADDERPC_OUTs_8_port, ADDERPC_OUTs_7_port, ADDERPC_OUTs_6_port, 
      ADDERPC_OUTs_5_port, ADDERPC_OUTs_4_port, ADDERPC_OUTs_3_port, 
      ADDERPC_OUTs_2_port, ADDERPC_OUTs_1_port, ADDERPC_OUTs_0_port, 
      DATAIN_RFs_31_port, DATAIN_RFs_30_port, DATAIN_RFs_29_port, 
      DATAIN_RFs_28_port, DATAIN_RFs_27_port, DATAIN_RFs_26_port, 
      DATAIN_RFs_25_port, DATAIN_RFs_24_port, DATAIN_RFs_23_port, 
      DATAIN_RFs_22_port, DATAIN_RFs_21_port, DATAIN_RFs_20_port, 
      DATAIN_RFs_19_port, DATAIN_RFs_18_port, DATAIN_RFs_17_port, 
      DATAIN_RFs_16_port, DATAIN_RFs_15_port, DATAIN_RFs_14_port, 
      DATAIN_RFs_13_port, DATAIN_RFs_12_port, DATAIN_RFs_11_port, 
      DATAIN_RFs_10_port, DATAIN_RFs_9_port, DATAIN_RFs_8_port, 
      DATAIN_RFs_7_port, DATAIN_RFs_6_port, DATAIN_RFs_5_port, 
      DATAIN_RFs_4_port, DATAIN_RFs_3_port, DATAIN_RFs_2_port, 
      DATAIN_RFs_1_port, DATAIN_RFs_0_port, A_outs_31_port, A_outs_30_port, 
      A_outs_29_port, A_outs_28_port, A_outs_27_port, A_outs_26_port, 
      A_outs_25_port, A_outs_24_port, A_outs_23_port, A_outs_22_port, 
      A_outs_21_port, A_outs_20_port, A_outs_19_port, A_outs_18_port, 
      A_outs_17_port, A_outs_16_port, A_outs_15_port, A_outs_14_port, 
      A_outs_13_port, A_outs_12_port, A_outs_11_port, A_outs_10_port, 
      A_outs_9_port, A_outs_8_port, A_outs_7_port, A_outs_6_port, A_outs_5_port
      , A_outs_4_port, A_outs_3_port, A_outs_2_port, A_outs_1_port, 
      A_outs_0_port, B_outs_31_port, B_outs_30_port, B_outs_29_port, 
      B_outs_28_port, B_outs_27_port, B_outs_26_port, B_outs_25_port, 
      B_outs_24_port, B_outs_23_port, B_outs_22_port, B_outs_21_port, 
      B_outs_20_port, B_outs_19_port, B_outs_18_port, B_outs_17_port, 
      B_outs_16_port, B_outs_15_port, B_outs_14_port, B_outs_13_port, 
      B_outs_12_port, B_outs_11_port, B_outs_10_port, B_outs_9_port, 
      B_outs_8_port, B_outs_7_port, B_outs_6_port, B_outs_5_port, B_outs_4_port
      , B_outs_3_port, B_outs_2_port, B_outs_1_port, B_outs_0_port, 
      Imm_outs_31_port, Imm_outs_30_port, Imm_outs_29_port, Imm_outs_28_port, 
      Imm_outs_27_port, Imm_outs_26_port, Imm_outs_25_port, Imm_outs_24_port, 
      Imm_outs_23_port, Imm_outs_22_port, Imm_outs_21_port, Imm_outs_20_port, 
      Imm_outs_19_port, Imm_outs_18_port, Imm_outs_17_port, Imm_outs_16_port, 
      Imm_outs_15_port, Imm_outs_14_port, Imm_outs_13_port, Imm_outs_12_port, 
      Imm_outs_11_port, Imm_outs_10_port, Imm_outs_9_port, Imm_outs_8_port, 
      Imm_outs_7_port, Imm_outs_6_port, Imm_outs_5_port, Imm_outs_4_port, 
      Imm_outs_3_port, Imm_outs_2_port, Imm_outs_1_port, Imm_outs_0_port, 
      IR_OUT4s_31_port, IR_OUT4s_30_port, IR_OUT4s_29_port, IR_OUT4s_28_port, 
      IR_OUT4s_27_port, IR_OUT4s_26_port, IR_OUT4s_25_port, IR_OUT4s_24_port, 
      IR_OUT4s_23_port, IR_OUT4s_22_port, IR_OUT4s_21_port, IR_OUT4s_20_port, 
      IR_OUT4s_19_port, IR_OUT4s_18_port, IR_OUT4s_17_port, IR_OUT4s_16_port, 
      IR_OUT4s_15_port, IR_OUT4s_14_port, IR_OUT4s_13_port, IR_OUT4s_12_port, 
      IR_OUT4s_11_port, IR_OUT4s_10_port, IR_OUT4s_9_port, IR_OUT4s_8_port, 
      IR_OUT4s_7_port, IR_OUT4s_6_port, IR_OUT4s_5_port, IR_OUT4s_4_port, 
      IR_OUT4s_3_port, IR_OUT4s_2_port, IR_OUT4s_1_port, IR_OUT4s_0_port, 
      IR_OUT2s_31_port, IR_OUT2s_30_port, IR_OUT2s_29_port, IR_OUT2s_28_port, 
      IR_OUT2s_27_port, IR_OUT2s_26_port, IR_OUT2s_25_port, IR_OUT2s_24_port, 
      IR_OUT2s_23_port, IR_OUT2s_22_port, IR_OUT2s_21_port, IR_OUT2s_20_port, 
      IR_OUT2s_19_port, IR_OUT2s_18_port, IR_OUT2s_17_port, IR_OUT2s_16_port, 
      IR_OUT2s_15_port, IR_OUT2s_14_port, IR_OUT2s_13_port, IR_OUT2s_12_port, 
      IR_OUT2s_11_port, IR_OUT2s_10_port, IR_OUT2s_9_port, IR_OUT2s_8_port, 
      IR_OUT2s_7_port, IR_OUT2s_6_port, IR_OUT2s_5_port, IR_OUT2s_4_port, 
      IR_OUT2s_3_port, IR_OUT2s_2_port, IR_OUT2s_1_port, IR_OUT2s_0_port, 
      NPC2_OUTs_31_port, NPC2_OUTs_30_port, NPC2_OUTs_29_port, 
      NPC2_OUTs_28_port, NPC2_OUTs_27_port, NPC2_OUTs_26_port, 
      NPC2_OUTs_25_port, NPC2_OUTs_24_port, NPC2_OUTs_23_port, 
      NPC2_OUTs_22_port, NPC2_OUTs_21_port, NPC2_OUTs_20_port, 
      NPC2_OUTs_19_port, NPC2_OUTs_18_port, NPC2_OUTs_17_port, 
      NPC2_OUTs_16_port, NPC2_OUTs_15_port, NPC2_OUTs_14_port, 
      NPC2_OUTs_13_port, NPC2_OUTs_12_port, NPC2_OUTs_11_port, 
      NPC2_OUTs_10_port, NPC2_OUTs_9_port, NPC2_OUTs_8_port, NPC2_OUTs_7_port, 
      NPC2_OUTs_6_port, NPC2_OUTs_5_port, NPC2_OUTs_4_port, NPC2_OUTs_3_port, 
      NPC2_OUTs_2_port, NPC2_OUTs_1_port, NPC2_OUTs_0_port, COND_OUTs, 
      IR_OUT3s_31_port, IR_OUT3s_30_port, IR_OUT3s_29_port, IR_OUT3s_28_port, 
      IR_OUT3s_27_port, IR_OUT3s_26_port, IR_OUT3s_25_port, IR_OUT3s_24_port, 
      IR_OUT3s_23_port, IR_OUT3s_22_port, IR_OUT3s_21_port, IR_OUT3s_20_port, 
      IR_OUT3s_19_port, IR_OUT3s_18_port, IR_OUT3s_17_port, IR_OUT3s_16_port, 
      IR_OUT3s_15_port, IR_OUT3s_14_port, IR_OUT3s_13_port, IR_OUT3s_12_port, 
      IR_OUT3s_11_port, IR_OUT3s_10_port, IR_OUT3s_9_port, IR_OUT3s_8_port, 
      IR_OUT3s_7_port, IR_OUT3s_6_port, IR_OUT3s_5_port, IR_OUT3s_4_port, 
      IR_OUT3s_3_port, IR_OUT3s_2_port, IR_OUT3s_1_port, IR_OUT3s_0_port, 
      LMD_OUTs_31_port, LMD_OUTs_30_port, LMD_OUTs_29_port, LMD_OUTs_28_port, 
      LMD_OUTs_27_port, LMD_OUTs_26_port, LMD_OUTs_25_port, LMD_OUTs_24_port, 
      LMD_OUTs_23_port, LMD_OUTs_22_port, LMD_OUTs_21_port, LMD_OUTs_20_port, 
      LMD_OUTs_19_port, LMD_OUTs_18_port, LMD_OUTs_17_port, LMD_OUTs_16_port, 
      LMD_OUTs_15_port, LMD_OUTs_14_port, LMD_OUTs_13_port, LMD_OUTs_12_port, 
      LMD_OUTs_11_port, LMD_OUTs_10_port, LMD_OUTs_9_port, LMD_OUTs_8_port, 
      LMD_OUTs_7_port, LMD_OUTs_6_port, LMD_OUTs_5_port, LMD_OUTs_4_port, 
      LMD_OUTs_3_port, LMD_OUTs_2_port, LMD_OUTs_1_port, LMD_OUTs_0_port, 
      ALU_OUT2s_31_port, ALU_OUT2s_30_port, ALU_OUT2s_29_port, 
      ALU_OUT2s_28_port, ALU_OUT2s_27_port, ALU_OUT2s_26_port, 
      ALU_OUT2s_25_port, ALU_OUT2s_24_port, ALU_OUT2s_23_port, 
      ALU_OUT2s_22_port, ALU_OUT2s_21_port, ALU_OUT2s_20_port, 
      ALU_OUT2s_19_port, ALU_OUT2s_18_port, ALU_OUT2s_17_port, 
      ALU_OUT2s_16_port, ALU_OUT2s_15_port, ALU_OUT2s_14_port, 
      ALU_OUT2s_13_port, ALU_OUT2s_12_port, ALU_OUT2s_11_port, 
      ALU_OUT2s_10_port, ALU_OUT2s_9_port, ALU_OUT2s_8_port, ALU_OUT2s_7_port, 
      ALU_OUT2s_6_port, ALU_OUT2s_5_port, ALU_OUT2s_4_port, ALU_OUT2s_3_port, 
      ALU_OUT2s_2_port, ALU_OUT2s_1_port, ALU_OUT2s_0_port, n3, n4 : std_logic;

begin
   ALU_OUT <= ( ALU_OUT_31_port, ALU_OUT_30_port, ALU_OUT_29_port, 
      ALU_OUT_28_port, ALU_OUT_27_port, ALU_OUT_26_port, ALU_OUT_25_port, 
      ALU_OUT_24_port, ALU_OUT_23_port, ALU_OUT_22_port, ALU_OUT_21_port, 
      ALU_OUT_20_port, ALU_OUT_19_port, ALU_OUT_18_port, ALU_OUT_17_port, 
      ALU_OUT_16_port, ALU_OUT_15_port, ALU_OUT_14_port, ALU_OUT_13_port, 
      ALU_OUT_12_port, ALU_OUT_11_port, ALU_OUT_10_port, ALU_OUT_9_port, 
      ALU_OUT_8_port, ALU_OUT_7_port, ALU_OUT_6_port, ALU_OUT_5_port, 
      ALU_OUT_4_port, ALU_OUT_3_port, ALU_OUT_2_port, ALU_OUT_1_port, 
      ALU_OUT_0_port );
   IR_OUT <= ( IR_OUT_31_port, IR_OUT_30_port, IR_OUT_29_port, IR_OUT_28_port, 
      IR_OUT_27_port, IR_OUT_26_port, IR_OUT_25_port, IR_OUT_24_port, 
      IR_OUT_23_port, IR_OUT_22_port, IR_OUT_21_port, IR_OUT_20_port, 
      IR_OUT_19_port, IR_OUT_18_port, IR_OUT_17_port, IR_OUT_16_port, 
      IR_OUT_15_port, IR_OUT_14_port, IR_OUT_13_port, IR_OUT_12_port, 
      IR_OUT_11_port, IR_OUT_10_port, IR_OUT_9_port, IR_OUT_8_port, 
      IR_OUT_7_port, IR_OUT_6_port, IR_OUT_5_port, IR_OUT_4_port, IR_OUT_3_port
      , IR_OUT_2_port, IR_OUT_1_port, IR_OUT_0_port );
   
   FETCH : fetchUnit_nbits32 port map( clk => n4, rst => n3, DATA_IRAM(31) => 
                           DATA_IRAM(31), DATA_IRAM(30) => DATA_IRAM(30), 
                           DATA_IRAM(29) => DATA_IRAM(29), DATA_IRAM(28) => 
                           DATA_IRAM(28), DATA_IRAM(27) => DATA_IRAM(27), 
                           DATA_IRAM(26) => DATA_IRAM(26), DATA_IRAM(25) => 
                           DATA_IRAM(25), DATA_IRAM(24) => DATA_IRAM(24), 
                           DATA_IRAM(23) => DATA_IRAM(23), DATA_IRAM(22) => 
                           DATA_IRAM(22), DATA_IRAM(21) => DATA_IRAM(21), 
                           DATA_IRAM(20) => DATA_IRAM(20), DATA_IRAM(19) => 
                           DATA_IRAM(19), DATA_IRAM(18) => DATA_IRAM(18), 
                           DATA_IRAM(17) => DATA_IRAM(17), DATA_IRAM(16) => 
                           DATA_IRAM(16), DATA_IRAM(15) => DATA_IRAM(15), 
                           DATA_IRAM(14) => DATA_IRAM(14), DATA_IRAM(13) => 
                           DATA_IRAM(13), DATA_IRAM(12) => DATA_IRAM(12), 
                           DATA_IRAM(11) => DATA_IRAM(11), DATA_IRAM(10) => 
                           DATA_IRAM(10), DATA_IRAM(9) => DATA_IRAM(9), 
                           DATA_IRAM(8) => DATA_IRAM(8), DATA_IRAM(7) => 
                           DATA_IRAM(7), DATA_IRAM(6) => DATA_IRAM(6), 
                           DATA_IRAM(5) => DATA_IRAM(5), DATA_IRAM(4) => 
                           DATA_IRAM(4), DATA_IRAM(3) => DATA_IRAM(3), 
                           DATA_IRAM(2) => DATA_IRAM(2), DATA_IRAM(1) => 
                           DATA_IRAM(1), DATA_IRAM(0) => DATA_IRAM(0), 
                           IR_LATCH_EN => IR_LATCH_EN, NPC_LATCH_EN => 
                           NPC_LATCH_EN, PC_LATCH_EN => PC_LATCH_EN, PC_IN(31) 
                           => TO_PC_OUTs_31_port, PC_IN(30) => 
                           TO_PC_OUTs_30_port, PC_IN(29) => TO_PC_OUTs_29_port,
                           PC_IN(28) => TO_PC_OUTs_28_port, PC_IN(27) => 
                           TO_PC_OUTs_27_port, PC_IN(26) => TO_PC_OUTs_26_port,
                           PC_IN(25) => TO_PC_OUTs_25_port, PC_IN(24) => 
                           TO_PC_OUTs_24_port, PC_IN(23) => TO_PC_OUTs_23_port,
                           PC_IN(22) => TO_PC_OUTs_22_port, PC_IN(21) => 
                           TO_PC_OUTs_21_port, PC_IN(20) => TO_PC_OUTs_20_port,
                           PC_IN(19) => TO_PC_OUTs_19_port, PC_IN(18) => 
                           TO_PC_OUTs_18_port, PC_IN(17) => TO_PC_OUTs_17_port,
                           PC_IN(16) => TO_PC_OUTs_16_port, PC_IN(15) => 
                           TO_PC_OUTs_15_port, PC_IN(14) => TO_PC_OUTs_14_port,
                           PC_IN(13) => TO_PC_OUTs_13_port, PC_IN(12) => 
                           TO_PC_OUTs_12_port, PC_IN(11) => TO_PC_OUTs_11_port,
                           PC_IN(10) => TO_PC_OUTs_10_port, PC_IN(9) => 
                           TO_PC_OUTs_9_port, PC_IN(8) => TO_PC_OUTs_8_port, 
                           PC_IN(7) => TO_PC_OUTs_7_port, PC_IN(6) => 
                           TO_PC_OUTs_6_port, PC_IN(5) => TO_PC_OUTs_5_port, 
                           PC_IN(4) => TO_PC_OUTs_4_port, PC_IN(3) => 
                           TO_PC_OUTs_3_port, PC_IN(2) => TO_PC_OUTs_2_port, 
                           PC_IN(1) => TO_PC_OUTs_1_port, PC_IN(0) => 
                           TO_PC_OUTs_0_port, ADDRESS_IRAM(31) => 
                           ADDRESS_IRAM(31), ADDRESS_IRAM(30) => 
                           ADDRESS_IRAM(30), ADDRESS_IRAM(29) => 
                           ADDRESS_IRAM(29), ADDRESS_IRAM(28) => 
                           ADDRESS_IRAM(28), ADDRESS_IRAM(27) => 
                           ADDRESS_IRAM(27), ADDRESS_IRAM(26) => 
                           ADDRESS_IRAM(26), ADDRESS_IRAM(25) => 
                           ADDRESS_IRAM(25), ADDRESS_IRAM(24) => 
                           ADDRESS_IRAM(24), ADDRESS_IRAM(23) => 
                           ADDRESS_IRAM(23), ADDRESS_IRAM(22) => 
                           ADDRESS_IRAM(22), ADDRESS_IRAM(21) => 
                           ADDRESS_IRAM(21), ADDRESS_IRAM(20) => 
                           ADDRESS_IRAM(20), ADDRESS_IRAM(19) => 
                           ADDRESS_IRAM(19), ADDRESS_IRAM(18) => 
                           ADDRESS_IRAM(18), ADDRESS_IRAM(17) => 
                           ADDRESS_IRAM(17), ADDRESS_IRAM(16) => 
                           ADDRESS_IRAM(16), ADDRESS_IRAM(15) => 
                           ADDRESS_IRAM(15), ADDRESS_IRAM(14) => 
                           ADDRESS_IRAM(14), ADDRESS_IRAM(13) => 
                           ADDRESS_IRAM(13), ADDRESS_IRAM(12) => 
                           ADDRESS_IRAM(12), ADDRESS_IRAM(11) => 
                           ADDRESS_IRAM(11), ADDRESS_IRAM(10) => 
                           ADDRESS_IRAM(10), ADDRESS_IRAM(9) => ADDRESS_IRAM(9)
                           , ADDRESS_IRAM(8) => ADDRESS_IRAM(8), 
                           ADDRESS_IRAM(7) => ADDRESS_IRAM(7), ADDRESS_IRAM(6) 
                           => ADDRESS_IRAM(6), ADDRESS_IRAM(5) => 
                           ADDRESS_IRAM(5), ADDRESS_IRAM(4) => ADDRESS_IRAM(4),
                           ADDRESS_IRAM(3) => ADDRESS_IRAM(3), ADDRESS_IRAM(2) 
                           => ADDRESS_IRAM(2), ADDRESS_IRAM(1) => 
                           ADDRESS_IRAM(1), ADDRESS_IRAM(0) => ADDRESS_IRAM(0),
                           NPC_OUT(31) => NPC_OUTs_31_port, NPC_OUT(30) => 
                           NPC_OUTs_30_port, NPC_OUT(29) => NPC_OUTs_29_port, 
                           NPC_OUT(28) => NPC_OUTs_28_port, NPC_OUT(27) => 
                           NPC_OUTs_27_port, NPC_OUT(26) => NPC_OUTs_26_port, 
                           NPC_OUT(25) => NPC_OUTs_25_port, NPC_OUT(24) => 
                           NPC_OUTs_24_port, NPC_OUT(23) => NPC_OUTs_23_port, 
                           NPC_OUT(22) => NPC_OUTs_22_port, NPC_OUT(21) => 
                           NPC_OUTs_21_port, NPC_OUT(20) => NPC_OUTs_20_port, 
                           NPC_OUT(19) => NPC_OUTs_19_port, NPC_OUT(18) => 
                           NPC_OUTs_18_port, NPC_OUT(17) => NPC_OUTs_17_port, 
                           NPC_OUT(16) => NPC_OUTs_16_port, NPC_OUT(15) => 
                           NPC_OUTs_15_port, NPC_OUT(14) => NPC_OUTs_14_port, 
                           NPC_OUT(13) => NPC_OUTs_13_port, NPC_OUT(12) => 
                           NPC_OUTs_12_port, NPC_OUT(11) => NPC_OUTs_11_port, 
                           NPC_OUT(10) => NPC_OUTs_10_port, NPC_OUT(9) => 
                           NPC_OUTs_9_port, NPC_OUT(8) => NPC_OUTs_8_port, 
                           NPC_OUT(7) => NPC_OUTs_7_port, NPC_OUT(6) => 
                           NPC_OUTs_6_port, NPC_OUT(5) => NPC_OUTs_5_port, 
                           NPC_OUT(4) => NPC_OUTs_4_port, NPC_OUT(3) => 
                           NPC_OUTs_3_port, NPC_OUT(2) => NPC_OUTs_2_port, 
                           NPC_OUT(1) => NPC_OUTs_1_port, NPC_OUT(0) => 
                           NPC_OUTs_0_port, IR_OUT(31) => IR_OUT_31_port, 
                           IR_OUT(30) => IR_OUT_30_port, IR_OUT(29) => 
                           IR_OUT_29_port, IR_OUT(28) => IR_OUT_28_port, 
                           IR_OUT(27) => IR_OUT_27_port, IR_OUT(26) => 
                           IR_OUT_26_port, IR_OUT(25) => IR_OUT_25_port, 
                           IR_OUT(24) => IR_OUT_24_port, IR_OUT(23) => 
                           IR_OUT_23_port, IR_OUT(22) => IR_OUT_22_port, 
                           IR_OUT(21) => IR_OUT_21_port, IR_OUT(20) => 
                           IR_OUT_20_port, IR_OUT(19) => IR_OUT_19_port, 
                           IR_OUT(18) => IR_OUT_18_port, IR_OUT(17) => 
                           IR_OUT_17_port, IR_OUT(16) => IR_OUT_16_port, 
                           IR_OUT(15) => IR_OUT_15_port, IR_OUT(14) => 
                           IR_OUT_14_port, IR_OUT(13) => IR_OUT_13_port, 
                           IR_OUT(12) => IR_OUT_12_port, IR_OUT(11) => 
                           IR_OUT_11_port, IR_OUT(10) => IR_OUT_10_port, 
                           IR_OUT(9) => IR_OUT_9_port, IR_OUT(8) => 
                           IR_OUT_8_port, IR_OUT(7) => IR_OUT_7_port, IR_OUT(6)
                           => IR_OUT_6_port, IR_OUT(5) => IR_OUT_5_port, 
                           IR_OUT(4) => IR_OUT_4_port, IR_OUT(3) => 
                           IR_OUT_3_port, IR_OUT(2) => IR_OUT_2_port, IR_OUT(1)
                           => IR_OUT_1_port, IR_OUT(0) => IR_OUT_0_port, 
                           ADDERPC_OUT(31) => ADDERPC_OUTs_31_port, 
                           ADDERPC_OUT(30) => ADDERPC_OUTs_30_port, 
                           ADDERPC_OUT(29) => ADDERPC_OUTs_29_port, 
                           ADDERPC_OUT(28) => ADDERPC_OUTs_28_port, 
                           ADDERPC_OUT(27) => ADDERPC_OUTs_27_port, 
                           ADDERPC_OUT(26) => ADDERPC_OUTs_26_port, 
                           ADDERPC_OUT(25) => ADDERPC_OUTs_25_port, 
                           ADDERPC_OUT(24) => ADDERPC_OUTs_24_port, 
                           ADDERPC_OUT(23) => ADDERPC_OUTs_23_port, 
                           ADDERPC_OUT(22) => ADDERPC_OUTs_22_port, 
                           ADDERPC_OUT(21) => ADDERPC_OUTs_21_port, 
                           ADDERPC_OUT(20) => ADDERPC_OUTs_20_port, 
                           ADDERPC_OUT(19) => ADDERPC_OUTs_19_port, 
                           ADDERPC_OUT(18) => ADDERPC_OUTs_18_port, 
                           ADDERPC_OUT(17) => ADDERPC_OUTs_17_port, 
                           ADDERPC_OUT(16) => ADDERPC_OUTs_16_port, 
                           ADDERPC_OUT(15) => ADDERPC_OUTs_15_port, 
                           ADDERPC_OUT(14) => ADDERPC_OUTs_14_port, 
                           ADDERPC_OUT(13) => ADDERPC_OUTs_13_port, 
                           ADDERPC_OUT(12) => ADDERPC_OUTs_12_port, 
                           ADDERPC_OUT(11) => ADDERPC_OUTs_11_port, 
                           ADDERPC_OUT(10) => ADDERPC_OUTs_10_port, 
                           ADDERPC_OUT(9) => ADDERPC_OUTs_9_port, 
                           ADDERPC_OUT(8) => ADDERPC_OUTs_8_port, 
                           ADDERPC_OUT(7) => ADDERPC_OUTs_7_port, 
                           ADDERPC_OUT(6) => ADDERPC_OUTs_6_port, 
                           ADDERPC_OUT(5) => ADDERPC_OUTs_5_port, 
                           ADDERPC_OUT(4) => ADDERPC_OUTs_4_port, 
                           ADDERPC_OUT(3) => ADDERPC_OUTs_3_port, 
                           ADDERPC_OUT(2) => ADDERPC_OUTs_2_port, 
                           ADDERPC_OUT(1) => ADDERPC_OUTs_1_port, 
                           ADDERPC_OUT(0) => ADDERPC_OUTs_0_port);
   DECODE : decodeUnit_nbits32 port map( clk => n4, rst => n3, RegA_LATCH_EN =>
                           RegA_LATCH_EN, RegB_LATCH_EN => RegB_LATCH_EN, 
                           RegIMM_LATCH_EN => RegIMM_LATCH_EN, RF_WE => RF_WE, 
                           DATAIN(31) => DATAIN_RFs_31_port, DATAIN(30) => 
                           DATAIN_RFs_30_port, DATAIN(29) => DATAIN_RFs_29_port
                           , DATAIN(28) => DATAIN_RFs_28_port, DATAIN(27) => 
                           DATAIN_RFs_27_port, DATAIN(26) => DATAIN_RFs_26_port
                           , DATAIN(25) => DATAIN_RFs_25_port, DATAIN(24) => 
                           DATAIN_RFs_24_port, DATAIN(23) => DATAIN_RFs_23_port
                           , DATAIN(22) => DATAIN_RFs_22_port, DATAIN(21) => 
                           DATAIN_RFs_21_port, DATAIN(20) => DATAIN_RFs_20_port
                           , DATAIN(19) => DATAIN_RFs_19_port, DATAIN(18) => 
                           DATAIN_RFs_18_port, DATAIN(17) => DATAIN_RFs_17_port
                           , DATAIN(16) => DATAIN_RFs_16_port, DATAIN(15) => 
                           DATAIN_RFs_15_port, DATAIN(14) => DATAIN_RFs_14_port
                           , DATAIN(13) => DATAIN_RFs_13_port, DATAIN(12) => 
                           DATAIN_RFs_12_port, DATAIN(11) => DATAIN_RFs_11_port
                           , DATAIN(10) => DATAIN_RFs_10_port, DATAIN(9) => 
                           DATAIN_RFs_9_port, DATAIN(8) => DATAIN_RFs_8_port, 
                           DATAIN(7) => DATAIN_RFs_7_port, DATAIN(6) => 
                           DATAIN_RFs_6_port, DATAIN(5) => DATAIN_RFs_5_port, 
                           DATAIN(4) => DATAIN_RFs_4_port, DATAIN(3) => 
                           DATAIN_RFs_3_port, DATAIN(2) => DATAIN_RFs_2_port, 
                           DATAIN(1) => DATAIN_RFs_1_port, DATAIN(0) => 
                           DATAIN_RFs_0_port, IR_OUT(31) => IR_OUT_31_port, 
                           IR_OUT(30) => IR_OUT_30_port, IR_OUT(29) => 
                           IR_OUT_29_port, IR_OUT(28) => IR_OUT_28_port, 
                           IR_OUT(27) => IR_OUT_27_port, IR_OUT(26) => 
                           IR_OUT_26_port, IR_OUT(25) => IR_OUT_25_port, 
                           IR_OUT(24) => IR_OUT_24_port, IR_OUT(23) => 
                           IR_OUT_23_port, IR_OUT(22) => IR_OUT_22_port, 
                           IR_OUT(21) => IR_OUT_21_port, IR_OUT(20) => 
                           IR_OUT_20_port, IR_OUT(19) => IR_OUT_19_port, 
                           IR_OUT(18) => IR_OUT_18_port, IR_OUT(17) => 
                           IR_OUT_17_port, IR_OUT(16) => IR_OUT_16_port, 
                           IR_OUT(15) => IR_OUT_15_port, IR_OUT(14) => 
                           IR_OUT_14_port, IR_OUT(13) => IR_OUT_13_port, 
                           IR_OUT(12) => IR_OUT_12_port, IR_OUT(11) => 
                           IR_OUT_11_port, IR_OUT(10) => IR_OUT_10_port, 
                           IR_OUT(9) => IR_OUT_9_port, IR_OUT(8) => 
                           IR_OUT_8_port, IR_OUT(7) => IR_OUT_7_port, IR_OUT(6)
                           => IR_OUT_6_port, IR_OUT(5) => IR_OUT_5_port, 
                           IR_OUT(4) => IR_OUT_4_port, IR_OUT(3) => 
                           IR_OUT_3_port, IR_OUT(2) => IR_OUT_2_port, IR_OUT(1)
                           => IR_OUT_1_port, IR_OUT(0) => IR_OUT_0_port, 
                           A_out(31) => A_outs_31_port, A_out(30) => 
                           A_outs_30_port, A_out(29) => A_outs_29_port, 
                           A_out(28) => A_outs_28_port, A_out(27) => 
                           A_outs_27_port, A_out(26) => A_outs_26_port, 
                           A_out(25) => A_outs_25_port, A_out(24) => 
                           A_outs_24_port, A_out(23) => A_outs_23_port, 
                           A_out(22) => A_outs_22_port, A_out(21) => 
                           A_outs_21_port, A_out(20) => A_outs_20_port, 
                           A_out(19) => A_outs_19_port, A_out(18) => 
                           A_outs_18_port, A_out(17) => A_outs_17_port, 
                           A_out(16) => A_outs_16_port, A_out(15) => 
                           A_outs_15_port, A_out(14) => A_outs_14_port, 
                           A_out(13) => A_outs_13_port, A_out(12) => 
                           A_outs_12_port, A_out(11) => A_outs_11_port, 
                           A_out(10) => A_outs_10_port, A_out(9) => 
                           A_outs_9_port, A_out(8) => A_outs_8_port, A_out(7) 
                           => A_outs_7_port, A_out(6) => A_outs_6_port, 
                           A_out(5) => A_outs_5_port, A_out(4) => A_outs_4_port
                           , A_out(3) => A_outs_3_port, A_out(2) => 
                           A_outs_2_port, A_out(1) => A_outs_1_port, A_out(0) 
                           => A_outs_0_port, B_out(31) => B_outs_31_port, 
                           B_out(30) => B_outs_30_port, B_out(29) => 
                           B_outs_29_port, B_out(28) => B_outs_28_port, 
                           B_out(27) => B_outs_27_port, B_out(26) => 
                           B_outs_26_port, B_out(25) => B_outs_25_port, 
                           B_out(24) => B_outs_24_port, B_out(23) => 
                           B_outs_23_port, B_out(22) => B_outs_22_port, 
                           B_out(21) => B_outs_21_port, B_out(20) => 
                           B_outs_20_port, B_out(19) => B_outs_19_port, 
                           B_out(18) => B_outs_18_port, B_out(17) => 
                           B_outs_17_port, B_out(16) => B_outs_16_port, 
                           B_out(15) => B_outs_15_port, B_out(14) => 
                           B_outs_14_port, B_out(13) => B_outs_13_port, 
                           B_out(12) => B_outs_12_port, B_out(11) => 
                           B_outs_11_port, B_out(10) => B_outs_10_port, 
                           B_out(9) => B_outs_9_port, B_out(8) => B_outs_8_port
                           , B_out(7) => B_outs_7_port, B_out(6) => 
                           B_outs_6_port, B_out(5) => B_outs_5_port, B_out(4) 
                           => B_outs_4_port, B_out(3) => B_outs_3_port, 
                           B_out(2) => B_outs_2_port, B_out(1) => B_outs_1_port
                           , B_out(0) => B_outs_0_port, Imm_out(31) => 
                           Imm_outs_31_port, Imm_out(30) => Imm_outs_30_port, 
                           Imm_out(29) => Imm_outs_29_port, Imm_out(28) => 
                           Imm_outs_28_port, Imm_out(27) => Imm_outs_27_port, 
                           Imm_out(26) => Imm_outs_26_port, Imm_out(25) => 
                           Imm_outs_25_port, Imm_out(24) => Imm_outs_24_port, 
                           Imm_out(23) => Imm_outs_23_port, Imm_out(22) => 
                           Imm_outs_22_port, Imm_out(21) => Imm_outs_21_port, 
                           Imm_out(20) => Imm_outs_20_port, Imm_out(19) => 
                           Imm_outs_19_port, Imm_out(18) => Imm_outs_18_port, 
                           Imm_out(17) => Imm_outs_17_port, Imm_out(16) => 
                           Imm_outs_16_port, Imm_out(15) => Imm_outs_15_port, 
                           Imm_out(14) => Imm_outs_14_port, Imm_out(13) => 
                           Imm_outs_13_port, Imm_out(12) => Imm_outs_12_port, 
                           Imm_out(11) => Imm_outs_11_port, Imm_out(10) => 
                           Imm_outs_10_port, Imm_out(9) => Imm_outs_9_port, 
                           Imm_out(8) => Imm_outs_8_port, Imm_out(7) => 
                           Imm_outs_7_port, Imm_out(6) => Imm_outs_6_port, 
                           Imm_out(5) => Imm_outs_5_port, Imm_out(4) => 
                           Imm_outs_4_port, Imm_out(3) => Imm_outs_3_port, 
                           Imm_out(2) => Imm_outs_2_port, Imm_out(1) => 
                           Imm_outs_1_port, Imm_out(0) => Imm_outs_0_port, 
                           IR_IN2(31) => IR_OUT4s_31_port, IR_IN2(30) => 
                           IR_OUT4s_30_port, IR_IN2(29) => IR_OUT4s_29_port, 
                           IR_IN2(28) => IR_OUT4s_28_port, IR_IN2(27) => 
                           IR_OUT4s_27_port, IR_IN2(26) => IR_OUT4s_26_port, 
                           IR_IN2(25) => IR_OUT4s_25_port, IR_IN2(24) => 
                           IR_OUT4s_24_port, IR_IN2(23) => IR_OUT4s_23_port, 
                           IR_IN2(22) => IR_OUT4s_22_port, IR_IN2(21) => 
                           IR_OUT4s_21_port, IR_IN2(20) => IR_OUT4s_20_port, 
                           IR_IN2(19) => IR_OUT4s_19_port, IR_IN2(18) => 
                           IR_OUT4s_18_port, IR_IN2(17) => IR_OUT4s_17_port, 
                           IR_IN2(16) => IR_OUT4s_16_port, IR_IN2(15) => 
                           IR_OUT4s_15_port, IR_IN2(14) => IR_OUT4s_14_port, 
                           IR_IN2(13) => IR_OUT4s_13_port, IR_IN2(12) => 
                           IR_OUT4s_12_port, IR_IN2(11) => IR_OUT4s_11_port, 
                           IR_IN2(10) => IR_OUT4s_10_port, IR_IN2(9) => 
                           IR_OUT4s_9_port, IR_IN2(8) => IR_OUT4s_8_port, 
                           IR_IN2(7) => IR_OUT4s_7_port, IR_IN2(6) => 
                           IR_OUT4s_6_port, IR_IN2(5) => IR_OUT4s_5_port, 
                           IR_IN2(4) => IR_OUT4s_4_port, IR_IN2(3) => 
                           IR_OUT4s_3_port, IR_IN2(2) => IR_OUT4s_2_port, 
                           IR_IN2(1) => IR_OUT4s_1_port, IR_IN2(0) => 
                           IR_OUT4s_0_port, IR_OUT2(31) => IR_OUT2s_31_port, 
                           IR_OUT2(30) => IR_OUT2s_30_port, IR_OUT2(29) => 
                           IR_OUT2s_29_port, IR_OUT2(28) => IR_OUT2s_28_port, 
                           IR_OUT2(27) => IR_OUT2s_27_port, IR_OUT2(26) => 
                           IR_OUT2s_26_port, IR_OUT2(25) => IR_OUT2s_25_port, 
                           IR_OUT2(24) => IR_OUT2s_24_port, IR_OUT2(23) => 
                           IR_OUT2s_23_port, IR_OUT2(22) => IR_OUT2s_22_port, 
                           IR_OUT2(21) => IR_OUT2s_21_port, IR_OUT2(20) => 
                           IR_OUT2s_20_port, IR_OUT2(19) => IR_OUT2s_19_port, 
                           IR_OUT2(18) => IR_OUT2s_18_port, IR_OUT2(17) => 
                           IR_OUT2s_17_port, IR_OUT2(16) => IR_OUT2s_16_port, 
                           IR_OUT2(15) => IR_OUT2s_15_port, IR_OUT2(14) => 
                           IR_OUT2s_14_port, IR_OUT2(13) => IR_OUT2s_13_port, 
                           IR_OUT2(12) => IR_OUT2s_12_port, IR_OUT2(11) => 
                           IR_OUT2s_11_port, IR_OUT2(10) => IR_OUT2s_10_port, 
                           IR_OUT2(9) => IR_OUT2s_9_port, IR_OUT2(8) => 
                           IR_OUT2s_8_port, IR_OUT2(7) => IR_OUT2s_7_port, 
                           IR_OUT2(6) => IR_OUT2s_6_port, IR_OUT2(5) => 
                           IR_OUT2s_5_port, IR_OUT2(4) => IR_OUT2s_4_port, 
                           IR_OUT2(3) => IR_OUT2s_3_port, IR_OUT2(2) => 
                           IR_OUT2s_2_port, IR_OUT2(1) => IR_OUT2s_1_port, 
                           IR_OUT2(0) => IR_OUT2s_0_port, NPC_IN(31) => 
                           NPC_OUTs_31_port, NPC_IN(30) => NPC_OUTs_30_port, 
                           NPC_IN(29) => NPC_OUTs_29_port, NPC_IN(28) => 
                           NPC_OUTs_28_port, NPC_IN(27) => NPC_OUTs_27_port, 
                           NPC_IN(26) => NPC_OUTs_26_port, NPC_IN(25) => 
                           NPC_OUTs_25_port, NPC_IN(24) => NPC_OUTs_24_port, 
                           NPC_IN(23) => NPC_OUTs_23_port, NPC_IN(22) => 
                           NPC_OUTs_22_port, NPC_IN(21) => NPC_OUTs_21_port, 
                           NPC_IN(20) => NPC_OUTs_20_port, NPC_IN(19) => 
                           NPC_OUTs_19_port, NPC_IN(18) => NPC_OUTs_18_port, 
                           NPC_IN(17) => NPC_OUTs_17_port, NPC_IN(16) => 
                           NPC_OUTs_16_port, NPC_IN(15) => NPC_OUTs_15_port, 
                           NPC_IN(14) => NPC_OUTs_14_port, NPC_IN(13) => 
                           NPC_OUTs_13_port, NPC_IN(12) => NPC_OUTs_12_port, 
                           NPC_IN(11) => NPC_OUTs_11_port, NPC_IN(10) => 
                           NPC_OUTs_10_port, NPC_IN(9) => NPC_OUTs_9_port, 
                           NPC_IN(8) => NPC_OUTs_8_port, NPC_IN(7) => 
                           NPC_OUTs_7_port, NPC_IN(6) => NPC_OUTs_6_port, 
                           NPC_IN(5) => NPC_OUTs_5_port, NPC_IN(4) => 
                           NPC_OUTs_4_port, NPC_IN(3) => NPC_OUTs_3_port, 
                           NPC_IN(2) => NPC_OUTs_2_port, NPC_IN(1) => 
                           NPC_OUTs_1_port, NPC_IN(0) => NPC_OUTs_0_port, 
                           NPC2_OUT(31) => NPC2_OUTs_31_port, NPC2_OUT(30) => 
                           NPC2_OUTs_30_port, NPC2_OUT(29) => NPC2_OUTs_29_port
                           , NPC2_OUT(28) => NPC2_OUTs_28_port, NPC2_OUT(27) =>
                           NPC2_OUTs_27_port, NPC2_OUT(26) => NPC2_OUTs_26_port
                           , NPC2_OUT(25) => NPC2_OUTs_25_port, NPC2_OUT(24) =>
                           NPC2_OUTs_24_port, NPC2_OUT(23) => NPC2_OUTs_23_port
                           , NPC2_OUT(22) => NPC2_OUTs_22_port, NPC2_OUT(21) =>
                           NPC2_OUTs_21_port, NPC2_OUT(20) => NPC2_OUTs_20_port
                           , NPC2_OUT(19) => NPC2_OUTs_19_port, NPC2_OUT(18) =>
                           NPC2_OUTs_18_port, NPC2_OUT(17) => NPC2_OUTs_17_port
                           , NPC2_OUT(16) => NPC2_OUTs_16_port, NPC2_OUT(15) =>
                           NPC2_OUTs_15_port, NPC2_OUT(14) => NPC2_OUTs_14_port
                           , NPC2_OUT(13) => NPC2_OUTs_13_port, NPC2_OUT(12) =>
                           NPC2_OUTs_12_port, NPC2_OUT(11) => NPC2_OUTs_11_port
                           , NPC2_OUT(10) => NPC2_OUTs_10_port, NPC2_OUT(9) => 
                           NPC2_OUTs_9_port, NPC2_OUT(8) => NPC2_OUTs_8_port, 
                           NPC2_OUT(7) => NPC2_OUTs_7_port, NPC2_OUT(6) => 
                           NPC2_OUTs_6_port, NPC2_OUT(5) => NPC2_OUTs_5_port, 
                           NPC2_OUT(4) => NPC2_OUTs_4_port, NPC2_OUT(3) => 
                           NPC2_OUTs_3_port, NPC2_OUT(2) => NPC2_OUTs_2_port, 
                           NPC2_OUT(1) => NPC2_OUTs_1_port, NPC2_OUT(0) => 
                           NPC2_OUTs_0_port);
   EXECUTE : executionUnit_nbits32 port map( clk => n4, rst => n3, 
                           ALU_OUTREG_ENABLE => ALU_OUTREG_EN, MUXA_SEL => 
                           MUXA_SEL, MUXB_SEL => MUXB_SEL, COND_ENABLE => 
                           EQ_COND, ALU_BITS(0) => ALU_OPCODE(0), ALU_BITS(1) 
                           => ALU_OPCODE(1), ALU_BITS(2) => ALU_OPCODE(2), 
                           ALU_BITS(3) => ALU_OPCODE(3), NPC_OUT(31) => 
                           NPC2_OUTs_31_port, NPC_OUT(30) => NPC2_OUTs_30_port,
                           NPC_OUT(29) => NPC2_OUTs_29_port, NPC_OUT(28) => 
                           NPC2_OUTs_28_port, NPC_OUT(27) => NPC2_OUTs_27_port,
                           NPC_OUT(26) => NPC2_OUTs_26_port, NPC_OUT(25) => 
                           NPC2_OUTs_25_port, NPC_OUT(24) => NPC2_OUTs_24_port,
                           NPC_OUT(23) => NPC2_OUTs_23_port, NPC_OUT(22) => 
                           NPC2_OUTs_22_port, NPC_OUT(21) => NPC2_OUTs_21_port,
                           NPC_OUT(20) => NPC2_OUTs_20_port, NPC_OUT(19) => 
                           NPC2_OUTs_19_port, NPC_OUT(18) => NPC2_OUTs_18_port,
                           NPC_OUT(17) => NPC2_OUTs_17_port, NPC_OUT(16) => 
                           NPC2_OUTs_16_port, NPC_OUT(15) => NPC2_OUTs_15_port,
                           NPC_OUT(14) => NPC2_OUTs_14_port, NPC_OUT(13) => 
                           NPC2_OUTs_13_port, NPC_OUT(12) => NPC2_OUTs_12_port,
                           NPC_OUT(11) => NPC2_OUTs_11_port, NPC_OUT(10) => 
                           NPC2_OUTs_10_port, NPC_OUT(9) => NPC2_OUTs_9_port, 
                           NPC_OUT(8) => NPC2_OUTs_8_port, NPC_OUT(7) => 
                           NPC2_OUTs_7_port, NPC_OUT(6) => NPC2_OUTs_6_port, 
                           NPC_OUT(5) => NPC2_OUTs_5_port, NPC_OUT(4) => 
                           NPC2_OUTs_4_port, NPC_OUT(3) => NPC2_OUTs_3_port, 
                           NPC_OUT(2) => NPC2_OUTs_2_port, NPC_OUT(1) => 
                           NPC2_OUTs_1_port, NPC_OUT(0) => NPC2_OUTs_0_port, 
                           A_out(31) => A_outs_31_port, A_out(30) => 
                           A_outs_30_port, A_out(29) => A_outs_29_port, 
                           A_out(28) => A_outs_28_port, A_out(27) => 
                           A_outs_27_port, A_out(26) => A_outs_26_port, 
                           A_out(25) => A_outs_25_port, A_out(24) => 
                           A_outs_24_port, A_out(23) => A_outs_23_port, 
                           A_out(22) => A_outs_22_port, A_out(21) => 
                           A_outs_21_port, A_out(20) => A_outs_20_port, 
                           A_out(19) => A_outs_19_port, A_out(18) => 
                           A_outs_18_port, A_out(17) => A_outs_17_port, 
                           A_out(16) => A_outs_16_port, A_out(15) => 
                           A_outs_15_port, A_out(14) => A_outs_14_port, 
                           A_out(13) => A_outs_13_port, A_out(12) => 
                           A_outs_12_port, A_out(11) => A_outs_11_port, 
                           A_out(10) => A_outs_10_port, A_out(9) => 
                           A_outs_9_port, A_out(8) => A_outs_8_port, A_out(7) 
                           => A_outs_7_port, A_out(6) => A_outs_6_port, 
                           A_out(5) => A_outs_5_port, A_out(4) => A_outs_4_port
                           , A_out(3) => A_outs_3_port, A_out(2) => 
                           A_outs_2_port, A_out(1) => A_outs_1_port, A_out(0) 
                           => A_outs_0_port, B_out(31) => B_outs_31_port, 
                           B_out(30) => B_outs_30_port, B_out(29) => 
                           B_outs_29_port, B_out(28) => B_outs_28_port, 
                           B_out(27) => B_outs_27_port, B_out(26) => 
                           B_outs_26_port, B_out(25) => B_outs_25_port, 
                           B_out(24) => B_outs_24_port, B_out(23) => 
                           B_outs_23_port, B_out(22) => B_outs_22_port, 
                           B_out(21) => B_outs_21_port, B_out(20) => 
                           B_outs_20_port, B_out(19) => B_outs_19_port, 
                           B_out(18) => B_outs_18_port, B_out(17) => 
                           B_outs_17_port, B_out(16) => B_outs_16_port, 
                           B_out(15) => B_outs_15_port, B_out(14) => 
                           B_outs_14_port, B_out(13) => B_outs_13_port, 
                           B_out(12) => B_outs_12_port, B_out(11) => 
                           B_outs_11_port, B_out(10) => B_outs_10_port, 
                           B_out(9) => B_outs_9_port, B_out(8) => B_outs_8_port
                           , B_out(7) => B_outs_7_port, B_out(6) => 
                           B_outs_6_port, B_out(5) => B_outs_5_port, B_out(4) 
                           => B_outs_4_port, B_out(3) => B_outs_3_port, 
                           B_out(2) => B_outs_2_port, B_out(1) => B_outs_1_port
                           , B_out(0) => B_outs_0_port, Imm_out(31) => 
                           Imm_outs_31_port, Imm_out(30) => Imm_outs_30_port, 
                           Imm_out(29) => Imm_outs_29_port, Imm_out(28) => 
                           Imm_outs_28_port, Imm_out(27) => Imm_outs_27_port, 
                           Imm_out(26) => Imm_outs_26_port, Imm_out(25) => 
                           Imm_outs_25_port, Imm_out(24) => Imm_outs_24_port, 
                           Imm_out(23) => Imm_outs_23_port, Imm_out(22) => 
                           Imm_outs_22_port, Imm_out(21) => Imm_outs_21_port, 
                           Imm_out(20) => Imm_outs_20_port, Imm_out(19) => 
                           Imm_outs_19_port, Imm_out(18) => Imm_outs_18_port, 
                           Imm_out(17) => Imm_outs_17_port, Imm_out(16) => 
                           Imm_outs_16_port, Imm_out(15) => Imm_outs_15_port, 
                           Imm_out(14) => Imm_outs_14_port, Imm_out(13) => 
                           Imm_outs_13_port, Imm_out(12) => Imm_outs_12_port, 
                           Imm_out(11) => Imm_outs_11_port, Imm_out(10) => 
                           Imm_outs_10_port, Imm_out(9) => Imm_outs_9_port, 
                           Imm_out(8) => Imm_outs_8_port, Imm_out(7) => 
                           Imm_outs_7_port, Imm_out(6) => Imm_outs_6_port, 
                           Imm_out(5) => Imm_outs_5_port, Imm_out(4) => 
                           Imm_outs_4_port, Imm_out(3) => Imm_outs_3_port, 
                           Imm_out(2) => Imm_outs_2_port, Imm_out(1) => 
                           Imm_outs_1_port, Imm_out(0) => Imm_outs_0_port, 
                           ALUREG_OUTPUT(31) => ALU_OUT_31_port, 
                           ALUREG_OUTPUT(30) => ALU_OUT_30_port, 
                           ALUREG_OUTPUT(29) => ALU_OUT_29_port, 
                           ALUREG_OUTPUT(28) => ALU_OUT_28_port, 
                           ALUREG_OUTPUT(27) => ALU_OUT_27_port, 
                           ALUREG_OUTPUT(26) => ALU_OUT_26_port, 
                           ALUREG_OUTPUT(25) => ALU_OUT_25_port, 
                           ALUREG_OUTPUT(24) => ALU_OUT_24_port, 
                           ALUREG_OUTPUT(23) => ALU_OUT_23_port, 
                           ALUREG_OUTPUT(22) => ALU_OUT_22_port, 
                           ALUREG_OUTPUT(21) => ALU_OUT_21_port, 
                           ALUREG_OUTPUT(20) => ALU_OUT_20_port, 
                           ALUREG_OUTPUT(19) => ALU_OUT_19_port, 
                           ALUREG_OUTPUT(18) => ALU_OUT_18_port, 
                           ALUREG_OUTPUT(17) => ALU_OUT_17_port, 
                           ALUREG_OUTPUT(16) => ALU_OUT_16_port, 
                           ALUREG_OUTPUT(15) => ALU_OUT_15_port, 
                           ALUREG_OUTPUT(14) => ALU_OUT_14_port, 
                           ALUREG_OUTPUT(13) => ALU_OUT_13_port, 
                           ALUREG_OUTPUT(12) => ALU_OUT_12_port, 
                           ALUREG_OUTPUT(11) => ALU_OUT_11_port, 
                           ALUREG_OUTPUT(10) => ALU_OUT_10_port, 
                           ALUREG_OUTPUT(9) => ALU_OUT_9_port, ALUREG_OUTPUT(8)
                           => ALU_OUT_8_port, ALUREG_OUTPUT(7) => 
                           ALU_OUT_7_port, ALUREG_OUTPUT(6) => ALU_OUT_6_port, 
                           ALUREG_OUTPUT(5) => ALU_OUT_5_port, ALUREG_OUTPUT(4)
                           => ALU_OUT_4_port, ALUREG_OUTPUT(3) => 
                           ALU_OUT_3_port, ALUREG_OUTPUT(2) => ALU_OUT_2_port, 
                           ALUREG_OUTPUT(1) => ALU_OUT_1_port, ALUREG_OUTPUT(0)
                           => ALU_OUT_0_port, COND_OUT => COND_OUTs, IR_IN3(31)
                           => IR_OUT2s_31_port, IR_IN3(30) => IR_OUT2s_30_port,
                           IR_IN3(29) => IR_OUT2s_29_port, IR_IN3(28) => 
                           IR_OUT2s_28_port, IR_IN3(27) => IR_OUT2s_27_port, 
                           IR_IN3(26) => IR_OUT2s_26_port, IR_IN3(25) => 
                           IR_OUT2s_25_port, IR_IN3(24) => IR_OUT2s_24_port, 
                           IR_IN3(23) => IR_OUT2s_23_port, IR_IN3(22) => 
                           IR_OUT2s_22_port, IR_IN3(21) => IR_OUT2s_21_port, 
                           IR_IN3(20) => IR_OUT2s_20_port, IR_IN3(19) => 
                           IR_OUT2s_19_port, IR_IN3(18) => IR_OUT2s_18_port, 
                           IR_IN3(17) => IR_OUT2s_17_port, IR_IN3(16) => 
                           IR_OUT2s_16_port, IR_IN3(15) => IR_OUT2s_15_port, 
                           IR_IN3(14) => IR_OUT2s_14_port, IR_IN3(13) => 
                           IR_OUT2s_13_port, IR_IN3(12) => IR_OUT2s_12_port, 
                           IR_IN3(11) => IR_OUT2s_11_port, IR_IN3(10) => 
                           IR_OUT2s_10_port, IR_IN3(9) => IR_OUT2s_9_port, 
                           IR_IN3(8) => IR_OUT2s_8_port, IR_IN3(7) => 
                           IR_OUT2s_7_port, IR_IN3(6) => IR_OUT2s_6_port, 
                           IR_IN3(5) => IR_OUT2s_5_port, IR_IN3(4) => 
                           IR_OUT2s_4_port, IR_IN3(3) => IR_OUT2s_3_port, 
                           IR_IN3(2) => IR_OUT2s_2_port, IR_IN3(1) => 
                           IR_OUT2s_1_port, IR_IN3(0) => IR_OUT2s_0_port, 
                           IR_OUT3(31) => IR_OUT3s_31_port, IR_OUT3(30) => 
                           IR_OUT3s_30_port, IR_OUT3(29) => IR_OUT3s_29_port, 
                           IR_OUT3(28) => IR_OUT3s_28_port, IR_OUT3(27) => 
                           IR_OUT3s_27_port, IR_OUT3(26) => IR_OUT3s_26_port, 
                           IR_OUT3(25) => IR_OUT3s_25_port, IR_OUT3(24) => 
                           IR_OUT3s_24_port, IR_OUT3(23) => IR_OUT3s_23_port, 
                           IR_OUT3(22) => IR_OUT3s_22_port, IR_OUT3(21) => 
                           IR_OUT3s_21_port, IR_OUT3(20) => IR_OUT3s_20_port, 
                           IR_OUT3(19) => IR_OUT3s_19_port, IR_OUT3(18) => 
                           IR_OUT3s_18_port, IR_OUT3(17) => IR_OUT3s_17_port, 
                           IR_OUT3(16) => IR_OUT3s_16_port, IR_OUT3(15) => 
                           IR_OUT3s_15_port, IR_OUT3(14) => IR_OUT3s_14_port, 
                           IR_OUT3(13) => IR_OUT3s_13_port, IR_OUT3(12) => 
                           IR_OUT3s_12_port, IR_OUT3(11) => IR_OUT3s_11_port, 
                           IR_OUT3(10) => IR_OUT3s_10_port, IR_OUT3(9) => 
                           IR_OUT3s_9_port, IR_OUT3(8) => IR_OUT3s_8_port, 
                           IR_OUT3(7) => IR_OUT3s_7_port, IR_OUT3(6) => 
                           IR_OUT3s_6_port, IR_OUT3(5) => IR_OUT3s_5_port, 
                           IR_OUT3(4) => IR_OUT3s_4_port, IR_OUT3(3) => 
                           IR_OUT3s_3_port, IR_OUT3(2) => IR_OUT3s_2_port, 
                           IR_OUT3(1) => IR_OUT3s_1_port, IR_OUT3(0) => 
                           IR_OUT3s_0_port, B_outreg(31) => B(31), B_outreg(30)
                           => B(30), B_outreg(29) => B(29), B_outreg(28) => 
                           B(28), B_outreg(27) => B(27), B_outreg(26) => B(26),
                           B_outreg(25) => B(25), B_outreg(24) => B(24), 
                           B_outreg(23) => B(23), B_outreg(22) => B(22), 
                           B_outreg(21) => B(21), B_outreg(20) => B(20), 
                           B_outreg(19) => B(19), B_outreg(18) => B(18), 
                           B_outreg(17) => B(17), B_outreg(16) => B(16), 
                           B_outreg(15) => B(15), B_outreg(14) => B(14), 
                           B_outreg(13) => B(13), B_outreg(12) => B(12), 
                           B_outreg(11) => B(11), B_outreg(10) => B(10), 
                           B_outreg(9) => B(9), B_outreg(8) => B(8), 
                           B_outreg(7) => B(7), B_outreg(6) => B(6), 
                           B_outreg(5) => B(5), B_outreg(4) => B(4), 
                           B_outreg(3) => B(3), B_outreg(2) => B(2), 
                           B_outreg(1) => B(1), B_outreg(0) => B(0));
   MEMORY : memoryUnit_nbits32 port map( clk => n4, rst => n3, LMD_LATCH_EN => 
                           LMD_LATCH_EN, JUMP_EN => JUMP_EN, DRAM_DATA(31) => 
                           DRAM_DATA(31), DRAM_DATA(30) => DRAM_DATA(30), 
                           DRAM_DATA(29) => DRAM_DATA(29), DRAM_DATA(28) => 
                           DRAM_DATA(28), DRAM_DATA(27) => DRAM_DATA(27), 
                           DRAM_DATA(26) => DRAM_DATA(26), DRAM_DATA(25) => 
                           DRAM_DATA(25), DRAM_DATA(24) => DRAM_DATA(24), 
                           DRAM_DATA(23) => DRAM_DATA(23), DRAM_DATA(22) => 
                           DRAM_DATA(22), DRAM_DATA(21) => DRAM_DATA(21), 
                           DRAM_DATA(20) => DRAM_DATA(20), DRAM_DATA(19) => 
                           DRAM_DATA(19), DRAM_DATA(18) => DRAM_DATA(18), 
                           DRAM_DATA(17) => DRAM_DATA(17), DRAM_DATA(16) => 
                           DRAM_DATA(16), DRAM_DATA(15) => DRAM_DATA(15), 
                           DRAM_DATA(14) => DRAM_DATA(14), DRAM_DATA(13) => 
                           DRAM_DATA(13), DRAM_DATA(12) => DRAM_DATA(12), 
                           DRAM_DATA(11) => DRAM_DATA(11), DRAM_DATA(10) => 
                           DRAM_DATA(10), DRAM_DATA(9) => DRAM_DATA(9), 
                           DRAM_DATA(8) => DRAM_DATA(8), DRAM_DATA(7) => 
                           DRAM_DATA(7), DRAM_DATA(6) => DRAM_DATA(6), 
                           DRAM_DATA(5) => DRAM_DATA(5), DRAM_DATA(4) => 
                           DRAM_DATA(4), DRAM_DATA(3) => DRAM_DATA(3), 
                           DRAM_DATA(2) => DRAM_DATA(2), DRAM_DATA(1) => 
                           DRAM_DATA(1), DRAM_DATA(0) => DRAM_DATA(0), 
                           ALUREG_OUTPUT(31) => ALU_OUT_31_port, 
                           ALUREG_OUTPUT(30) => ALU_OUT_30_port, 
                           ALUREG_OUTPUT(29) => ALU_OUT_29_port, 
                           ALUREG_OUTPUT(28) => ALU_OUT_28_port, 
                           ALUREG_OUTPUT(27) => ALU_OUT_27_port, 
                           ALUREG_OUTPUT(26) => ALU_OUT_26_port, 
                           ALUREG_OUTPUT(25) => ALU_OUT_25_port, 
                           ALUREG_OUTPUT(24) => ALU_OUT_24_port, 
                           ALUREG_OUTPUT(23) => ALU_OUT_23_port, 
                           ALUREG_OUTPUT(22) => ALU_OUT_22_port, 
                           ALUREG_OUTPUT(21) => ALU_OUT_21_port, 
                           ALUREG_OUTPUT(20) => ALU_OUT_20_port, 
                           ALUREG_OUTPUT(19) => ALU_OUT_19_port, 
                           ALUREG_OUTPUT(18) => ALU_OUT_18_port, 
                           ALUREG_OUTPUT(17) => ALU_OUT_17_port, 
                           ALUREG_OUTPUT(16) => ALU_OUT_16_port, 
                           ALUREG_OUTPUT(15) => ALU_OUT_15_port, 
                           ALUREG_OUTPUT(14) => ALU_OUT_14_port, 
                           ALUREG_OUTPUT(13) => ALU_OUT_13_port, 
                           ALUREG_OUTPUT(12) => ALU_OUT_12_port, 
                           ALUREG_OUTPUT(11) => ALU_OUT_11_port, 
                           ALUREG_OUTPUT(10) => ALU_OUT_10_port, 
                           ALUREG_OUTPUT(9) => ALU_OUT_9_port, ALUREG_OUTPUT(8)
                           => ALU_OUT_8_port, ALUREG_OUTPUT(7) => 
                           ALU_OUT_7_port, ALUREG_OUTPUT(6) => ALU_OUT_6_port, 
                           ALUREG_OUTPUT(5) => ALU_OUT_5_port, ALUREG_OUTPUT(4)
                           => ALU_OUT_4_port, ALUREG_OUTPUT(3) => 
                           ALU_OUT_3_port, ALUREG_OUTPUT(2) => ALU_OUT_2_port, 
                           ALUREG_OUTPUT(1) => ALU_OUT_1_port, ALUREG_OUTPUT(0)
                           => ALU_OUT_0_port, NPC_OUT(31) => 
                           ADDERPC_OUTs_31_port, NPC_OUT(30) => 
                           ADDERPC_OUTs_30_port, NPC_OUT(29) => 
                           ADDERPC_OUTs_29_port, NPC_OUT(28) => 
                           ADDERPC_OUTs_28_port, NPC_OUT(27) => 
                           ADDERPC_OUTs_27_port, NPC_OUT(26) => 
                           ADDERPC_OUTs_26_port, NPC_OUT(25) => 
                           ADDERPC_OUTs_25_port, NPC_OUT(24) => 
                           ADDERPC_OUTs_24_port, NPC_OUT(23) => 
                           ADDERPC_OUTs_23_port, NPC_OUT(22) => 
                           ADDERPC_OUTs_22_port, NPC_OUT(21) => 
                           ADDERPC_OUTs_21_port, NPC_OUT(20) => 
                           ADDERPC_OUTs_20_port, NPC_OUT(19) => 
                           ADDERPC_OUTs_19_port, NPC_OUT(18) => 
                           ADDERPC_OUTs_18_port, NPC_OUT(17) => 
                           ADDERPC_OUTs_17_port, NPC_OUT(16) => 
                           ADDERPC_OUTs_16_port, NPC_OUT(15) => 
                           ADDERPC_OUTs_15_port, NPC_OUT(14) => 
                           ADDERPC_OUTs_14_port, NPC_OUT(13) => 
                           ADDERPC_OUTs_13_port, NPC_OUT(12) => 
                           ADDERPC_OUTs_12_port, NPC_OUT(11) => 
                           ADDERPC_OUTs_11_port, NPC_OUT(10) => 
                           ADDERPC_OUTs_10_port, NPC_OUT(9) => 
                           ADDERPC_OUTs_9_port, NPC_OUT(8) => 
                           ADDERPC_OUTs_8_port, NPC_OUT(7) => 
                           ADDERPC_OUTs_7_port, NPC_OUT(6) => 
                           ADDERPC_OUTs_6_port, NPC_OUT(5) => 
                           ADDERPC_OUTs_5_port, NPC_OUT(4) => 
                           ADDERPC_OUTs_4_port, NPC_OUT(3) => 
                           ADDERPC_OUTs_3_port, NPC_OUT(2) => 
                           ADDERPC_OUTs_2_port, NPC_OUT(1) => 
                           ADDERPC_OUTs_1_port, NPC_OUT(0) => 
                           ADDERPC_OUTs_0_port, COND_OUT => COND_OUTs, 
                           DRAM_DATAout(31) => LMD_OUTs_31_port, 
                           DRAM_DATAout(30) => LMD_OUTs_30_port, 
                           DRAM_DATAout(29) => LMD_OUTs_29_port, 
                           DRAM_DATAout(28) => LMD_OUTs_28_port, 
                           DRAM_DATAout(27) => LMD_OUTs_27_port, 
                           DRAM_DATAout(26) => LMD_OUTs_26_port, 
                           DRAM_DATAout(25) => LMD_OUTs_25_port, 
                           DRAM_DATAout(24) => LMD_OUTs_24_port, 
                           DRAM_DATAout(23) => LMD_OUTs_23_port, 
                           DRAM_DATAout(22) => LMD_OUTs_22_port, 
                           DRAM_DATAout(21) => LMD_OUTs_21_port, 
                           DRAM_DATAout(20) => LMD_OUTs_20_port, 
                           DRAM_DATAout(19) => LMD_OUTs_19_port, 
                           DRAM_DATAout(18) => LMD_OUTs_18_port, 
                           DRAM_DATAout(17) => LMD_OUTs_17_port, 
                           DRAM_DATAout(16) => LMD_OUTs_16_port, 
                           DRAM_DATAout(15) => LMD_OUTs_15_port, 
                           DRAM_DATAout(14) => LMD_OUTs_14_port, 
                           DRAM_DATAout(13) => LMD_OUTs_13_port, 
                           DRAM_DATAout(12) => LMD_OUTs_12_port, 
                           DRAM_DATAout(11) => LMD_OUTs_11_port, 
                           DRAM_DATAout(10) => LMD_OUTs_10_port, 
                           DRAM_DATAout(9) => LMD_OUTs_9_port, DRAM_DATAout(8) 
                           => LMD_OUTs_8_port, DRAM_DATAout(7) => 
                           LMD_OUTs_7_port, DRAM_DATAout(6) => LMD_OUTs_6_port,
                           DRAM_DATAout(5) => LMD_OUTs_5_port, DRAM_DATAout(4) 
                           => LMD_OUTs_4_port, DRAM_DATAout(3) => 
                           LMD_OUTs_3_port, DRAM_DATAout(2) => LMD_OUTs_2_port,
                           DRAM_DATAout(1) => LMD_OUTs_1_port, DRAM_DATAout(0) 
                           => LMD_OUTs_0_port, TO_PC_OUT(31) => 
                           TO_PC_OUTs_31_port, TO_PC_OUT(30) => 
                           TO_PC_OUTs_30_port, TO_PC_OUT(29) => 
                           TO_PC_OUTs_29_port, TO_PC_OUT(28) => 
                           TO_PC_OUTs_28_port, TO_PC_OUT(27) => 
                           TO_PC_OUTs_27_port, TO_PC_OUT(26) => 
                           TO_PC_OUTs_26_port, TO_PC_OUT(25) => 
                           TO_PC_OUTs_25_port, TO_PC_OUT(24) => 
                           TO_PC_OUTs_24_port, TO_PC_OUT(23) => 
                           TO_PC_OUTs_23_port, TO_PC_OUT(22) => 
                           TO_PC_OUTs_22_port, TO_PC_OUT(21) => 
                           TO_PC_OUTs_21_port, TO_PC_OUT(20) => 
                           TO_PC_OUTs_20_port, TO_PC_OUT(19) => 
                           TO_PC_OUTs_19_port, TO_PC_OUT(18) => 
                           TO_PC_OUTs_18_port, TO_PC_OUT(17) => 
                           TO_PC_OUTs_17_port, TO_PC_OUT(16) => 
                           TO_PC_OUTs_16_port, TO_PC_OUT(15) => 
                           TO_PC_OUTs_15_port, TO_PC_OUT(14) => 
                           TO_PC_OUTs_14_port, TO_PC_OUT(13) => 
                           TO_PC_OUTs_13_port, TO_PC_OUT(12) => 
                           TO_PC_OUTs_12_port, TO_PC_OUT(11) => 
                           TO_PC_OUTs_11_port, TO_PC_OUT(10) => 
                           TO_PC_OUTs_10_port, TO_PC_OUT(9) => 
                           TO_PC_OUTs_9_port, TO_PC_OUT(8) => TO_PC_OUTs_8_port
                           , TO_PC_OUT(7) => TO_PC_OUTs_7_port, TO_PC_OUT(6) =>
                           TO_PC_OUTs_6_port, TO_PC_OUT(5) => TO_PC_OUTs_5_port
                           , TO_PC_OUT(4) => TO_PC_OUTs_4_port, TO_PC_OUT(3) =>
                           TO_PC_OUTs_3_port, TO_PC_OUT(2) => TO_PC_OUTs_2_port
                           , TO_PC_OUT(1) => TO_PC_OUTs_1_port, TO_PC_OUT(0) =>
                           TO_PC_OUTs_0_port, ALU_OUT2(31) => ALU_OUT2s_31_port
                           , ALU_OUT2(30) => ALU_OUT2s_30_port, ALU_OUT2(29) =>
                           ALU_OUT2s_29_port, ALU_OUT2(28) => ALU_OUT2s_28_port
                           , ALU_OUT2(27) => ALU_OUT2s_27_port, ALU_OUT2(26) =>
                           ALU_OUT2s_26_port, ALU_OUT2(25) => ALU_OUT2s_25_port
                           , ALU_OUT2(24) => ALU_OUT2s_24_port, ALU_OUT2(23) =>
                           ALU_OUT2s_23_port, ALU_OUT2(22) => ALU_OUT2s_22_port
                           , ALU_OUT2(21) => ALU_OUT2s_21_port, ALU_OUT2(20) =>
                           ALU_OUT2s_20_port, ALU_OUT2(19) => ALU_OUT2s_19_port
                           , ALU_OUT2(18) => ALU_OUT2s_18_port, ALU_OUT2(17) =>
                           ALU_OUT2s_17_port, ALU_OUT2(16) => ALU_OUT2s_16_port
                           , ALU_OUT2(15) => ALU_OUT2s_15_port, ALU_OUT2(14) =>
                           ALU_OUT2s_14_port, ALU_OUT2(13) => ALU_OUT2s_13_port
                           , ALU_OUT2(12) => ALU_OUT2s_12_port, ALU_OUT2(11) =>
                           ALU_OUT2s_11_port, ALU_OUT2(10) => ALU_OUT2s_10_port
                           , ALU_OUT2(9) => ALU_OUT2s_9_port, ALU_OUT2(8) => 
                           ALU_OUT2s_8_port, ALU_OUT2(7) => ALU_OUT2s_7_port, 
                           ALU_OUT2(6) => ALU_OUT2s_6_port, ALU_OUT2(5) => 
                           ALU_OUT2s_5_port, ALU_OUT2(4) => ALU_OUT2s_4_port, 
                           ALU_OUT2(3) => ALU_OUT2s_3_port, ALU_OUT2(2) => 
                           ALU_OUT2s_2_port, ALU_OUT2(1) => ALU_OUT2s_1_port, 
                           ALU_OUT2(0) => ALU_OUT2s_0_port, IR_IN4(31) => 
                           IR_OUT3s_31_port, IR_IN4(30) => IR_OUT3s_30_port, 
                           IR_IN4(29) => IR_OUT3s_29_port, IR_IN4(28) => 
                           IR_OUT3s_28_port, IR_IN4(27) => IR_OUT3s_27_port, 
                           IR_IN4(26) => IR_OUT3s_26_port, IR_IN4(25) => 
                           IR_OUT3s_25_port, IR_IN4(24) => IR_OUT3s_24_port, 
                           IR_IN4(23) => IR_OUT3s_23_port, IR_IN4(22) => 
                           IR_OUT3s_22_port, IR_IN4(21) => IR_OUT3s_21_port, 
                           IR_IN4(20) => IR_OUT3s_20_port, IR_IN4(19) => 
                           IR_OUT3s_19_port, IR_IN4(18) => IR_OUT3s_18_port, 
                           IR_IN4(17) => IR_OUT3s_17_port, IR_IN4(16) => 
                           IR_OUT3s_16_port, IR_IN4(15) => IR_OUT3s_15_port, 
                           IR_IN4(14) => IR_OUT3s_14_port, IR_IN4(13) => 
                           IR_OUT3s_13_port, IR_IN4(12) => IR_OUT3s_12_port, 
                           IR_IN4(11) => IR_OUT3s_11_port, IR_IN4(10) => 
                           IR_OUT3s_10_port, IR_IN4(9) => IR_OUT3s_9_port, 
                           IR_IN4(8) => IR_OUT3s_8_port, IR_IN4(7) => 
                           IR_OUT3s_7_port, IR_IN4(6) => IR_OUT3s_6_port, 
                           IR_IN4(5) => IR_OUT3s_5_port, IR_IN4(4) => 
                           IR_OUT3s_4_port, IR_IN4(3) => IR_OUT3s_3_port, 
                           IR_IN4(2) => IR_OUT3s_2_port, IR_IN4(1) => 
                           IR_OUT3s_1_port, IR_IN4(0) => IR_OUT3s_0_port, 
                           IR_OUT4(31) => IR_OUT4s_31_port, IR_OUT4(30) => 
                           IR_OUT4s_30_port, IR_OUT4(29) => IR_OUT4s_29_port, 
                           IR_OUT4(28) => IR_OUT4s_28_port, IR_OUT4(27) => 
                           IR_OUT4s_27_port, IR_OUT4(26) => IR_OUT4s_26_port, 
                           IR_OUT4(25) => IR_OUT4s_25_port, IR_OUT4(24) => 
                           IR_OUT4s_24_port, IR_OUT4(23) => IR_OUT4s_23_port, 
                           IR_OUT4(22) => IR_OUT4s_22_port, IR_OUT4(21) => 
                           IR_OUT4s_21_port, IR_OUT4(20) => IR_OUT4s_20_port, 
                           IR_OUT4(19) => IR_OUT4s_19_port, IR_OUT4(18) => 
                           IR_OUT4s_18_port, IR_OUT4(17) => IR_OUT4s_17_port, 
                           IR_OUT4(16) => IR_OUT4s_16_port, IR_OUT4(15) => 
                           IR_OUT4s_15_port, IR_OUT4(14) => IR_OUT4s_14_port, 
                           IR_OUT4(13) => IR_OUT4s_13_port, IR_OUT4(12) => 
                           IR_OUT4s_12_port, IR_OUT4(11) => IR_OUT4s_11_port, 
                           IR_OUT4(10) => IR_OUT4s_10_port, IR_OUT4(9) => 
                           IR_OUT4s_9_port, IR_OUT4(8) => IR_OUT4s_8_port, 
                           IR_OUT4(7) => IR_OUT4s_7_port, IR_OUT4(6) => 
                           IR_OUT4s_6_port, IR_OUT4(5) => IR_OUT4s_5_port, 
                           IR_OUT4(4) => IR_OUT4s_4_port, IR_OUT4(3) => 
                           IR_OUT4s_3_port, IR_OUT4(2) => IR_OUT4s_2_port, 
                           IR_OUT4(1) => IR_OUT4s_1_port, IR_OUT4(0) => 
                           IR_OUT4s_0_port);
   WB : writeBack_nbits32 port map( LMD_OUT(31) => LMD_OUTs_31_port, 
                           LMD_OUT(30) => LMD_OUTs_30_port, LMD_OUT(29) => 
                           LMD_OUTs_29_port, LMD_OUT(28) => LMD_OUTs_28_port, 
                           LMD_OUT(27) => LMD_OUTs_27_port, LMD_OUT(26) => 
                           LMD_OUTs_26_port, LMD_OUT(25) => LMD_OUTs_25_port, 
                           LMD_OUT(24) => LMD_OUTs_24_port, LMD_OUT(23) => 
                           LMD_OUTs_23_port, LMD_OUT(22) => LMD_OUTs_22_port, 
                           LMD_OUT(21) => LMD_OUTs_21_port, LMD_OUT(20) => 
                           LMD_OUTs_20_port, LMD_OUT(19) => LMD_OUTs_19_port, 
                           LMD_OUT(18) => LMD_OUTs_18_port, LMD_OUT(17) => 
                           LMD_OUTs_17_port, LMD_OUT(16) => LMD_OUTs_16_port, 
                           LMD_OUT(15) => LMD_OUTs_15_port, LMD_OUT(14) => 
                           LMD_OUTs_14_port, LMD_OUT(13) => LMD_OUTs_13_port, 
                           LMD_OUT(12) => LMD_OUTs_12_port, LMD_OUT(11) => 
                           LMD_OUTs_11_port, LMD_OUT(10) => LMD_OUTs_10_port, 
                           LMD_OUT(9) => LMD_OUTs_9_port, LMD_OUT(8) => 
                           LMD_OUTs_8_port, LMD_OUT(7) => LMD_OUTs_7_port, 
                           LMD_OUT(6) => LMD_OUTs_6_port, LMD_OUT(5) => 
                           LMD_OUTs_5_port, LMD_OUT(4) => LMD_OUTs_4_port, 
                           LMD_OUT(3) => LMD_OUTs_3_port, LMD_OUT(2) => 
                           LMD_OUTs_2_port, LMD_OUT(1) => LMD_OUTs_1_port, 
                           LMD_OUT(0) => LMD_OUTs_0_port, ALUREG_OUTPUT(31) => 
                           ALU_OUT2s_31_port, ALUREG_OUTPUT(30) => 
                           ALU_OUT2s_30_port, ALUREG_OUTPUT(29) => 
                           ALU_OUT2s_29_port, ALUREG_OUTPUT(28) => 
                           ALU_OUT2s_28_port, ALUREG_OUTPUT(27) => 
                           ALU_OUT2s_27_port, ALUREG_OUTPUT(26) => 
                           ALU_OUT2s_26_port, ALUREG_OUTPUT(25) => 
                           ALU_OUT2s_25_port, ALUREG_OUTPUT(24) => 
                           ALU_OUT2s_24_port, ALUREG_OUTPUT(23) => 
                           ALU_OUT2s_23_port, ALUREG_OUTPUT(22) => 
                           ALU_OUT2s_22_port, ALUREG_OUTPUT(21) => 
                           ALU_OUT2s_21_port, ALUREG_OUTPUT(20) => 
                           ALU_OUT2s_20_port, ALUREG_OUTPUT(19) => 
                           ALU_OUT2s_19_port, ALUREG_OUTPUT(18) => 
                           ALU_OUT2s_18_port, ALUREG_OUTPUT(17) => 
                           ALU_OUT2s_17_port, ALUREG_OUTPUT(16) => 
                           ALU_OUT2s_16_port, ALUREG_OUTPUT(15) => 
                           ALU_OUT2s_15_port, ALUREG_OUTPUT(14) => 
                           ALU_OUT2s_14_port, ALUREG_OUTPUT(13) => 
                           ALU_OUT2s_13_port, ALUREG_OUTPUT(12) => 
                           ALU_OUT2s_12_port, ALUREG_OUTPUT(11) => 
                           ALU_OUT2s_11_port, ALUREG_OUTPUT(10) => 
                           ALU_OUT2s_10_port, ALUREG_OUTPUT(9) => 
                           ALU_OUT2s_9_port, ALUREG_OUTPUT(8) => 
                           ALU_OUT2s_8_port, ALUREG_OUTPUT(7) => 
                           ALU_OUT2s_7_port, ALUREG_OUTPUT(6) => 
                           ALU_OUT2s_6_port, ALUREG_OUTPUT(5) => 
                           ALU_OUT2s_5_port, ALUREG_OUTPUT(4) => 
                           ALU_OUT2s_4_port, ALUREG_OUTPUT(3) => 
                           ALU_OUT2s_3_port, ALUREG_OUTPUT(2) => 
                           ALU_OUT2s_2_port, ALUREG_OUTPUT(1) => 
                           ALU_OUT2s_1_port, ALUREG_OUTPUT(0) => 
                           ALU_OUT2s_0_port, WB_MUX_SEL => WB_MUX_SEL, 
                           DATAIN_RF(31) => DATAIN_RFs_31_port, DATAIN_RF(30) 
                           => DATAIN_RFs_30_port, DATAIN_RF(29) => 
                           DATAIN_RFs_29_port, DATAIN_RF(28) => 
                           DATAIN_RFs_28_port, DATAIN_RF(27) => 
                           DATAIN_RFs_27_port, DATAIN_RF(26) => 
                           DATAIN_RFs_26_port, DATAIN_RF(25) => 
                           DATAIN_RFs_25_port, DATAIN_RF(24) => 
                           DATAIN_RFs_24_port, DATAIN_RF(23) => 
                           DATAIN_RFs_23_port, DATAIN_RF(22) => 
                           DATAIN_RFs_22_port, DATAIN_RF(21) => 
                           DATAIN_RFs_21_port, DATAIN_RF(20) => 
                           DATAIN_RFs_20_port, DATAIN_RF(19) => 
                           DATAIN_RFs_19_port, DATAIN_RF(18) => 
                           DATAIN_RFs_18_port, DATAIN_RF(17) => 
                           DATAIN_RFs_17_port, DATAIN_RF(16) => 
                           DATAIN_RFs_16_port, DATAIN_RF(15) => 
                           DATAIN_RFs_15_port, DATAIN_RF(14) => 
                           DATAIN_RFs_14_port, DATAIN_RF(13) => 
                           DATAIN_RFs_13_port, DATAIN_RF(12) => 
                           DATAIN_RFs_12_port, DATAIN_RF(11) => 
                           DATAIN_RFs_11_port, DATAIN_RF(10) => 
                           DATAIN_RFs_10_port, DATAIN_RF(9) => 
                           DATAIN_RFs_9_port, DATAIN_RF(8) => DATAIN_RFs_8_port
                           , DATAIN_RF(7) => DATAIN_RFs_7_port, DATAIN_RF(6) =>
                           DATAIN_RFs_6_port, DATAIN_RF(5) => DATAIN_RFs_5_port
                           , DATAIN_RF(4) => DATAIN_RFs_4_port, DATAIN_RF(3) =>
                           DATAIN_RFs_3_port, DATAIN_RF(2) => DATAIN_RFs_2_port
                           , DATAIN_RF(1) => DATAIN_RFs_1_port, DATAIN_RF(0) =>
                           DATAIN_RFs_0_port);
   U1 : BUF_X1 port map( A => rst, Z => n3);
   U2 : BUF_X1 port map( A => clk, Z => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
         std_logic;  ALU_OPCODE : out std_logic_vector (0 to 3);  DRAM_WE, 
         LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, WB_MUX_SEL, RF_WE : out std_logic
         );

end dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, aluOpcode_i_3_port, aluOpcode_i_2_port, 
      aluOpcode_i_1_port, aluOpcode_i_0_port, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n_2045, 
      n_2046, n_2047, n_2048 : std_logic;

begin
   IR_LATCH_EN <= X_Logic1_port;
   NPC_LATCH_EN <= X_Logic1_port;
   PC_LATCH_EN <= X_Logic1_port;
   
   X_Logic1_port <= '1';
   RegIMM_LATCH_EN <= '0';
   RegB_LATCH_EN <= '0';
   RegA_LATCH_EN <= '0';
   aluOpcode1_reg_3_inst : DFFS_X1 port map( D => aluOpcode_i_3_port, CK => Clk
                           , SN => n59, Q => ALU_OPCODE(0), QN => n_2045);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => aluOpcode_i_2_port, CK => Clk
                           , RN => n59, Q => ALU_OPCODE(1), QN => n_2046);
   aluOpcode1_reg_1_inst : DFFS_X1 port map( D => aluOpcode_i_1_port, CK => Clk
                           , SN => n59, Q => ALU_OPCODE(2), QN => n_2047);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => aluOpcode_i_0_port, CK => Clk
                           , RN => n59, Q => ALU_OPCODE(3), QN => n_2048);
   RF_WE <= '0';
   WB_MUX_SEL <= '0';
   JUMP_EN <= '0';
   LMD_LATCH_EN <= '0';
   DRAM_WE <= '0';
   EQ_COND <= '0';
   ALU_OUTREG_EN <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   U3 : INV_X1 port map( A => Rst, ZN => n59);
   U13 : NAND3_X1 port map( A1 => n60, A2 => n61, A3 => n62, ZN => 
                           aluOpcode_i_3_port);
   U14 : AOI22_X1 port map( A1 => n63, A2 => IR_IN(2), B1 => IR_IN(28), B2 => 
                           n64, ZN => n62);
   U15 : OAI21_X1 port map( B1 => n65, B2 => n66, A => n67, ZN => n64);
   U16 : NOR2_X1 port map( A1 => n68, A2 => n69, ZN => n63);
   U17 : INV_X1 port map( A => n70, ZN => n61);
   U18 : XOR2_X1 port map( A => n71, B => n72, Z => n60);
   U19 : OAI211_X1 port map( C1 => n71, C2 => n73, A => n74, B => n75, ZN => 
                           aluOpcode_i_2_port);
   U20 : NAND3_X1 port map( A1 => n76, A2 => n77, A3 => n78, ZN => n74);
   U21 : MUX2_X1 port map( A => n79, B => n80, S => IR_IN(3), Z => n78);
   U22 : NOR3_X1 port map( A1 => n81, A2 => IR_IN(2), A3 => n82, ZN => n80);
   U23 : AOI21_X1 port map( B1 => n81, B2 => n83, A => n84, ZN => n79);
   U24 : NAND2_X1 port map( A1 => IR_IN(5), A2 => n82, ZN => n83);
   U25 : NAND4_X1 port map( A1 => n85, A2 => n86, A3 => n87, A4 => n88, ZN => 
                           aluOpcode_i_1_port);
   U26 : AND4_X1 port map( A1 => n72, A2 => n67, A3 => n89, A4 => n75, ZN => 
                           n88);
   U27 : INV_X1 port map( A => n71, ZN => n67);
   U28 : AOI21_X1 port map( B1 => n90, B2 => IR_IN(27), A => n70, ZN => n87);
   U29 : OAI21_X1 port map( B1 => n91, B2 => n69, A => n92, ZN => n70);
   U30 : MUX2_X1 port map( A => n93, B => n94, S => IR_IN(30), Z => n92);
   U31 : AOI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n94);
   U32 : MUX2_X1 port map( A => IR_IN(26), B => IR_IN(27), S => IR_IN(29), Z =>
                           n97);
   U33 : AOI22_X1 port map( A1 => n98, A2 => IR_IN(27), B1 => n99, B2 => n96, 
                           ZN => n93);
   U34 : NOR2_X1 port map( A1 => IR_IN(29), A2 => n71, ZN => n98);
   U35 : NOR2_X1 port map( A1 => n100, A2 => n95, ZN => n71);
   U36 : AND3_X1 port map( A1 => n77, A2 => n101, A3 => n102, ZN => n91);
   U37 : OAI21_X1 port map( B1 => IR_IN(0), B2 => IR_IN(3), A => n81, ZN => 
                           n102);
   U38 : INV_X1 port map( A => n103, ZN => n101);
   U39 : AOI21_X1 port map( B1 => n104, B2 => IR_IN(5), A => IR_IN(2), ZN => 
                           n103);
   U40 : XOR2_X1 port map( A => n82, B => IR_IN(3), Z => n104);
   U41 : INV_X1 port map( A => IR_IN(0), ZN => n82);
   U42 : OAI211_X1 port map( C1 => IR_IN(1), C2 => n84, A => IR_IN(5), B => n76
                           , ZN => n86);
   U43 : NAND3_X1 port map( A1 => n65, A2 => n66, A3 => IR_IN(28), ZN => n85);
   U44 : NAND3_X1 port map( A1 => n105, A2 => n75, A3 => n106, ZN => 
                           aluOpcode_i_0_port);
   U45 : AOI22_X1 port map( A1 => n107, A2 => n72, B1 => n90, B2 => n99, ZN => 
                           n106);
   U46 : INV_X1 port map( A => n108, ZN => n99);
   U47 : INV_X1 port map( A => n73, ZN => n90);
   U48 : NAND4_X1 port map( A1 => IR_IN(28), A2 => IR_IN(29), A3 => n66, A4 => 
                           n72, ZN => n73);
   U49 : INV_X1 port map( A => IR_IN(31), ZN => n72);
   U50 : OAI33_X1 port map( A1 => n109, A2 => n66, A3 => n96, B1 => n89, B2 => 
                           IR_IN(26), B3 => n100, ZN => n107);
   U51 : NAND3_X1 port map( A1 => n96, A2 => n66, A3 => IR_IN(29), ZN => n89);
   U52 : INV_X1 port map( A => IR_IN(28), ZN => n96);
   U53 : MUX2_X1 port map( A => n110, B => n108, S => IR_IN(29), Z => n109);
   U54 : NAND2_X1 port map( A1 => IR_IN(26), A2 => n100, ZN => n108);
   U55 : INV_X1 port map( A => IR_IN(27), ZN => n100);
   U56 : NAND2_X1 port map( A1 => IR_IN(27), A2 => n95, ZN => n110);
   U57 : NAND4_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), A3 => IR_IN(26), 
                           A4 => n111, ZN => n75);
   U58 : NAND3_X1 port map( A1 => n76, A2 => n77, A3 => n112, ZN => n105);
   U59 : MUX2_X1 port map( A => n113, B => n114, S => IR_IN(0), Z => n112);
   U60 : AOI21_X1 port map( B1 => n68, B2 => n84, A => n81, ZN => n114);
   U61 : NAND2_X1 port map( A1 => IR_IN(5), A2 => n115, ZN => n81);
   U62 : INV_X1 port map( A => IR_IN(3), ZN => n68);
   U63 : NOR3_X1 port map( A1 => n115, A2 => IR_IN(3), A3 => n116, ZN => n113);
   U64 : XOR2_X1 port map( A => IR_IN(5), B => n84, Z => n116);
   U65 : INV_X1 port map( A => IR_IN(2), ZN => n84);
   U66 : INV_X1 port map( A => IR_IN(1), ZN => n115);
   U67 : NOR4_X1 port map( A1 => IR_IN(6), A2 => IR_IN(4), A3 => IR_IN(10), A4 
                           => n117, ZN => n77);
   U68 : OR3_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), ZN =>
                           n117);
   U69 : INV_X1 port map( A => n69, ZN => n76);
   U70 : NAND4_X1 port map( A1 => n111, A2 => n95, A3 => n65, A4 => n66, ZN => 
                           n69);
   U71 : INV_X1 port map( A => IR_IN(30), ZN => n66);
   U72 : INV_X1 port map( A => IR_IN(29), ZN => n65);
   U73 : INV_X1 port map( A => IR_IN(26), ZN => n95);
   U74 : NOR3_X1 port map( A1 => IR_IN(28), A2 => IR_IN(31), A3 => IR_IN(27), 
                           ZN => n111);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity dlx is

   port( Clk_port, Rst_port : in std_logic;  DATA_IRAM_port, DATAread_DRAM_port
         : in std_logic_vector (31 downto 0);  WE_DRAM_port : out std_logic;  
         ADDRESS_DRAM_port, DATAwrite_DRAM_port, ADDRESS_IRAM_port : out 
         std_logic_vector (31 downto 0));

end dlx;

architecture SYN_STRUCTURAL of dlx is

   component datapath_nbits32
      port( clk, rst : in std_logic;  DATA_IRAM : in std_logic_vector (31 
            downto 0);  IR_LATCH_EN, NPC_LATCH_EN, PC_LATCH_EN, RegA_LATCH_EN, 
            RegB_LATCH_EN, RegIMM_LATCH_EN, RF_WE, MUXA_SEL, MUXB_SEL, 
            ALU_OUTREG_EN, EQ_COND : in std_logic;  ALU_OPCODE : in 
            std_logic_vector (0 to 3);  DRAM_DATA : in std_logic_vector (31 
            downto 0);  LMD_LATCH_EN, JUMP_EN, WB_MUX_SEL : in std_logic;  B, 
            ALU_OUT, ADDRESS_IRAM, IR_OUT : out std_logic_vector (31 downto 0)
            );
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
            std_logic;  ALU_OPCODE : out std_logic_vector (0 to 3);  DRAM_WE, 
            LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, WB_MUX_SEL, RF_WE : out 
            std_logic);
   end component;
   
   signal IR_OUT_signal_31_port, IR_OUT_signal_30_port, IR_OUT_signal_29_port, 
      IR_OUT_signal_28_port, IR_OUT_signal_27_port, IR_OUT_signal_26_port, 
      IR_OUT_signal_25_port, IR_OUT_signal_24_port, IR_OUT_signal_23_port, 
      IR_OUT_signal_22_port, IR_OUT_signal_21_port, IR_OUT_signal_20_port, 
      IR_OUT_signal_19_port, IR_OUT_signal_18_port, IR_OUT_signal_17_port, 
      IR_OUT_signal_16_port, IR_OUT_signal_15_port, IR_OUT_signal_14_port, 
      IR_OUT_signal_13_port, IR_OUT_signal_12_port, IR_OUT_signal_11_port, 
      IR_OUT_signal_10_port, IR_OUT_signal_9_port, IR_OUT_signal_8_port, 
      IR_OUT_signal_7_port, IR_OUT_signal_6_port, IR_OUT_signal_5_port, 
      IR_OUT_signal_4_port, IR_OUT_signal_3_port, IR_OUT_signal_2_port, 
      IR_OUT_signal_1_port, IR_OUT_signal_0_port, IR_LATCH_EN_signal, 
      NPC_LATCH_EN_signal, RegA_LATCH_EN_signal, RegB_LATCH_EN_signal, 
      RegIMM_LATCH_EN_signal, MUXA_SEL_signal, MUXB_SEL_signal, 
      ALU_OUTREG_EN_signal, EQ_COND_signal, ALU_OPCODE_signal_0_port, 
      ALU_OPCODE_signal_1_port, ALU_OPCODE_signal_2_port, 
      ALU_OPCODE_signal_3_port, LMD_LATCH_EN_signal, JUMP_EN_signal, 
      PC_LATCH_EN_signal, WB_MUX_SEL_signal, RF_WE_signal, n_2049, n_2050, 
      n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, 
      n_2060, n_2061, n_2062, n_2063 : std_logic;

begin
   
   RF_WE_signal <= '0';
   WB_MUX_SEL_signal <= '0';
   PC_LATCH_EN_signal <= '1';
   JUMP_EN_signal <= '0';
   LMD_LATCH_EN_signal <= '0';
   WE_DRAM_port <= '0';
   EQ_COND_signal <= '0';
   ALU_OUTREG_EN_signal <= '0';
   MUXB_SEL_signal <= '0';
   MUXA_SEL_signal <= '0';
   RegIMM_LATCH_EN_signal <= '0';
   RegB_LATCH_EN_signal <= '0';
   RegA_LATCH_EN_signal <= '0';
   NPC_LATCH_EN_signal <= '1';
   IR_LATCH_EN_signal <= '1';
   CONTROL_UNIT : 
                           dlx_cu_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 
                           port map( Clk => Clk_port, Rst => Rst_port, 
                           IR_IN(31) => IR_OUT_signal_31_port, IR_IN(30) => 
                           IR_OUT_signal_30_port, IR_IN(29) => 
                           IR_OUT_signal_29_port, IR_IN(28) => 
                           IR_OUT_signal_28_port, IR_IN(27) => 
                           IR_OUT_signal_27_port, IR_IN(26) => 
                           IR_OUT_signal_26_port, IR_IN(25) => 
                           IR_OUT_signal_25_port, IR_IN(24) => 
                           IR_OUT_signal_24_port, IR_IN(23) => 
                           IR_OUT_signal_23_port, IR_IN(22) => 
                           IR_OUT_signal_22_port, IR_IN(21) => 
                           IR_OUT_signal_21_port, IR_IN(20) => 
                           IR_OUT_signal_20_port, IR_IN(19) => 
                           IR_OUT_signal_19_port, IR_IN(18) => 
                           IR_OUT_signal_18_port, IR_IN(17) => 
                           IR_OUT_signal_17_port, IR_IN(16) => 
                           IR_OUT_signal_16_port, IR_IN(15) => 
                           IR_OUT_signal_15_port, IR_IN(14) => 
                           IR_OUT_signal_14_port, IR_IN(13) => 
                           IR_OUT_signal_13_port, IR_IN(12) => 
                           IR_OUT_signal_12_port, IR_IN(11) => 
                           IR_OUT_signal_11_port, IR_IN(10) => 
                           IR_OUT_signal_10_port, IR_IN(9) => 
                           IR_OUT_signal_9_port, IR_IN(8) => 
                           IR_OUT_signal_8_port, IR_IN(7) => 
                           IR_OUT_signal_7_port, IR_IN(6) => 
                           IR_OUT_signal_6_port, IR_IN(5) => 
                           IR_OUT_signal_5_port, IR_IN(4) => 
                           IR_OUT_signal_4_port, IR_IN(3) => 
                           IR_OUT_signal_3_port, IR_IN(2) => 
                           IR_OUT_signal_2_port, IR_IN(1) => 
                           IR_OUT_signal_1_port, IR_IN(0) => 
                           IR_OUT_signal_0_port, IR_LATCH_EN => n_2049, 
                           NPC_LATCH_EN => n_2050, RegA_LATCH_EN => n_2051, 
                           RegB_LATCH_EN => n_2052, RegIMM_LATCH_EN => n_2053, 
                           MUXA_SEL => n_2054, MUXB_SEL => n_2055, 
                           ALU_OUTREG_EN => n_2056, EQ_COND => n_2057, 
                           ALU_OPCODE(0) => ALU_OPCODE_signal_0_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_signal_1_port, 
                           ALU_OPCODE(2) => ALU_OPCODE_signal_2_port, 
                           ALU_OPCODE(3) => ALU_OPCODE_signal_3_port, DRAM_WE 
                           => n_2058, LMD_LATCH_EN => n_2059, JUMP_EN => n_2060
                           , PC_LATCH_EN => n_2061, WB_MUX_SEL => n_2062, RF_WE
                           => n_2063);
   DATA_PATH : datapath_nbits32 port map( clk => Clk_port, rst => Rst_port, 
                           DATA_IRAM(31) => DATA_IRAM_port(31), DATA_IRAM(30) 
                           => DATA_IRAM_port(30), DATA_IRAM(29) => 
                           DATA_IRAM_port(29), DATA_IRAM(28) => 
                           DATA_IRAM_port(28), DATA_IRAM(27) => 
                           DATA_IRAM_port(27), DATA_IRAM(26) => 
                           DATA_IRAM_port(26), DATA_IRAM(25) => 
                           DATA_IRAM_port(25), DATA_IRAM(24) => 
                           DATA_IRAM_port(24), DATA_IRAM(23) => 
                           DATA_IRAM_port(23), DATA_IRAM(22) => 
                           DATA_IRAM_port(22), DATA_IRAM(21) => 
                           DATA_IRAM_port(21), DATA_IRAM(20) => 
                           DATA_IRAM_port(20), DATA_IRAM(19) => 
                           DATA_IRAM_port(19), DATA_IRAM(18) => 
                           DATA_IRAM_port(18), DATA_IRAM(17) => 
                           DATA_IRAM_port(17), DATA_IRAM(16) => 
                           DATA_IRAM_port(16), DATA_IRAM(15) => 
                           DATA_IRAM_port(15), DATA_IRAM(14) => 
                           DATA_IRAM_port(14), DATA_IRAM(13) => 
                           DATA_IRAM_port(13), DATA_IRAM(12) => 
                           DATA_IRAM_port(12), DATA_IRAM(11) => 
                           DATA_IRAM_port(11), DATA_IRAM(10) => 
                           DATA_IRAM_port(10), DATA_IRAM(9) => 
                           DATA_IRAM_port(9), DATA_IRAM(8) => DATA_IRAM_port(8)
                           , DATA_IRAM(7) => DATA_IRAM_port(7), DATA_IRAM(6) =>
                           DATA_IRAM_port(6), DATA_IRAM(5) => DATA_IRAM_port(5)
                           , DATA_IRAM(4) => DATA_IRAM_port(4), DATA_IRAM(3) =>
                           DATA_IRAM_port(3), DATA_IRAM(2) => DATA_IRAM_port(2)
                           , DATA_IRAM(1) => DATA_IRAM_port(1), DATA_IRAM(0) =>
                           DATA_IRAM_port(0), IR_LATCH_EN => IR_LATCH_EN_signal
                           , NPC_LATCH_EN => NPC_LATCH_EN_signal, PC_LATCH_EN 
                           => PC_LATCH_EN_signal, RegA_LATCH_EN => 
                           RegA_LATCH_EN_signal, RegB_LATCH_EN => 
                           RegB_LATCH_EN_signal, RegIMM_LATCH_EN => 
                           RegIMM_LATCH_EN_signal, RF_WE => RF_WE_signal, 
                           MUXA_SEL => MUXA_SEL_signal, MUXB_SEL => 
                           MUXB_SEL_signal, ALU_OUTREG_EN => 
                           ALU_OUTREG_EN_signal, EQ_COND => EQ_COND_signal, 
                           ALU_OPCODE(0) => ALU_OPCODE_signal_0_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_signal_1_port, 
                           ALU_OPCODE(2) => ALU_OPCODE_signal_2_port, 
                           ALU_OPCODE(3) => ALU_OPCODE_signal_3_port, 
                           DRAM_DATA(31) => DATAread_DRAM_port(31), 
                           DRAM_DATA(30) => DATAread_DRAM_port(30), 
                           DRAM_DATA(29) => DATAread_DRAM_port(29), 
                           DRAM_DATA(28) => DATAread_DRAM_port(28), 
                           DRAM_DATA(27) => DATAread_DRAM_port(27), 
                           DRAM_DATA(26) => DATAread_DRAM_port(26), 
                           DRAM_DATA(25) => DATAread_DRAM_port(25), 
                           DRAM_DATA(24) => DATAread_DRAM_port(24), 
                           DRAM_DATA(23) => DATAread_DRAM_port(23), 
                           DRAM_DATA(22) => DATAread_DRAM_port(22), 
                           DRAM_DATA(21) => DATAread_DRAM_port(21), 
                           DRAM_DATA(20) => DATAread_DRAM_port(20), 
                           DRAM_DATA(19) => DATAread_DRAM_port(19), 
                           DRAM_DATA(18) => DATAread_DRAM_port(18), 
                           DRAM_DATA(17) => DATAread_DRAM_port(17), 
                           DRAM_DATA(16) => DATAread_DRAM_port(16), 
                           DRAM_DATA(15) => DATAread_DRAM_port(15), 
                           DRAM_DATA(14) => DATAread_DRAM_port(14), 
                           DRAM_DATA(13) => DATAread_DRAM_port(13), 
                           DRAM_DATA(12) => DATAread_DRAM_port(12), 
                           DRAM_DATA(11) => DATAread_DRAM_port(11), 
                           DRAM_DATA(10) => DATAread_DRAM_port(10), 
                           DRAM_DATA(9) => DATAread_DRAM_port(9), DRAM_DATA(8) 
                           => DATAread_DRAM_port(8), DRAM_DATA(7) => 
                           DATAread_DRAM_port(7), DRAM_DATA(6) => 
                           DATAread_DRAM_port(6), DRAM_DATA(5) => 
                           DATAread_DRAM_port(5), DRAM_DATA(4) => 
                           DATAread_DRAM_port(4), DRAM_DATA(3) => 
                           DATAread_DRAM_port(3), DRAM_DATA(2) => 
                           DATAread_DRAM_port(2), DRAM_DATA(1) => 
                           DATAread_DRAM_port(1), DRAM_DATA(0) => 
                           DATAread_DRAM_port(0), LMD_LATCH_EN => 
                           LMD_LATCH_EN_signal, JUMP_EN => JUMP_EN_signal, 
                           WB_MUX_SEL => WB_MUX_SEL_signal, B(31) => 
                           DATAwrite_DRAM_port(31), B(30) => 
                           DATAwrite_DRAM_port(30), B(29) => 
                           DATAwrite_DRAM_port(29), B(28) => 
                           DATAwrite_DRAM_port(28), B(27) => 
                           DATAwrite_DRAM_port(27), B(26) => 
                           DATAwrite_DRAM_port(26), B(25) => 
                           DATAwrite_DRAM_port(25), B(24) => 
                           DATAwrite_DRAM_port(24), B(23) => 
                           DATAwrite_DRAM_port(23), B(22) => 
                           DATAwrite_DRAM_port(22), B(21) => 
                           DATAwrite_DRAM_port(21), B(20) => 
                           DATAwrite_DRAM_port(20), B(19) => 
                           DATAwrite_DRAM_port(19), B(18) => 
                           DATAwrite_DRAM_port(18), B(17) => 
                           DATAwrite_DRAM_port(17), B(16) => 
                           DATAwrite_DRAM_port(16), B(15) => 
                           DATAwrite_DRAM_port(15), B(14) => 
                           DATAwrite_DRAM_port(14), B(13) => 
                           DATAwrite_DRAM_port(13), B(12) => 
                           DATAwrite_DRAM_port(12), B(11) => 
                           DATAwrite_DRAM_port(11), B(10) => 
                           DATAwrite_DRAM_port(10), B(9) => 
                           DATAwrite_DRAM_port(9), B(8) => 
                           DATAwrite_DRAM_port(8), B(7) => 
                           DATAwrite_DRAM_port(7), B(6) => 
                           DATAwrite_DRAM_port(6), B(5) => 
                           DATAwrite_DRAM_port(5), B(4) => 
                           DATAwrite_DRAM_port(4), B(3) => 
                           DATAwrite_DRAM_port(3), B(2) => 
                           DATAwrite_DRAM_port(2), B(1) => 
                           DATAwrite_DRAM_port(1), B(0) => 
                           DATAwrite_DRAM_port(0), ALU_OUT(31) => 
                           ADDRESS_DRAM_port(31), ALU_OUT(30) => 
                           ADDRESS_DRAM_port(30), ALU_OUT(29) => 
                           ADDRESS_DRAM_port(29), ALU_OUT(28) => 
                           ADDRESS_DRAM_port(28), ALU_OUT(27) => 
                           ADDRESS_DRAM_port(27), ALU_OUT(26) => 
                           ADDRESS_DRAM_port(26), ALU_OUT(25) => 
                           ADDRESS_DRAM_port(25), ALU_OUT(24) => 
                           ADDRESS_DRAM_port(24), ALU_OUT(23) => 
                           ADDRESS_DRAM_port(23), ALU_OUT(22) => 
                           ADDRESS_DRAM_port(22), ALU_OUT(21) => 
                           ADDRESS_DRAM_port(21), ALU_OUT(20) => 
                           ADDRESS_DRAM_port(20), ALU_OUT(19) => 
                           ADDRESS_DRAM_port(19), ALU_OUT(18) => 
                           ADDRESS_DRAM_port(18), ALU_OUT(17) => 
                           ADDRESS_DRAM_port(17), ALU_OUT(16) => 
                           ADDRESS_DRAM_port(16), ALU_OUT(15) => 
                           ADDRESS_DRAM_port(15), ALU_OUT(14) => 
                           ADDRESS_DRAM_port(14), ALU_OUT(13) => 
                           ADDRESS_DRAM_port(13), ALU_OUT(12) => 
                           ADDRESS_DRAM_port(12), ALU_OUT(11) => 
                           ADDRESS_DRAM_port(11), ALU_OUT(10) => 
                           ADDRESS_DRAM_port(10), ALU_OUT(9) => 
                           ADDRESS_DRAM_port(9), ALU_OUT(8) => 
                           ADDRESS_DRAM_port(8), ALU_OUT(7) => 
                           ADDRESS_DRAM_port(7), ALU_OUT(6) => 
                           ADDRESS_DRAM_port(6), ALU_OUT(5) => 
                           ADDRESS_DRAM_port(5), ALU_OUT(4) => 
                           ADDRESS_DRAM_port(4), ALU_OUT(3) => 
                           ADDRESS_DRAM_port(3), ALU_OUT(2) => 
                           ADDRESS_DRAM_port(2), ALU_OUT(1) => 
                           ADDRESS_DRAM_port(1), ALU_OUT(0) => 
                           ADDRESS_DRAM_port(0), ADDRESS_IRAM(31) => 
                           ADDRESS_IRAM_port(31), ADDRESS_IRAM(30) => 
                           ADDRESS_IRAM_port(30), ADDRESS_IRAM(29) => 
                           ADDRESS_IRAM_port(29), ADDRESS_IRAM(28) => 
                           ADDRESS_IRAM_port(28), ADDRESS_IRAM(27) => 
                           ADDRESS_IRAM_port(27), ADDRESS_IRAM(26) => 
                           ADDRESS_IRAM_port(26), ADDRESS_IRAM(25) => 
                           ADDRESS_IRAM_port(25), ADDRESS_IRAM(24) => 
                           ADDRESS_IRAM_port(24), ADDRESS_IRAM(23) => 
                           ADDRESS_IRAM_port(23), ADDRESS_IRAM(22) => 
                           ADDRESS_IRAM_port(22), ADDRESS_IRAM(21) => 
                           ADDRESS_IRAM_port(21), ADDRESS_IRAM(20) => 
                           ADDRESS_IRAM_port(20), ADDRESS_IRAM(19) => 
                           ADDRESS_IRAM_port(19), ADDRESS_IRAM(18) => 
                           ADDRESS_IRAM_port(18), ADDRESS_IRAM(17) => 
                           ADDRESS_IRAM_port(17), ADDRESS_IRAM(16) => 
                           ADDRESS_IRAM_port(16), ADDRESS_IRAM(15) => 
                           ADDRESS_IRAM_port(15), ADDRESS_IRAM(14) => 
                           ADDRESS_IRAM_port(14), ADDRESS_IRAM(13) => 
                           ADDRESS_IRAM_port(13), ADDRESS_IRAM(12) => 
                           ADDRESS_IRAM_port(12), ADDRESS_IRAM(11) => 
                           ADDRESS_IRAM_port(11), ADDRESS_IRAM(10) => 
                           ADDRESS_IRAM_port(10), ADDRESS_IRAM(9) => 
                           ADDRESS_IRAM_port(9), ADDRESS_IRAM(8) => 
                           ADDRESS_IRAM_port(8), ADDRESS_IRAM(7) => 
                           ADDRESS_IRAM_port(7), ADDRESS_IRAM(6) => 
                           ADDRESS_IRAM_port(6), ADDRESS_IRAM(5) => 
                           ADDRESS_IRAM_port(5), ADDRESS_IRAM(4) => 
                           ADDRESS_IRAM_port(4), ADDRESS_IRAM(3) => 
                           ADDRESS_IRAM_port(3), ADDRESS_IRAM(2) => 
                           ADDRESS_IRAM_port(2), ADDRESS_IRAM(1) => 
                           ADDRESS_IRAM_port(1), ADDRESS_IRAM(0) => 
                           ADDRESS_IRAM_port(0), IR_OUT(31) => 
                           IR_OUT_signal_31_port, IR_OUT(30) => 
                           IR_OUT_signal_30_port, IR_OUT(29) => 
                           IR_OUT_signal_29_port, IR_OUT(28) => 
                           IR_OUT_signal_28_port, IR_OUT(27) => 
                           IR_OUT_signal_27_port, IR_OUT(26) => 
                           IR_OUT_signal_26_port, IR_OUT(25) => 
                           IR_OUT_signal_25_port, IR_OUT(24) => 
                           IR_OUT_signal_24_port, IR_OUT(23) => 
                           IR_OUT_signal_23_port, IR_OUT(22) => 
                           IR_OUT_signal_22_port, IR_OUT(21) => 
                           IR_OUT_signal_21_port, IR_OUT(20) => 
                           IR_OUT_signal_20_port, IR_OUT(19) => 
                           IR_OUT_signal_19_port, IR_OUT(18) => 
                           IR_OUT_signal_18_port, IR_OUT(17) => 
                           IR_OUT_signal_17_port, IR_OUT(16) => 
                           IR_OUT_signal_16_port, IR_OUT(15) => 
                           IR_OUT_signal_15_port, IR_OUT(14) => 
                           IR_OUT_signal_14_port, IR_OUT(13) => 
                           IR_OUT_signal_13_port, IR_OUT(12) => 
                           IR_OUT_signal_12_port, IR_OUT(11) => 
                           IR_OUT_signal_11_port, IR_OUT(10) => 
                           IR_OUT_signal_10_port, IR_OUT(9) => 
                           IR_OUT_signal_9_port, IR_OUT(8) => 
                           IR_OUT_signal_8_port, IR_OUT(7) => 
                           IR_OUT_signal_7_port, IR_OUT(6) => 
                           IR_OUT_signal_6_port, IR_OUT(5) => 
                           IR_OUT_signal_5_port, IR_OUT(4) => 
                           IR_OUT_signal_4_port, IR_OUT(3) => 
                           IR_OUT_signal_3_port, IR_OUT(2) => 
                           IR_OUT_signal_2_port, IR_OUT(1) => 
                           IR_OUT_signal_1_port, IR_OUT(0) => 
                           IR_OUT_signal_0_port);

end SYN_STRUCTURAL;
